

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733;

  INV_X2 U372 ( .A(n573), .ZN(n619) );
  OR2_X2 U373 ( .A1(n660), .A2(n573), .ZN(n487) );
  XNOR2_X2 U374 ( .A(n520), .B(KEYINPUT32), .ZN(n733) );
  XOR2_X2 U375 ( .A(n376), .B(n375), .Z(n533) );
  XNOR2_X2 U376 ( .A(n512), .B(n511), .ZN(n732) );
  OR2_X1 U377 ( .A1(n501), .A2(n664), .ZN(n417) );
  INV_X1 U378 ( .A(n702), .ZN(n351) );
  AND2_X2 U379 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U380 ( .A(n455), .B(n454), .ZN(n656) );
  XNOR2_X1 U381 ( .A(n437), .B(n436), .ZN(n683) );
  XNOR2_X1 U382 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n396) );
  XNOR2_X2 U383 ( .A(n487), .B(n486), .ZN(n565) );
  NOR2_X1 U384 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U385 ( .A1(n647), .A2(n646), .ZN(n650) );
  XNOR2_X1 U386 ( .A(n465), .B(KEYINPUT94), .ZN(n359) );
  XNOR2_X1 U387 ( .A(G119), .B(G128), .ZN(n456) );
  XNOR2_X1 U388 ( .A(n372), .B(n371), .ZN(n461) );
  NAND2_X2 U389 ( .A1(n363), .A2(n362), .ZN(n687) );
  NAND2_X1 U390 ( .A1(n641), .A2(n356), .ZN(n362) );
  NAND2_X1 U391 ( .A1(n353), .A2(n364), .ZN(n363) );
  INV_X1 U392 ( .A(KEYINPUT45), .ZN(n554) );
  NOR2_X1 U393 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U394 ( .A1(G902), .A2(n693), .ZN(n375) );
  BUF_X1 U395 ( .A(n687), .Z(n697) );
  XNOR2_X1 U396 ( .A(n435), .B(n434), .ZN(n436) );
  AND2_X1 U397 ( .A1(n477), .A2(n596), .ZN(n701) );
  NOR2_X1 U398 ( .A1(n575), .A2(n620), .ZN(n576) );
  XOR2_X1 U399 ( .A(KEYINPUT96), .B(G131), .Z(n443) );
  XNOR2_X1 U400 ( .A(G137), .B(G116), .ZN(n442) );
  XOR2_X1 U401 ( .A(KEYINPUT4), .B(KEYINPUT67), .Z(n719) );
  INV_X1 U402 ( .A(G146), .ZN(n429) );
  XOR2_X1 U403 ( .A(G131), .B(G140), .Z(n432) );
  XNOR2_X1 U404 ( .A(n638), .B(KEYINPUT78), .ZN(n364) );
  NOR2_X1 U405 ( .A1(n590), .A2(KEYINPUT2), .ZN(n361) );
  XNOR2_X1 U406 ( .A(n429), .B(G125), .ZN(n400) );
  OR2_X1 U407 ( .A1(n550), .A2(KEYINPUT89), .ZN(n551) );
  XNOR2_X1 U408 ( .A(n718), .B(n429), .ZN(n444) );
  NAND2_X1 U409 ( .A1(n351), .A2(n589), .ZN(n641) );
  XNOR2_X1 U410 ( .A(n453), .B(G472), .ZN(n454) );
  NOR2_X1 U411 ( .A1(n650), .A2(n496), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n360), .B(n358), .ZN(n698) );
  XNOR2_X1 U413 ( .A(n359), .B(n354), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n460), .B(n464), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n374), .B(n373), .ZN(n693) );
  XNOR2_X1 U416 ( .A(n564), .B(n563), .ZN(n731) );
  OR2_X1 U417 ( .A1(n584), .A2(n561), .ZN(n564) );
  AND2_X1 U418 ( .A1(n510), .A2(n509), .ZN(n512) );
  XNOR2_X1 U419 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U420 ( .A(n683), .B(n682), .ZN(n684) );
  OR2_X1 U421 ( .A1(n698), .A2(G902), .ZN(n352) );
  AND2_X1 U422 ( .A1(n351), .A2(n361), .ZN(n353) );
  XOR2_X1 U423 ( .A(n463), .B(n462), .Z(n354) );
  XNOR2_X1 U424 ( .A(G107), .B(KEYINPUT7), .ZN(n355) );
  INV_X1 U425 ( .A(n590), .ZN(n591) );
  AND2_X1 U426 ( .A1(n591), .A2(KEYINPUT2), .ZN(n356) );
  NAND2_X1 U427 ( .A1(n357), .A2(n528), .ZN(n529) );
  NAND2_X1 U428 ( .A1(n500), .A2(n357), .ZN(n559) );
  XNOR2_X1 U429 ( .A(n433), .B(n717), .ZN(n434) );
  XNOR2_X2 U430 ( .A(n417), .B(KEYINPUT19), .ZN(n574) );
  NOR2_X1 U431 ( .A1(n649), .A2(n650), .ZN(n503) );
  XNOR2_X2 U432 ( .A(n428), .B(n427), .ZN(n539) );
  XOR2_X1 U433 ( .A(n468), .B(n467), .Z(n365) );
  OR2_X1 U434 ( .A1(n557), .A2(n559), .ZN(n366) );
  XNOR2_X1 U435 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n383) );
  XNOR2_X1 U436 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n498) );
  INV_X1 U437 ( .A(G134), .ZN(n367) );
  XNOR2_X1 U438 ( .A(n431), .B(KEYINPUT80), .ZN(n433) );
  XNOR2_X1 U439 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U440 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U441 ( .A(KEYINPUT87), .ZN(n588) );
  XNOR2_X1 U442 ( .A(n370), .B(n355), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n438), .B(G469), .ZN(n439) );
  XNOR2_X1 U444 ( .A(n693), .B(KEYINPUT122), .ZN(n694) );
  XNOR2_X1 U445 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U446 ( .A(KEYINPUT103), .B(G478), .ZN(n376) );
  XOR2_X2 U447 ( .A(G143), .B(G128), .Z(n398) );
  XNOR2_X2 U448 ( .A(n398), .B(n367), .ZN(n718) );
  XOR2_X1 U449 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n368) );
  XNOR2_X1 U450 ( .A(G122), .B(G116), .ZN(n406) );
  XOR2_X1 U451 ( .A(n368), .B(n406), .Z(n369) );
  XNOR2_X1 U452 ( .A(n718), .B(n369), .ZN(n370) );
  XOR2_X1 U453 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n372) );
  XNOR2_X2 U454 ( .A(KEYINPUT64), .B(G953), .ZN(n477) );
  INV_X1 U455 ( .A(n477), .ZN(n722) );
  NAND2_X1 U456 ( .A1(G234), .A2(n722), .ZN(n371) );
  NAND2_X1 U457 ( .A1(G217), .A2(n461), .ZN(n373) );
  XNOR2_X1 U458 ( .A(KEYINPUT13), .B(G475), .ZN(n389) );
  XOR2_X1 U459 ( .A(G113), .B(G104), .Z(n378) );
  NOR2_X1 U460 ( .A1(G953), .A2(G237), .ZN(n446) );
  NAND2_X1 U461 ( .A1(G214), .A2(n446), .ZN(n377) );
  XNOR2_X1 U462 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U463 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n380) );
  XNOR2_X1 U464 ( .A(KEYINPUT11), .B(KEYINPUT101), .ZN(n379) );
  XNOR2_X1 U465 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U466 ( .A(n382), .B(n381), .Z(n387) );
  XNOR2_X1 U467 ( .A(n400), .B(n383), .ZN(n458) );
  XNOR2_X1 U468 ( .A(G143), .B(G122), .ZN(n384) );
  XNOR2_X1 U469 ( .A(n384), .B(n432), .ZN(n385) );
  XNOR2_X1 U470 ( .A(n458), .B(n385), .ZN(n386) );
  XNOR2_X1 U471 ( .A(n387), .B(n386), .ZN(n688) );
  NOR2_X1 U472 ( .A1(G902), .A2(n688), .ZN(n388) );
  XNOR2_X1 U473 ( .A(n389), .B(n388), .ZN(n532) );
  INV_X1 U474 ( .A(n532), .ZN(n390) );
  NAND2_X1 U475 ( .A1(n533), .A2(n390), .ZN(n392) );
  INV_X1 U476 ( .A(KEYINPUT106), .ZN(n391) );
  XNOR2_X2 U477 ( .A(n392), .B(n391), .ZN(n667) );
  XNOR2_X1 U478 ( .A(KEYINPUT15), .B(G902), .ZN(n590) );
  NAND2_X1 U479 ( .A1(G234), .A2(n590), .ZN(n393) );
  XNOR2_X1 U480 ( .A(KEYINPUT20), .B(n393), .ZN(n466) );
  NAND2_X1 U481 ( .A1(n466), .A2(G221), .ZN(n394) );
  XOR2_X1 U482 ( .A(n394), .B(KEYINPUT21), .Z(n646) );
  NAND2_X1 U483 ( .A1(n667), .A2(n646), .ZN(n395) );
  XNOR2_X1 U484 ( .A(n395), .B(KEYINPUT107), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n396), .B(KEYINPUT81), .ZN(n397) );
  XNOR2_X1 U486 ( .A(n398), .B(n397), .ZN(n403) );
  INV_X1 U487 ( .A(G224), .ZN(n399) );
  NOR2_X1 U488 ( .A1(n477), .A2(n399), .ZN(n401) );
  XNOR2_X1 U489 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U490 ( .A(n403), .B(n402), .ZN(n408) );
  XNOR2_X1 U491 ( .A(G110), .B(G107), .ZN(n404) );
  XNOR2_X1 U492 ( .A(n404), .B(G104), .ZN(n430) );
  XNOR2_X1 U493 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n405) );
  XNOR2_X1 U494 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U495 ( .A(n430), .B(n407), .ZN(n711) );
  XNOR2_X1 U496 ( .A(n408), .B(n711), .ZN(n410) );
  XNOR2_X1 U497 ( .A(n719), .B(G101), .ZN(n435) );
  XNOR2_X1 U498 ( .A(G113), .B(KEYINPUT3), .ZN(n409) );
  XNOR2_X1 U499 ( .A(n409), .B(G119), .ZN(n710) );
  XNOR2_X1 U500 ( .A(n435), .B(n710), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n410), .B(n450), .ZN(n603) );
  NAND2_X1 U502 ( .A1(n603), .A2(n590), .ZN(n415) );
  INV_X1 U503 ( .A(G902), .ZN(n412) );
  INV_X1 U504 ( .A(G237), .ZN(n411) );
  NAND2_X1 U505 ( .A1(n412), .A2(n411), .ZN(n416) );
  NAND2_X1 U506 ( .A1(n416), .A2(G210), .ZN(n413) );
  XNOR2_X1 U507 ( .A(n413), .B(KEYINPUT92), .ZN(n414) );
  XNOR2_X2 U508 ( .A(n415), .B(n414), .ZN(n501) );
  NAND2_X1 U509 ( .A1(n416), .A2(G214), .ZN(n497) );
  INV_X1 U510 ( .A(n497), .ZN(n664) );
  NAND2_X1 U511 ( .A1(G234), .A2(G237), .ZN(n418) );
  XNOR2_X1 U512 ( .A(n418), .B(KEYINPUT14), .ZN(n419) );
  XNOR2_X1 U513 ( .A(KEYINPUT76), .B(n419), .ZN(n420) );
  NAND2_X1 U514 ( .A1(G952), .A2(n420), .ZN(n677) );
  NOR2_X1 U515 ( .A1(n677), .A2(G953), .ZN(n481) );
  NAND2_X1 U516 ( .A1(G902), .A2(n420), .ZN(n476) );
  INV_X1 U517 ( .A(G953), .ZN(n635) );
  OR2_X1 U518 ( .A1(n635), .A2(G898), .ZN(n714) );
  NOR2_X1 U519 ( .A1(n476), .A2(n714), .ZN(n421) );
  OR2_X1 U520 ( .A1(n481), .A2(n421), .ZN(n422) );
  NAND2_X1 U521 ( .A1(n574), .A2(n422), .ZN(n424) );
  INV_X1 U522 ( .A(KEYINPUT0), .ZN(n423) );
  XNOR2_X2 U523 ( .A(n424), .B(n423), .ZN(n526) );
  NAND2_X1 U524 ( .A1(n425), .A2(n526), .ZN(n428) );
  XNOR2_X1 U525 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U526 ( .A(n426), .B(KEYINPUT65), .ZN(n427) );
  XNOR2_X1 U527 ( .A(n430), .B(n444), .ZN(n437) );
  NAND2_X1 U528 ( .A1(n722), .A2(G227), .ZN(n431) );
  XOR2_X1 U529 ( .A(G137), .B(KEYINPUT70), .Z(n459) );
  XNOR2_X1 U530 ( .A(n432), .B(n459), .ZN(n717) );
  NOR2_X2 U531 ( .A1(G902), .A2(n683), .ZN(n440) );
  XNOR2_X1 U532 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n438) );
  XNOR2_X2 U533 ( .A(n440), .B(n439), .ZN(n495) );
  XNOR2_X1 U534 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n441) );
  XNOR2_X2 U535 ( .A(n495), .B(n441), .ZN(n571) );
  XNOR2_X1 U536 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U537 ( .A(n445), .B(n444), .ZN(n452) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n448) );
  NAND2_X1 U539 ( .A1(n446), .A2(G210), .ZN(n447) );
  XNOR2_X1 U540 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U541 ( .A(n452), .B(n451), .ZN(n593) );
  NOR2_X1 U542 ( .A1(G902), .A2(n593), .ZN(n455) );
  XNOR2_X1 U543 ( .A(KEYINPUT73), .B(KEYINPUT98), .ZN(n453) );
  XOR2_X1 U544 ( .A(G140), .B(G110), .Z(n457) );
  XNOR2_X1 U545 ( .A(n457), .B(n456), .ZN(n465) );
  XNOR2_X1 U546 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U547 ( .A1(G221), .A2(n461), .ZN(n464) );
  XOR2_X1 U548 ( .A(KEYINPUT95), .B(KEYINPUT24), .Z(n463) );
  XNOR2_X1 U549 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n462) );
  XOR2_X1 U550 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n468) );
  NAND2_X1 U551 ( .A1(n466), .A2(G217), .ZN(n467) );
  XNOR2_X2 U552 ( .A(n352), .B(n365), .ZN(n647) );
  OR2_X1 U553 ( .A1(n656), .A2(n647), .ZN(n469) );
  NOR2_X1 U554 ( .A1(n571), .A2(n469), .ZN(n470) );
  NAND2_X1 U555 ( .A1(n539), .A2(n470), .ZN(n471) );
  XNOR2_X1 U556 ( .A(n471), .B(KEYINPUT108), .ZN(n521) );
  XNOR2_X1 U557 ( .A(n521), .B(G110), .ZN(G12) );
  XNOR2_X1 U558 ( .A(n501), .B(KEYINPUT38), .ZN(n556) );
  NAND2_X1 U559 ( .A1(n556), .A2(n497), .ZN(n472) );
  XNOR2_X1 U560 ( .A(n472), .B(KEYINPUT113), .ZN(n663) );
  NAND2_X1 U561 ( .A1(n663), .A2(n667), .ZN(n475) );
  INV_X1 U562 ( .A(KEYINPUT114), .ZN(n473) );
  XNOR2_X1 U563 ( .A(n473), .B(KEYINPUT41), .ZN(n474) );
  XNOR2_X1 U564 ( .A(n475), .B(n474), .ZN(n660) );
  INV_X1 U565 ( .A(n647), .ZN(n516) );
  INV_X1 U566 ( .A(n646), .ZN(n482) );
  NOR2_X1 U567 ( .A1(G900), .A2(n476), .ZN(n478) );
  NAND2_X1 U568 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U569 ( .A(KEYINPUT109), .B(n479), .ZN(n480) );
  NOR2_X1 U570 ( .A1(n481), .A2(n480), .ZN(n557) );
  NOR2_X1 U571 ( .A1(n482), .A2(n557), .ZN(n483) );
  NAND2_X1 U572 ( .A1(n516), .A2(n483), .ZN(n490) );
  INV_X1 U573 ( .A(n656), .ZN(n528) );
  NOR2_X1 U574 ( .A1(n490), .A2(n528), .ZN(n484) );
  XNOR2_X1 U575 ( .A(n484), .B(KEYINPUT28), .ZN(n485) );
  NAND2_X1 U576 ( .A1(n485), .A2(n495), .ZN(n573) );
  INV_X1 U577 ( .A(KEYINPUT42), .ZN(n486) );
  XOR2_X1 U578 ( .A(G137), .B(n565), .Z(G39) );
  XNOR2_X1 U579 ( .A(n656), .B(KEYINPUT6), .ZN(n515) );
  INV_X1 U580 ( .A(KEYINPUT105), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n504) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n561) );
  INV_X1 U583 ( .A(n561), .ZN(n624) );
  NAND2_X1 U584 ( .A1(n624), .A2(n497), .ZN(n488) );
  OR2_X1 U585 ( .A1(n504), .A2(n488), .ZN(n489) );
  NOR2_X1 U586 ( .A1(n490), .A2(n489), .ZN(n569) );
  INV_X1 U587 ( .A(n571), .ZN(n649) );
  NAND2_X1 U588 ( .A1(n569), .A2(n649), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n491), .B(KEYINPUT110), .ZN(n492) );
  XNOR2_X1 U590 ( .A(n492), .B(KEYINPUT43), .ZN(n493) );
  NAND2_X1 U591 ( .A1(n493), .A2(n501), .ZN(n585) );
  XNOR2_X1 U592 ( .A(n585), .B(G140), .ZN(G42) );
  INV_X1 U593 ( .A(n533), .ZN(n494) );
  NAND2_X1 U594 ( .A1(n494), .A2(n532), .ZN(n508) );
  INV_X1 U595 ( .A(n495), .ZN(n496) );
  NAND2_X1 U596 ( .A1(n656), .A2(n497), .ZN(n499) );
  NOR2_X1 U597 ( .A1(n508), .A2(n366), .ZN(n502) );
  INV_X1 U598 ( .A(n501), .ZN(n568) );
  NAND2_X1 U599 ( .A1(n502), .A2(n568), .ZN(n577) );
  XNOR2_X1 U600 ( .A(n577), .B(G143), .ZN(G45) );
  XNOR2_X1 U601 ( .A(n503), .B(KEYINPUT77), .ZN(n525) );
  NOR2_X1 U602 ( .A1(n525), .A2(n504), .ZN(n505) );
  XNOR2_X1 U603 ( .A(n505), .B(KEYINPUT33), .ZN(n672) );
  INV_X1 U604 ( .A(n526), .ZN(n530) );
  NOR2_X1 U605 ( .A1(n672), .A2(n530), .ZN(n507) );
  XOR2_X1 U606 ( .A(KEYINPUT34), .B(KEYINPUT83), .Z(n506) );
  XNOR2_X1 U607 ( .A(n507), .B(n506), .ZN(n510) );
  INV_X1 U608 ( .A(n508), .ZN(n509) );
  XNOR2_X1 U609 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n511) );
  NOR2_X1 U610 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n524) );
  OR2_X1 U611 ( .A1(KEYINPUT89), .A2(n524), .ZN(n513) );
  NOR2_X1 U612 ( .A1(n732), .A2(n513), .ZN(n544) );
  INV_X1 U613 ( .A(KEYINPUT44), .ZN(n522) );
  XOR2_X1 U614 ( .A(n515), .B(n514), .Z(n537) );
  NAND2_X1 U615 ( .A1(n516), .A2(n571), .ZN(n517) );
  NOR2_X1 U616 ( .A1(n537), .A2(n517), .ZN(n518) );
  XNOR2_X1 U617 ( .A(KEYINPUT84), .B(n518), .ZN(n519) );
  NAND2_X1 U618 ( .A1(n539), .A2(n519), .ZN(n520) );
  NAND2_X1 U619 ( .A1(n733), .A2(n521), .ZN(n547) );
  NOR2_X1 U620 ( .A1(n522), .A2(n547), .ZN(n523) );
  OR2_X1 U621 ( .A1(n524), .A2(n523), .ZN(n542) );
  NOR2_X1 U622 ( .A1(n525), .A2(n528), .ZN(n658) );
  NAND2_X1 U623 ( .A1(n658), .A2(n526), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n527), .B(KEYINPUT31), .ZN(n626) );
  NOR2_X1 U625 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U626 ( .A(KEYINPUT99), .B(n531), .Z(n611) );
  OR2_X1 U627 ( .A1(n626), .A2(n611), .ZN(n535) );
  NOR2_X1 U628 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U629 ( .A(KEYINPUT104), .B(n534), .ZN(n627) );
  OR2_X1 U630 ( .A1(n627), .A2(n624), .ZN(n662) );
  NAND2_X1 U631 ( .A1(n535), .A2(n662), .ZN(n540) );
  NAND2_X1 U632 ( .A1(n649), .A2(n647), .ZN(n536) );
  NOR2_X1 U633 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U634 ( .A1(n539), .A2(n538), .ZN(n609) );
  AND2_X1 U635 ( .A1(n540), .A2(n609), .ZN(n541) );
  NAND2_X1 U636 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U637 ( .A1(n544), .A2(n543), .ZN(n553) );
  NOR2_X1 U638 ( .A1(n547), .A2(KEYINPUT44), .ZN(n546) );
  INV_X1 U639 ( .A(KEYINPUT90), .ZN(n545) );
  NOR2_X1 U640 ( .A1(n546), .A2(n545), .ZN(n549) );
  NOR2_X1 U641 ( .A1(n547), .A2(KEYINPUT90), .ZN(n548) );
  NOR2_X1 U642 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U643 ( .A1(n551), .A2(n732), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X2 U645 ( .A(n555), .B(n554), .ZN(n702) );
  INV_X1 U646 ( .A(n556), .ZN(n665) );
  OR2_X1 U647 ( .A1(n665), .A2(n557), .ZN(n558) );
  XNOR2_X1 U648 ( .A(n560), .B(KEYINPUT39), .ZN(n584) );
  INV_X1 U649 ( .A(KEYINPUT112), .ZN(n562) );
  XNOR2_X1 U650 ( .A(n562), .B(KEYINPUT40), .ZN(n563) );
  NOR2_X1 U651 ( .A1(n731), .A2(n565), .ZN(n567) );
  INV_X1 U652 ( .A(KEYINPUT46), .ZN(n566) );
  XNOR2_X1 U653 ( .A(n567), .B(n566), .ZN(n581) );
  AND2_X1 U654 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U655 ( .A(n570), .B(KEYINPUT36), .ZN(n572) );
  NAND2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n630) );
  NAND2_X1 U657 ( .A1(n619), .A2(n662), .ZN(n575) );
  INV_X1 U658 ( .A(n574), .ZN(n620) );
  XNOR2_X1 U659 ( .A(n576), .B(KEYINPUT47), .ZN(n578) );
  AND2_X1 U660 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n630), .A2(n579), .ZN(n580) );
  XNOR2_X1 U662 ( .A(n582), .B(KEYINPUT48), .ZN(n587) );
  INV_X1 U663 ( .A(n627), .ZN(n583) );
  OR2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n631) );
  AND2_X1 U665 ( .A1(n585), .A2(n631), .ZN(n586) );
  XNOR2_X2 U666 ( .A(n589), .B(n588), .ZN(n638) );
  NAND2_X1 U667 ( .A1(n687), .A2(G472), .ZN(n595) );
  XOR2_X1 U668 ( .A(KEYINPUT115), .B(KEYINPUT62), .Z(n592) );
  XNOR2_X1 U669 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U670 ( .A(n595), .B(n594), .ZN(n597) );
  INV_X1 U671 ( .A(G952), .ZN(n596) );
  NOR2_X2 U672 ( .A1(n597), .A2(n701), .ZN(n599) );
  XNOR2_X1 U673 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n598) );
  XNOR2_X1 U674 ( .A(n599), .B(n598), .ZN(G57) );
  NAND2_X1 U675 ( .A1(n687), .A2(G210), .ZN(n605) );
  XNOR2_X1 U676 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n601) );
  XNOR2_X1 U677 ( .A(KEYINPUT55), .B(KEYINPUT85), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n605), .B(n604), .ZN(n606) );
  NOR2_X2 U681 ( .A1(n606), .A2(n701), .ZN(n608) );
  XNOR2_X1 U682 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n608), .B(n607), .ZN(G51) );
  XNOR2_X1 U684 ( .A(G101), .B(n609), .ZN(G3) );
  NAND2_X1 U685 ( .A1(n611), .A2(n624), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n610), .B(G104), .ZN(G6) );
  XNOR2_X1 U687 ( .A(G107), .B(KEYINPUT27), .ZN(n615) );
  XOR2_X1 U688 ( .A(KEYINPUT116), .B(KEYINPUT26), .Z(n613) );
  NAND2_X1 U689 ( .A1(n611), .A2(n627), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n615), .B(n614), .ZN(G9) );
  NAND2_X1 U692 ( .A1(n619), .A2(n627), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n616), .A2(n620), .ZN(n618) );
  XNOR2_X1 U694 ( .A(G128), .B(KEYINPUT29), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n618), .B(n617), .ZN(G30) );
  NAND2_X1 U696 ( .A1(n619), .A2(n624), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U698 ( .A(G146), .B(KEYINPUT117), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n623), .B(n622), .ZN(G48) );
  NAND2_X1 U700 ( .A1(n626), .A2(n624), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n625), .B(G113), .ZN(G15) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(G116), .ZN(G18) );
  XOR2_X1 U704 ( .A(G125), .B(KEYINPUT37), .Z(n629) );
  XNOR2_X1 U705 ( .A(n630), .B(n629), .ZN(G27) );
  INV_X1 U706 ( .A(n631), .ZN(n632) );
  XOR2_X1 U707 ( .A(G134), .B(n632), .Z(G36) );
  NOR2_X1 U708 ( .A1(n672), .A2(n660), .ZN(n634) );
  NOR2_X1 U709 ( .A1(KEYINPUT2), .A2(KEYINPUT86), .ZN(n633) );
  NOR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n645) );
  AND2_X1 U712 ( .A1(n589), .A2(KEYINPUT2), .ZN(n637) );
  NOR2_X1 U713 ( .A1(n702), .A2(n637), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n643) );
  AND2_X1 U715 ( .A1(KEYINPUT2), .A2(KEYINPUT86), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n680) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U720 ( .A(KEYINPUT49), .B(n648), .ZN(n654) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n651), .B(KEYINPUT50), .ZN(n652) );
  XNOR2_X1 U723 ( .A(KEYINPUT118), .B(n652), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT51), .B(n659), .Z(n661) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n674) );
  NAND2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n669) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n668) );
  AND2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U733 ( .A(KEYINPUT119), .B(n670), .Z(n671) );
  NOR2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U736 ( .A(KEYINPUT52), .B(n675), .ZN(n676) );
  NOR2_X1 U737 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U738 ( .A(KEYINPUT120), .B(n678), .Z(n679) );
  NAND2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U740 ( .A(KEYINPUT53), .B(n681), .Z(G75) );
  NAND2_X1 U741 ( .A1(n697), .A2(G469), .ZN(n685) );
  XOR2_X1 U742 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n682) );
  NOR2_X1 U743 ( .A1(n701), .A2(n686), .ZN(G54) );
  NAND2_X1 U744 ( .A1(n687), .A2(G475), .ZN(n690) );
  XOR2_X1 U745 ( .A(n688), .B(KEYINPUT59), .Z(n689) );
  XNOR2_X1 U746 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X2 U747 ( .A1(n691), .A2(n701), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n692), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U749 ( .A1(n697), .A2(G478), .ZN(n695) );
  NOR2_X1 U750 ( .A1(n701), .A2(n696), .ZN(G63) );
  NAND2_X1 U751 ( .A1(n697), .A2(G217), .ZN(n699) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n701), .A2(n700), .ZN(G66) );
  NOR2_X1 U754 ( .A1(n702), .A2(G953), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n703), .B(KEYINPUT123), .ZN(n707) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n704) );
  XNOR2_X1 U757 ( .A(KEYINPUT61), .B(n704), .ZN(n705) );
  NAND2_X1 U758 ( .A1(n705), .A2(G898), .ZN(n706) );
  NAND2_X1 U759 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n708), .B(KEYINPUT124), .ZN(n716) );
  XOR2_X1 U761 ( .A(G101), .B(KEYINPUT125), .Z(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U764 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U765 ( .A(n716), .B(n715), .Z(G69) );
  XNOR2_X1 U766 ( .A(n717), .B(n458), .ZN(n721) );
  XNOR2_X1 U767 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U768 ( .A(n721), .B(n720), .ZN(n724) );
  XNOR2_X1 U769 ( .A(n638), .B(n724), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n723), .A2(n722), .ZN(n730) );
  XOR2_X1 U771 ( .A(n724), .B(KEYINPUT126), .Z(n725) );
  XNOR2_X1 U772 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n727), .A2(G953), .ZN(n728) );
  XOR2_X1 U775 ( .A(KEYINPUT127), .B(n728), .Z(n729) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U777 ( .A(n731), .B(G131), .Z(G33) );
  XNOR2_X1 U778 ( .A(G122), .B(n732), .ZN(G24) );
  XNOR2_X1 U779 ( .A(G119), .B(n733), .ZN(G21) );
endmodule

