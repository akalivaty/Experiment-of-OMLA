

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(KEYINPUT91), .B(n734), .ZN(n705) );
  INV_X1 U556 ( .A(KEYINPUT97), .ZN(n761) );
  NOR2_X1 U557 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U558 ( .A1(n887), .A2(n676), .ZN(n680) );
  XOR2_X1 U559 ( .A(KEYINPUT1), .B(n534), .Z(n647) );
  XOR2_X1 U560 ( .A(KEYINPUT23), .B(n530), .Z(n523) );
  AND2_X1 U561 ( .A1(n755), .A2(n773), .ZN(n524) );
  INV_X1 U562 ( .A(KEYINPUT93), .ZN(n692) );
  XNOR2_X1 U563 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U564 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n722) );
  XNOR2_X1 U565 ( .A(n723), .B(n722), .ZN(n724) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n717) );
  NAND2_X2 U567 ( .A1(n780), .A2(n684), .ZN(n734) );
  XNOR2_X1 U568 ( .A(n762), .B(n761), .ZN(n763) );
  AND2_X1 U569 ( .A1(n681), .A2(G40), .ZN(n682) );
  NAND2_X1 U570 ( .A1(n683), .A2(n682), .ZN(n779) );
  XNOR2_X1 U571 ( .A(n560), .B(KEYINPUT14), .ZN(n561) );
  NOR2_X1 U572 ( .A1(G2104), .A2(n529), .ZN(n890) );
  INV_X1 U573 ( .A(KEYINPUT101), .ZN(n815) );
  XNOR2_X1 U574 ( .A(n562), .B(n561), .ZN(n564) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n635) );
  AND2_X1 U576 ( .A1(n529), .A2(G2104), .ZN(n886) );
  XNOR2_X1 U577 ( .A(n816), .B(n815), .ZN(n829) );
  NOR2_X1 U578 ( .A1(n643), .A2(G651), .ZN(n648) );
  XNOR2_X1 U579 ( .A(KEYINPUT17), .B(n526), .ZN(n887) );
  NOR2_X1 U580 ( .A1(n571), .A2(n570), .ZN(n1015) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X1 U582 ( .A(KEYINPUT64), .B(n525), .Z(n526) );
  NAND2_X1 U583 ( .A1(n887), .A2(G137), .ZN(n683) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NAND2_X1 U585 ( .A1(G113), .A2(n892), .ZN(n528) );
  INV_X1 U586 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U587 ( .A1(G125), .A2(n890), .ZN(n527) );
  AND2_X1 U588 ( .A1(n528), .A2(n527), .ZN(n531) );
  NAND2_X1 U589 ( .A1(G101), .A2(n886), .ZN(n530) );
  AND2_X1 U590 ( .A1(n531), .A2(n523), .ZN(n681) );
  AND2_X1 U591 ( .A1(n683), .A2(n681), .ZN(G160) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G132), .ZN(G219) );
  INV_X1 U594 ( .A(G82), .ZN(G220) );
  INV_X1 U595 ( .A(G57), .ZN(G237) );
  XOR2_X1 U596 ( .A(KEYINPUT0), .B(G543), .Z(n643) );
  XNOR2_X1 U597 ( .A(KEYINPUT65), .B(G651), .ZN(n533) );
  NOR2_X1 U598 ( .A1(n643), .A2(n533), .ZN(n633) );
  NAND2_X1 U599 ( .A1(n633), .A2(G75), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(KEYINPUT81), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n648), .A2(G50), .ZN(n536) );
  NOR2_X1 U602 ( .A1(G543), .A2(n533), .ZN(n534) );
  NAND2_X1 U603 ( .A1(G62), .A2(n647), .ZN(n535) );
  NAND2_X1 U604 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U605 ( .A(KEYINPUT80), .B(n537), .Z(n539) );
  NAND2_X1 U606 ( .A1(n635), .A2(G88), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(G166) );
  NAND2_X1 U609 ( .A1(n635), .A2(G89), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U611 ( .A1(G76), .A2(n633), .ZN(n543) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(KEYINPUT5), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n648), .A2(G51), .ZN(n547) );
  NAND2_X1 U615 ( .A1(G63), .A2(n647), .ZN(n546) );
  NAND2_X1 U616 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n548), .Z(n549) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U621 ( .A1(G138), .A2(n887), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G102), .A2(n886), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G114), .A2(n892), .ZN(n553) );
  NAND2_X1 U624 ( .A1(G126), .A2(n890), .ZN(n552) );
  AND2_X1 U625 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U626 ( .A1(n555), .A2(n554), .ZN(n677) );
  NOR2_X1 U627 ( .A1(n556), .A2(n677), .ZN(G164) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U629 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U630 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n559) );
  INV_X1 U631 ( .A(G223), .ZN(n831) );
  NAND2_X1 U632 ( .A1(G567), .A2(n831), .ZN(n558) );
  XNOR2_X1 U633 ( .A(n559), .B(n558), .ZN(G234) );
  NAND2_X1 U634 ( .A1(n647), .A2(G56), .ZN(n562) );
  INV_X1 U635 ( .A(KEYINPUT71), .ZN(n560) );
  NAND2_X1 U636 ( .A1(G43), .A2(n648), .ZN(n563) );
  NAND2_X1 U637 ( .A1(n564), .A2(n563), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n635), .A2(G81), .ZN(n565) );
  XNOR2_X1 U639 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U640 ( .A1(G68), .A2(n633), .ZN(n566) );
  NAND2_X1 U641 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U642 ( .A(KEYINPUT72), .B(n568), .Z(n569) );
  XNOR2_X1 U643 ( .A(KEYINPUT13), .B(n569), .ZN(n570) );
  NAND2_X1 U644 ( .A1(n1015), .A2(G860), .ZN(G153) );
  NAND2_X1 U645 ( .A1(n648), .A2(G52), .ZN(n573) );
  NAND2_X1 U646 ( .A1(G64), .A2(n647), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G90), .A2(n635), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G77), .A2(n633), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U651 ( .A(KEYINPUT9), .B(n576), .Z(n577) );
  NOR2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U653 ( .A(KEYINPUT68), .B(n579), .ZN(G171) );
  XNOR2_X1 U654 ( .A(KEYINPUT73), .B(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n635), .A2(G92), .ZN(n581) );
  NAND2_X1 U657 ( .A1(G66), .A2(n647), .ZN(n580) );
  NAND2_X1 U658 ( .A1(n581), .A2(n580), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G79), .A2(n633), .ZN(n582) );
  XNOR2_X1 U660 ( .A(n582), .B(KEYINPUT74), .ZN(n584) );
  NAND2_X1 U661 ( .A1(G54), .A2(n648), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U663 ( .A(KEYINPUT75), .B(n585), .Z(n586) );
  NOR2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U665 ( .A(KEYINPUT15), .B(n588), .Z(n857) );
  INV_X1 U666 ( .A(n857), .ZN(n1006) );
  INV_X1 U667 ( .A(G868), .ZN(n658) );
  NAND2_X1 U668 ( .A1(n1006), .A2(n658), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U670 ( .A1(n648), .A2(G53), .ZN(n592) );
  NAND2_X1 U671 ( .A1(G65), .A2(n647), .ZN(n591) );
  NAND2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U673 ( .A(KEYINPUT69), .B(n593), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n633), .A2(G78), .ZN(n595) );
  NAND2_X1 U675 ( .A1(G91), .A2(n635), .ZN(n594) );
  AND2_X1 U676 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U678 ( .A1(G286), .A2(n658), .ZN(n599) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U680 ( .A1(n599), .A2(n598), .ZN(G297) );
  INV_X1 U681 ( .A(G860), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n601), .A2(n857), .ZN(n602) );
  XNOR2_X1 U684 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U685 ( .A1(n857), .A2(G868), .ZN(n603) );
  NOR2_X1 U686 ( .A1(G559), .A2(n603), .ZN(n605) );
  AND2_X1 U687 ( .A1(n658), .A2(n1015), .ZN(n604) );
  NOR2_X1 U688 ( .A1(n605), .A2(n604), .ZN(G282) );
  XOR2_X1 U689 ( .A(G2100), .B(KEYINPUT78), .Z(n616) );
  NAND2_X1 U690 ( .A1(G123), .A2(n890), .ZN(n606) );
  XNOR2_X1 U691 ( .A(n606), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U692 ( .A1(G99), .A2(n886), .ZN(n608) );
  NAND2_X1 U693 ( .A1(G135), .A2(n887), .ZN(n607) );
  NAND2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n892), .A2(G111), .ZN(n609) );
  XOR2_X1 U696 ( .A(KEYINPUT76), .B(n609), .Z(n610) );
  NOR2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n940) );
  XNOR2_X1 U699 ( .A(KEYINPUT77), .B(n940), .ZN(n614) );
  XNOR2_X1 U700 ( .A(n614), .B(G2096), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U702 ( .A1(G559), .A2(n857), .ZN(n617) );
  XOR2_X1 U703 ( .A(n1015), .B(n617), .Z(n656) );
  NOR2_X1 U704 ( .A1(n656), .A2(G860), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n648), .A2(G55), .ZN(n619) );
  NAND2_X1 U706 ( .A1(G67), .A2(n647), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U708 ( .A1(G93), .A2(n635), .ZN(n621) );
  NAND2_X1 U709 ( .A1(G80), .A2(n633), .ZN(n620) );
  NAND2_X1 U710 ( .A1(n621), .A2(n620), .ZN(n622) );
  OR2_X1 U711 ( .A1(n623), .A2(n622), .ZN(n659) );
  XOR2_X1 U712 ( .A(n624), .B(n659), .Z(G145) );
  NAND2_X1 U713 ( .A1(G47), .A2(n648), .ZN(n625) );
  XNOR2_X1 U714 ( .A(n625), .B(KEYINPUT66), .ZN(n627) );
  NAND2_X1 U715 ( .A1(G60), .A2(n647), .ZN(n626) );
  NAND2_X1 U716 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U717 ( .A1(G85), .A2(n635), .ZN(n629) );
  NAND2_X1 U718 ( .A1(G72), .A2(n633), .ZN(n628) );
  NAND2_X1 U719 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U720 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U721 ( .A(KEYINPUT67), .B(n632), .ZN(G290) );
  NAND2_X1 U722 ( .A1(n633), .A2(G73), .ZN(n634) );
  XNOR2_X1 U723 ( .A(n634), .B(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n635), .A2(G86), .ZN(n637) );
  NAND2_X1 U725 ( .A1(G61), .A2(n647), .ZN(n636) );
  NAND2_X1 U726 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U727 ( .A1(G48), .A2(n648), .ZN(n638) );
  XNOR2_X1 U728 ( .A(KEYINPUT79), .B(n638), .ZN(n639) );
  NOR2_X1 U729 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U732 ( .A1(G87), .A2(n643), .ZN(n644) );
  NAND2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U734 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n648), .A2(G49), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G288) );
  INV_X1 U737 ( .A(G299), .ZN(n1001) );
  XNOR2_X1 U738 ( .A(G166), .B(n1001), .ZN(n655) );
  XNOR2_X1 U739 ( .A(G290), .B(G305), .ZN(n653) );
  XOR2_X1 U740 ( .A(KEYINPUT19), .B(n659), .Z(n651) );
  XNOR2_X1 U741 ( .A(n651), .B(G288), .ZN(n652) );
  XNOR2_X1 U742 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U743 ( .A(n655), .B(n654), .ZN(n860) );
  XNOR2_X1 U744 ( .A(n656), .B(n860), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U747 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U752 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G120), .A2(G69), .ZN(n666) );
  NOR2_X1 U755 ( .A1(G237), .A2(n666), .ZN(n667) );
  XNOR2_X1 U756 ( .A(KEYINPUT82), .B(n667), .ZN(n668) );
  NAND2_X1 U757 ( .A1(n668), .A2(G108), .ZN(n835) );
  NAND2_X1 U758 ( .A1(n835), .A2(G567), .ZN(n673) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U761 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U762 ( .A1(G96), .A2(n671), .ZN(n836) );
  NAND2_X1 U763 ( .A1(n836), .A2(G2106), .ZN(n672) );
  NAND2_X1 U764 ( .A1(n673), .A2(n672), .ZN(n837) );
  NAND2_X1 U765 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U766 ( .A1(n837), .A2(n674), .ZN(n834) );
  NAND2_X1 U767 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U768 ( .A(G166), .ZN(G303) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n675) );
  XNOR2_X1 U770 ( .A(n675), .B(KEYINPUT24), .ZN(n686) );
  INV_X1 U771 ( .A(G1384), .ZN(n678) );
  AND2_X1 U772 ( .A1(G138), .A2(n678), .ZN(n676) );
  AND2_X1 U773 ( .A1(n678), .A2(n677), .ZN(n679) );
  OR2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n780) );
  INV_X1 U775 ( .A(n779), .ZN(n684) );
  NAND2_X1 U776 ( .A1(n734), .A2(G8), .ZN(n685) );
  XNOR2_X1 U777 ( .A(n685), .B(KEYINPUT88), .ZN(n688) );
  BUF_X1 U778 ( .A(n688), .Z(n773) );
  INV_X1 U779 ( .A(n773), .ZN(n764) );
  NAND2_X1 U780 ( .A1(n686), .A2(n764), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n687), .B(KEYINPUT89), .ZN(n757) );
  NOR2_X1 U782 ( .A1(n688), .A2(G1966), .ZN(n730) );
  XNOR2_X1 U783 ( .A(G2078), .B(KEYINPUT25), .ZN(n952) );
  NAND2_X1 U784 ( .A1(n705), .A2(n952), .ZN(n690) );
  XOR2_X1 U785 ( .A(KEYINPUT90), .B(G1961), .Z(n989) );
  NAND2_X1 U786 ( .A1(n989), .A2(n734), .ZN(n689) );
  NAND2_X1 U787 ( .A1(n690), .A2(n689), .ZN(n725) );
  NAND2_X1 U788 ( .A1(n725), .A2(G171), .ZN(n720) );
  NAND2_X1 U789 ( .A1(n705), .A2(G2072), .ZN(n691) );
  XNOR2_X1 U790 ( .A(KEYINPUT27), .B(n691), .ZN(n695) );
  XOR2_X1 U791 ( .A(KEYINPUT92), .B(G1956), .Z(n976) );
  NOR2_X1 U792 ( .A1(n705), .A2(n976), .ZN(n693) );
  NOR2_X1 U793 ( .A1(n695), .A2(n694), .ZN(n697) );
  NOR2_X1 U794 ( .A1(n697), .A2(n1001), .ZN(n696) );
  XOR2_X1 U795 ( .A(n696), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U796 ( .A1(n697), .A2(n1001), .ZN(n714) );
  NAND2_X1 U797 ( .A1(n734), .A2(G1341), .ZN(n698) );
  XNOR2_X1 U798 ( .A(n698), .B(KEYINPUT94), .ZN(n699) );
  NAND2_X1 U799 ( .A1(n699), .A2(n1015), .ZN(n703) );
  INV_X1 U800 ( .A(n734), .ZN(n700) );
  NAND2_X1 U801 ( .A1(G1996), .A2(n700), .ZN(n701) );
  XOR2_X1 U802 ( .A(KEYINPUT26), .B(n701), .Z(n702) );
  NOR2_X1 U803 ( .A1(n703), .A2(n702), .ZN(n704) );
  OR2_X1 U804 ( .A1(n857), .A2(n704), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n857), .A2(n704), .ZN(n710) );
  NAND2_X1 U806 ( .A1(G2067), .A2(n705), .ZN(n707) );
  NAND2_X1 U807 ( .A1(G1348), .A2(n734), .ZN(n706) );
  NAND2_X1 U808 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U809 ( .A(KEYINPUT95), .B(n708), .Z(n709) );
  NAND2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U813 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U814 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n741) );
  NOR2_X1 U816 ( .A1(G2084), .A2(n734), .ZN(n731) );
  NOR2_X1 U817 ( .A1(n730), .A2(n731), .ZN(n721) );
  NAND2_X1 U818 ( .A1(G8), .A2(n721), .ZN(n723) );
  NOR2_X1 U819 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U820 ( .A1(n725), .A2(G171), .ZN(n726) );
  NOR2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U822 ( .A(n728), .B(KEYINPUT31), .Z(n740) );
  AND2_X1 U823 ( .A1(n741), .A2(n740), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U825 ( .A1(G8), .A2(n731), .ZN(n732) );
  NAND2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n750) );
  INV_X1 U827 ( .A(G8), .ZN(n739) );
  NOR2_X1 U828 ( .A1(n773), .A2(G1971), .ZN(n736) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U831 ( .A1(n737), .A2(G303), .ZN(n738) );
  OR2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n743) );
  AND2_X1 U833 ( .A1(n740), .A2(n743), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n747) );
  INV_X1 U835 ( .A(n743), .ZN(n745) );
  AND2_X1 U836 ( .A1(G286), .A2(G8), .ZN(n744) );
  OR2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U839 ( .A(n748), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n760) );
  INV_X1 U841 ( .A(n760), .ZN(n753) );
  NAND2_X1 U842 ( .A1(G8), .A2(G166), .ZN(n751) );
  NOR2_X1 U843 ( .A1(G2090), .A2(n751), .ZN(n752) );
  XNOR2_X1 U844 ( .A(n754), .B(KEYINPUT99), .ZN(n755) );
  XNOR2_X1 U845 ( .A(n524), .B(KEYINPUT100), .ZN(n756) );
  NOR2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n778) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n1007) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n769) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U850 ( .A1(n769), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(KEYINPUT98), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n1019) );
  NAND2_X1 U854 ( .A1(n1019), .A2(n764), .ZN(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U856 ( .A1(KEYINPUT33), .A2(n767), .ZN(n775) );
  NAND2_X1 U857 ( .A1(KEYINPUT33), .A2(KEYINPUT98), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n771) );
  INV_X1 U859 ( .A(n769), .ZN(n1018) );
  NAND2_X1 U860 ( .A1(KEYINPUT98), .A2(n1018), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n1007), .A2(n776), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n814) );
  NOR2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n826) );
  XNOR2_X1 U867 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NAND2_X1 U868 ( .A1(G104), .A2(n886), .ZN(n782) );
  NAND2_X1 U869 ( .A1(G140), .A2(n887), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n783), .ZN(n789) );
  NAND2_X1 U872 ( .A1(G116), .A2(n892), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G128), .A2(n890), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U875 ( .A(KEYINPUT35), .B(n786), .ZN(n787) );
  XNOR2_X1 U876 ( .A(KEYINPUT83), .B(n787), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U878 ( .A(KEYINPUT36), .B(n790), .ZN(n904) );
  NOR2_X1 U879 ( .A1(n824), .A2(n904), .ZN(n942) );
  NAND2_X1 U880 ( .A1(n826), .A2(n942), .ZN(n822) );
  NAND2_X1 U881 ( .A1(n886), .A2(G95), .ZN(n791) );
  XNOR2_X1 U882 ( .A(n791), .B(KEYINPUT84), .ZN(n793) );
  NAND2_X1 U883 ( .A1(G107), .A2(n892), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n890), .A2(G119), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G131), .A2(n887), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n796) );
  OR2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n899) );
  AND2_X1 U889 ( .A1(n899), .A2(G1991), .ZN(n808) );
  NAND2_X1 U890 ( .A1(n892), .A2(G117), .ZN(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT85), .B(n798), .Z(n800) );
  NAND2_X1 U892 ( .A1(n890), .A2(G129), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U894 ( .A(KEYINPUT86), .B(n801), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n886), .A2(G105), .ZN(n802) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(n802), .Z(n803) );
  NOR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U898 ( .A1(G141), .A2(n887), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n873) );
  AND2_X1 U900 ( .A1(n873), .A2(G1996), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n925) );
  INV_X1 U902 ( .A(n826), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n925), .A2(n809), .ZN(n819) );
  XNOR2_X1 U904 ( .A(KEYINPUT87), .B(n819), .ZN(n811) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n1005) );
  NAND2_X1 U906 ( .A1(n826), .A2(n1005), .ZN(n810) );
  AND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U908 ( .A1(n822), .A2(n812), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n816) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n873), .ZN(n932) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n899), .ZN(n939) );
  NOR2_X1 U913 ( .A1(n817), .A2(n939), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n932), .A2(n820), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n824), .A2(n904), .ZN(n924) );
  NAND2_X1 U919 ( .A1(n825), .A2(n924), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U922 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U925 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n837), .ZN(G319) );
  XOR2_X1 U936 ( .A(G2678), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT104), .B(KEYINPUT103), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2090), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2100), .B(G2096), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U945 ( .A(G2078), .B(G2084), .Z(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1971), .B(G1976), .Z(n849) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1981), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n850), .B(G2474), .Z(n852) );
  XNOR2_X1 U951 ( .A(G1966), .B(G1956), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT41), .B(G1961), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(G229) );
  XNOR2_X1 U957 ( .A(n1015), .B(G286), .ZN(n859) );
  XNOR2_X1 U958 ( .A(G171), .B(n857), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  NOR2_X1 U961 ( .A1(G37), .A2(n862), .ZN(G397) );
  NAND2_X1 U962 ( .A1(n887), .A2(G136), .ZN(n871) );
  NAND2_X1 U963 ( .A1(G124), .A2(n890), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n863), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G100), .A2(n886), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n864), .B(KEYINPUT106), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G112), .A2(n892), .ZN(n867) );
  XNOR2_X1 U969 ( .A(KEYINPUT105), .B(n867), .ZN(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT107), .ZN(G162) );
  XOR2_X1 U973 ( .A(n873), .B(G162), .Z(n903) );
  NAND2_X1 U974 ( .A1(G106), .A2(n886), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G142), .A2(n887), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT45), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G118), .A2(n892), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G130), .A2(n890), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(KEYINPUT108), .B(n879), .Z(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n882), .B(G164), .ZN(n883) );
  XNOR2_X1 U984 ( .A(KEYINPUT48), .B(n883), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n940), .B(KEYINPUT46), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n898) );
  NAND2_X1 U987 ( .A1(G103), .A2(n886), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G139), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n897) );
  NAND2_X1 U990 ( .A1(n890), .A2(G127), .ZN(n891) );
  XOR2_X1 U991 ( .A(KEYINPUT109), .B(n891), .Z(n894) );
  NAND2_X1 U992 ( .A1(n892), .A2(G115), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n926) );
  XOR2_X1 U996 ( .A(n898), .B(n926), .Z(n901) );
  XOR2_X1 U997 ( .A(G160), .B(n899), .Z(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n906), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT110), .B(n907), .ZN(G395) );
  XOR2_X1 U1003 ( .A(G2438), .B(G2435), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G2443), .B(G2430), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n910), .B(G2454), .Z(n912) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1009 ( .A(G2451), .B(G2427), .Z(n914) );
  XNOR2_X1 U1010 ( .A(KEYINPUT102), .B(G2446), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1012 ( .A(n916), .B(n915), .Z(n917) );
  NAND2_X1 U1013 ( .A1(G14), .A2(n917), .ZN(n923) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G397), .A2(G395), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(n923), .ZN(G401) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n937) );
  XOR2_X1 U1023 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT112), .B(n929), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n930), .B(KEYINPUT50), .ZN(n935) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n946) );
  XOR2_X1 U1033 ( .A(G160), .B(G2084), .Z(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT111), .B(n944), .Z(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(n947), .B(KEYINPUT52), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n948), .A2(G29), .ZN(n972) );
  XNOR2_X1 U1041 ( .A(G1991), .B(G25), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n957) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n951) );
  NAND2_X1 U1045 ( .A1(n951), .A2(G28), .ZN(n955) );
  XOR2_X1 U1046 ( .A(G27), .B(n952), .Z(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT114), .B(n953), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1050 ( .A(KEYINPUT115), .B(G1996), .Z(n958) );
  XNOR2_X1 U1051 ( .A(G32), .B(n958), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1053 ( .A(KEYINPUT53), .B(n961), .Z(n964) );
  XOR2_X1 U1054 ( .A(G34), .B(KEYINPUT54), .Z(n962) );
  XNOR2_X1 U1055 ( .A(G2084), .B(n962), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(n967), .B(KEYINPUT116), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n968), .ZN(n969) );
  XOR2_X1 U1061 ( .A(n969), .B(KEYINPUT55), .Z(n970) );
  XNOR2_X1 U1062 ( .A(KEYINPUT113), .B(n970), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n1033) );
  XOR2_X1 U1064 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n974) );
  XNOR2_X1 U1065 ( .A(KEYINPUT59), .B(G4), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1067 ( .A(G1348), .B(n975), .Z(n983) );
  XOR2_X1 U1068 ( .A(G1981), .B(G6), .Z(n978) );
  XNOR2_X1 U1069 ( .A(n976), .B(G20), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G19), .B(G1341), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1075 ( .A(n984), .B(KEYINPUT60), .Z(n985) );
  XNOR2_X1 U1076 ( .A(KEYINPUT124), .B(n985), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(G21), .B(G1966), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT125), .B(n988), .Z(n991) );
  XNOR2_X1 U1080 ( .A(n989), .B(G5), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n998) );
  XNOR2_X1 U1082 ( .A(G1976), .B(G23), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1971), .B(G22), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1085 ( .A(G1986), .B(G24), .Z(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT58), .B(n996), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1089 ( .A(KEYINPUT61), .B(n999), .Z(n1000) );
  NOR2_X1 U1090 ( .A1(G16), .A2(n1000), .ZN(n1030) );
  XOR2_X1 U1091 ( .A(G16), .B(KEYINPUT56), .Z(n1027) );
  XNOR2_X1 U1092 ( .A(n1001), .B(G1956), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(G171), .B(G1961), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1014) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G1348), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G168), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(KEYINPUT117), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT57), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1025) );
  XOR2_X1 U1103 ( .A(n1015), .B(G1341), .Z(n1017) );
  XOR2_X1 U1104 ( .A(G1971), .B(G166), .Z(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(n1018), .B(KEYINPUT118), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1021), .B(KEYINPUT119), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(n1028), .B(KEYINPUT120), .ZN(n1029) );
  NOR2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1114 ( .A(KEYINPUT126), .B(n1031), .Z(n1032) );
  NOR2_X1 U1115 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1116 ( .A1(n1034), .A2(G11), .ZN(n1035) );
  XNOR2_X1 U1117 ( .A(n1035), .B(KEYINPUT127), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1036), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

