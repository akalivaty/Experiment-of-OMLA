//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n596, new_n597, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT67), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n454), .B2(G2106), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT71), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n463), .B2(new_n465), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT71), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n461), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n462), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT72), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n483), .A3(G101), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n479), .A2(G2105), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n473), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n467), .B1(new_n463), .B2(new_n465), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(G124), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n471), .A2(G136), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND2_X1  g070(.A1(new_n480), .A2(G102), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n466), .B2(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n496), .B1(new_n499), .B2(new_n467), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n467), .A2(G138), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT3), .B1(new_n464), .B2(G2104), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n463), .B2(new_n465), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n509), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n500), .B1(new_n510), .B2(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n515), .B1(new_n521), .B2(new_n523), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT74), .B(G651), .Z(new_n528));
  INV_X1    g103(.A(new_n517), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(G62), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n531), .A2(new_n532), .B1(G75), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G62), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n516), .B2(new_n517), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT75), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n528), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n525), .B(new_n527), .C1(new_n537), .C2(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n533), .A2(new_n536), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(new_n520), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT77), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n541), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n546));
  AOI22_X1  g121(.A1(G88), .A2(new_n524), .B1(new_n526), .B2(G50), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(G166));
  NAND2_X1  g124(.A1(new_n526), .A2(G51), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n553));
  AND2_X1   g128(.A1(G63), .A2(G651), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n552), .A2(new_n553), .B1(new_n518), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n524), .A2(G89), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(G286));
  INV_X1    g133(.A(G286), .ZN(G168));
  AOI22_X1  g134(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n528), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT78), .ZN(new_n562));
  AOI22_X1  g137(.A1(G90), .A2(new_n524), .B1(new_n526), .B2(G52), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G171));
  NAND2_X1  g140(.A1(G68), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G56), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n519), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n526), .A2(G43), .B1(new_n568), .B2(new_n520), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n524), .A2(G81), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT79), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT80), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND4_X1  g153(.A1(G319), .A2(G483), .A3(G661), .A4(new_n578), .ZN(G188));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n526), .B2(G53), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n526), .A2(new_n581), .A3(G53), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G65), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n519), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n524), .A2(G91), .B1(new_n588), .B2(G651), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n580), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n584), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n580), .B(new_n589), .C1(new_n591), .C2(new_n582), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(G299));
  NAND2_X1  g169(.A1(new_n564), .A2(KEYINPUT82), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n564), .A2(KEYINPUT82), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(G301));
  INV_X1    g173(.A(G166), .ZN(G303));
  NAND2_X1  g174(.A1(new_n524), .A2(G87), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n526), .A2(G49), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G288));
  NAND2_X1  g178(.A1(new_n524), .A2(G86), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n526), .A2(G48), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n528), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(G72), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G60), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n519), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n528), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(new_n611), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n524), .A2(G85), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n526), .A2(G47), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n617), .A2(KEYINPUT84), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n617), .A2(KEYINPUT84), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(new_n524), .A2(G92), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT10), .Z(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  INV_X1    g198(.A(G66), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n519), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n526), .A2(G54), .B1(new_n625), .B2(G651), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  MUX2_X1   g202(.A(new_n627), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g203(.A(new_n627), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(new_n627), .ZN(new_n634));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G860), .ZN(G148));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n571), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n638), .B1(new_n640), .B2(new_n637), .ZN(G323));
  XOR2_X1   g216(.A(G323), .B(KEYINPUT85), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g218(.A1(new_n475), .A2(new_n476), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n480), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT13), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n471), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n491), .A2(G123), .ZN(new_n651));
  NOR2_X1   g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n656), .ZN(G156));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT88), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT87), .B(KEYINPUT16), .Z(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2072), .B(G2078), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(KEYINPUT89), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n682));
  OAI22_X1  g257(.A1(new_n681), .A2(new_n682), .B1(new_n676), .B2(new_n677), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  OAI221_X1 g259(.A(new_n678), .B1(new_n677), .B2(new_n680), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n676), .A2(new_n679), .A3(new_n677), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT18), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(new_n655), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2100), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT90), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1961), .B(G1966), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT20), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n694), .B(new_n695), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n698), .B(new_n699), .C1(new_n693), .C2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1986), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT91), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1981), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n704), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G4), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n634), .B2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(G21), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G168), .B2(new_n713), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT100), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n717), .B1(new_n720), .B2(G1966), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G33), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n644), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI21_X1  g299(.A(G2105), .B1(new_n724), .B2(KEYINPUT98), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(KEYINPUT98), .B2(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT25), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n471), .A2(G139), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n723), .B1(new_n731), .B2(new_n722), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n722), .A2(G35), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G162), .B2(new_n722), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT29), .B(G2090), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT24), .B(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(new_n722), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT99), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n486), .B2(new_n722), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n732), .A2(G2072), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n733), .A2(new_n737), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G171), .A2(new_n713), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G5), .B2(new_n713), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n572), .A2(new_n713), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n713), .B2(G19), .ZN(new_n751));
  INV_X1    g326(.A(G1341), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(new_n742), .B2(new_n741), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n747), .A2(new_n748), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n749), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n721), .A2(new_n745), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(KEYINPUT30), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n654), .B2(new_n722), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n722), .A2(G26), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT28), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n471), .A2(G140), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n491), .A2(G128), .ZN(new_n767));
  NOR2_X1   g342(.A1(G104), .A2(G2105), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT97), .B(G2067), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n763), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n751), .B2(new_n752), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT26), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(G105), .B2(new_n480), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n471), .A2(G141), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n491), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G32), .B(new_n783), .S(G29), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT27), .B(G1996), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n722), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n722), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2078), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n774), .A2(new_n775), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n720), .A2(G1966), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT101), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n713), .A2(G20), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT23), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n631), .B2(new_n713), .ZN(new_n795));
  INV_X1    g370(.A(G1956), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n756), .A2(new_n790), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G24), .ZN(new_n799));
  INV_X1    g374(.A(G290), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n801), .A2(G1986), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n722), .A2(G25), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT92), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n471), .A2(G131), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n491), .A2(G119), .ZN(new_n806));
  OR2_X1    g381(.A1(G95), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT93), .Z(new_n810));
  OAI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(new_n722), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n801), .A2(G1986), .ZN(new_n815));
  OR3_X1    g390(.A1(new_n802), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n713), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n713), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT33), .B(G1976), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n713), .A2(G6), .ZN(new_n822));
  INV_X1    g397(.A(G305), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n713), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT32), .B(G1981), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n826), .A2(new_n827), .ZN(new_n832));
  INV_X1    g407(.A(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n821), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(G16), .A2(G22), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G166), .B2(G16), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT96), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(KEYINPUT96), .ZN(new_n840));
  INV_X1    g415(.A(G1971), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n839), .B2(new_n840), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n835), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n816), .B1(new_n844), .B2(KEYINPUT34), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT34), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n835), .A2(new_n846), .A3(new_n842), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT36), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT36), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n798), .B1(new_n849), .B2(new_n851), .ZN(G311));
  INV_X1    g427(.A(new_n798), .ZN(new_n853));
  INV_X1    g428(.A(new_n851), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n850), .B1(new_n845), .B2(new_n847), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(G150));
  NAND2_X1  g431(.A1(new_n524), .A2(G93), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n526), .A2(G55), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n857), .B(new_n858), .C1(new_n528), .C2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n571), .B(new_n860), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n634), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT102), .B(G860), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(G145));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT4), .B1(new_n508), .B2(KEYINPUT73), .ZN(new_n874));
  AOI211_X1 g449(.A(new_n506), .B(new_n501), .C1(new_n463), .C2(new_n465), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n512), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n496), .ZN(new_n877));
  OAI21_X1  g452(.A(G126), .B1(new_n503), .B2(new_n504), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n497), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n879), .B2(G2105), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n885));
  NOR2_X1   g460(.A1(G106), .A2(G2105), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n491), .B2(G130), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n471), .A2(G142), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n809), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n809), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n645), .B(new_n646), .Z(new_n894));
  NOR3_X1   g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n806), .A2(new_n808), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n896), .A2(new_n805), .A3(new_n889), .A4(new_n888), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n647), .B1(new_n897), .B2(new_n891), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n882), .B(new_n884), .C1(new_n895), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n770), .B(new_n783), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n647), .A3(new_n891), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n894), .B1(new_n892), .B2(new_n893), .ZN(new_n903));
  INV_X1    g478(.A(new_n882), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(new_n883), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n899), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n901), .B1(new_n899), .B2(new_n905), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n906), .A2(new_n907), .B1(new_n726), .B2(new_n730), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n899), .A2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n900), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n899), .A2(new_n901), .A3(new_n905), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n731), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G160), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n494), .B(new_n654), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n908), .A2(new_n912), .A3(new_n913), .A4(new_n486), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n873), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n915), .A2(new_n917), .ZN(new_n923));
  INV_X1    g498(.A(new_n916), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(KEYINPUT105), .A3(new_n919), .A4(new_n918), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n922), .A2(KEYINPUT40), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT40), .B1(new_n922), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(G395));
  NAND2_X1  g504(.A1(G290), .A2(G288), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n818), .B(new_n614), .C1(new_n618), .C2(new_n619), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  NOR2_X1   g508(.A1(G303), .A2(G305), .ZN(new_n934));
  NOR2_X1   g509(.A1(G166), .A2(new_n823), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n935), .B2(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OR3_X1    g516(.A1(new_n941), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n942));
  NOR2_X1   g517(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT107), .B1(new_n590), .B2(new_n593), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n589), .B1(new_n591), .B2(new_n582), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT81), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n592), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n634), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(G299), .A2(new_n951), .A3(new_n627), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT41), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(KEYINPUT41), .A3(new_n954), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n861), .B(KEYINPUT106), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(new_n640), .ZN(new_n962));
  MUX2_X1   g537(.A(new_n956), .B(new_n960), .S(new_n962), .Z(new_n963));
  AND2_X1   g538(.A1(new_n947), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n947), .A2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n860), .A2(new_n637), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  INV_X1    g544(.A(KEYINPUT82), .ZN(new_n970));
  NAND2_X1  g545(.A1(G171), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G286), .B1(new_n971), .B2(new_n595), .ZN(new_n972));
  NOR2_X1   g547(.A1(G171), .A2(G168), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n861), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n861), .ZN(new_n975));
  INV_X1    g550(.A(new_n973), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n975), .B(new_n976), .C1(G301), .C2(G286), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n958), .A2(new_n959), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n977), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n956), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n941), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n978), .A2(new_n980), .A3(new_n938), .A4(new_n940), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT44), .B1(new_n986), .B2(KEYINPUT110), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(G397));
  OR2_X1    g568(.A1(G290), .A2(G1986), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT112), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT111), .B(G1384), .Z(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(G164), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n473), .A2(G40), .A3(new_n485), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  INV_X1    g580(.A(G2067), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n770), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n783), .B(G1996), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n809), .B(new_n812), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n1000), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1004), .A2(new_n1005), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n810), .A2(new_n812), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1010), .A3(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n770), .A2(G2067), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1001), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n1001), .A2(new_n1021), .A3(G1996), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1000), .B1(new_n783), .B2(new_n1008), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1001), .B2(G1996), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1020), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1014), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n473), .A2(G40), .A3(new_n485), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n876), .B2(new_n880), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n604), .A2(new_n605), .A3(new_n607), .A4(new_n1035), .ZN(new_n1036));
  OR2_X1    g611(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1034), .A2(KEYINPUT116), .A3(KEYINPUT49), .A4(new_n1036), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1033), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n818), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1036), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1033), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1031), .B1(new_n1032), .B2(KEYINPUT45), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n996), .B(new_n997), .C1(new_n876), .C2(new_n880), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n996), .B1(G164), .B2(G1384), .ZN(new_n1051));
  INV_X1    g626(.A(new_n997), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n881), .A2(KEYINPUT45), .A3(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1051), .A2(KEYINPUT113), .A3(new_n1031), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n841), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1384), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT4), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n505), .B2(new_n506), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n511), .B1(new_n1058), .B2(new_n509), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1059), .B2(new_n500), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n999), .B1(new_n1060), .B2(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1032), .A2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT114), .B(G2090), .Z(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1030), .B1(new_n1055), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n543), .A2(G8), .A3(new_n548), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n600), .A2(new_n601), .A3(G1976), .A4(new_n602), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT115), .ZN(new_n1072));
  OAI21_X1  g647(.A(G8), .B1(new_n1060), .B2(new_n999), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT52), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1071), .A2(KEYINPUT115), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(KEYINPUT115), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1033), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1042), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1046), .B1(new_n1070), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1067), .B(KEYINPUT55), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1063), .A2(KEYINPUT117), .ZN(new_n1082));
  AOI211_X1 g657(.A(KEYINPUT50), .B(G1384), .C1(new_n876), .C2(new_n880), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(new_n1061), .A4(new_n1064), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1055), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1081), .B1(new_n1087), .B2(new_n1030), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1079), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1089));
  INV_X1    g664(.A(G1966), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n996), .B(G1384), .C1(new_n876), .C2(new_n880), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n1048), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1060), .A2(KEYINPUT50), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(new_n742), .A3(new_n1063), .A4(new_n1031), .ZN(new_n1094));
  AOI211_X1 g669(.A(new_n1030), .B(G286), .C1(new_n1092), .C2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1095), .A2(KEYINPUT63), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1089), .B(new_n1099), .C1(new_n1069), .C2(new_n1066), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1080), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1092), .A2(new_n1094), .A3(G168), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT51), .ZN(new_n1104));
  AOI21_X1  g679(.A(G168), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  OAI211_X1 g681(.A(G8), .B(new_n1102), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1031), .B1(new_n1032), .B2(new_n1062), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n748), .B1(new_n1110), .B2(new_n1083), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1032), .A2(KEYINPUT45), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G2078), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1051), .A2(new_n1112), .A3(new_n1031), .A4(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1111), .A2(KEYINPUT122), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT122), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G2078), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n999), .B1(new_n1060), .B2(new_n996), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT113), .B1(new_n1120), .B2(new_n1053), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1048), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1113), .ZN(new_n1124));
  AOI21_X1  g699(.A(G301), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1109), .A2(new_n1125), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1126), .A2(KEYINPUT126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1104), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1107), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT62), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1126), .B2(KEYINPUT126), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1101), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1082), .A2(new_n1085), .A3(new_n1061), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n796), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n949), .B(KEYINPUT57), .Z(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1120), .A2(new_n1053), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1060), .A2(new_n999), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1139), .A2(new_n716), .B1(new_n1006), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n627), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT119), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1135), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1138), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1138), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1147), .B2(new_n1144), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1144), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT61), .A3(new_n1138), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1048), .A2(G1996), .A3(new_n1049), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT58), .B(G1341), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1140), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n572), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1148), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n634), .B1(new_n1141), .B2(KEYINPUT60), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT121), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1162), .B(new_n634), .C1(new_n1141), .C2(KEYINPUT60), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1158), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1145), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1088), .B(new_n1089), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(G301), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1118), .A2(new_n1124), .A3(new_n1171), .A4(G301), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT53), .B1(new_n1119), .B2(KEYINPUT123), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(KEYINPUT123), .B2(new_n1119), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1053), .A2(new_n1031), .A3(new_n1176), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n748), .A2(new_n1139), .B1(new_n1177), .B2(new_n998), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1124), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1174), .B1(new_n1179), .B2(new_n564), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT54), .B1(new_n1173), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1124), .A2(G301), .A3(new_n1178), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1182), .A2(KEYINPUT124), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1125), .A2(KEYINPUT54), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(KEYINPUT124), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1170), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1132), .B1(new_n1169), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1012), .B1(G1986), .B2(G290), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1001), .B1(new_n995), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1029), .B1(new_n1188), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g766(.A1(new_n922), .A2(new_n926), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n674), .A2(G319), .ZN(new_n1194));
  NOR4_X1   g768(.A1(new_n709), .A2(new_n710), .A3(G227), .A4(new_n1194), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1193), .A2(new_n988), .A3(new_n1195), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


