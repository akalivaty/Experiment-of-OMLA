

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775;

  XNOR2_X1 U380 ( .A(n537), .B(n362), .ZN(n596) );
  XNOR2_X1 U381 ( .A(n469), .B(n527), .ZN(n506) );
  XNOR2_X1 U382 ( .A(n463), .B(n462), .ZN(n433) );
  AND2_X1 U383 ( .A1(n455), .A2(n456), .ZN(n454) );
  XNOR2_X1 U384 ( .A(n559), .B(KEYINPUT19), .ZN(n600) );
  NOR2_X1 U385 ( .A1(n601), .A2(n600), .ZN(n603) );
  XNOR2_X1 U386 ( .A(n746), .B(KEYINPUT124), .ZN(n747) );
  INV_X1 U387 ( .A(n680), .ZN(n523) );
  AND2_X1 U388 ( .A1(n649), .A2(G475), .ZN(n439) );
  OR2_X1 U389 ( .A1(n717), .A2(n590), .ZN(n572) );
  XNOR2_X2 U390 ( .A(n403), .B(n488), .ZN(n763) );
  XNOR2_X2 U391 ( .A(n516), .B(KEYINPUT4), .ZN(n403) );
  NAND2_X1 U392 ( .A1(n703), .A2(n752), .ZN(n701) );
  INV_X1 U393 ( .A(KEYINPUT3), .ZN(n389) );
  INV_X1 U394 ( .A(KEYINPUT106), .ZN(n390) );
  INV_X1 U395 ( .A(n701), .ZN(n358) );
  AND2_X1 U396 ( .A1(n394), .A2(n643), .ZN(n378) );
  XNOR2_X1 U397 ( .A(n436), .B(n435), .ZN(n595) );
  NAND2_X1 U398 ( .A1(n437), .A2(n551), .ZN(n436) );
  XNOR2_X1 U399 ( .A(n603), .B(n602), .ZN(n691) );
  NAND2_X1 U400 ( .A1(n399), .A2(n558), .ZN(n398) );
  XNOR2_X1 U401 ( .A(n452), .B(n574), .ZN(n599) );
  XNOR2_X1 U402 ( .A(n397), .B(KEYINPUT0), .ZN(n640) );
  NOR2_X1 U403 ( .A1(n600), .A2(n564), .ZN(n397) );
  XNOR2_X1 U404 ( .A(n572), .B(KEYINPUT95), .ZN(n639) );
  OR2_X1 U405 ( .A1(n584), .A2(n579), .ZN(n680) );
  XNOR2_X1 U406 ( .A(n714), .B(n390), .ZN(n587) );
  AND2_X1 U407 ( .A1(n458), .A2(n457), .ZN(n456) );
  XNOR2_X1 U408 ( .A(n388), .B(n387), .ZN(n531) );
  XNOR2_X1 U409 ( .A(n389), .B(KEYINPUT71), .ZN(n388) );
  XOR2_X1 U410 ( .A(G116), .B(G107), .Z(n528) );
  XNOR2_X1 U411 ( .A(KEYINPUT15), .B(G902), .ZN(n647) );
  XNOR2_X1 U412 ( .A(G113), .B(G101), .ZN(n387) );
  NAND2_X1 U413 ( .A1(n358), .A2(n368), .ZN(n453) );
  OR2_X1 U414 ( .A1(n591), .A2(n590), .ZN(n601) );
  XNOR2_X2 U415 ( .A(n763), .B(G146), .ZN(n550) );
  INV_X1 U416 ( .A(KEYINPUT48), .ZN(n428) );
  XNOR2_X1 U417 ( .A(n382), .B(G104), .ZN(n530) );
  INV_X1 U418 ( .A(G122), .ZN(n382) );
  XOR2_X1 U419 ( .A(G146), .B(G125), .Z(n527) );
  XNOR2_X1 U420 ( .A(n539), .B(KEYINPUT91), .ZN(n727) );
  NAND2_X1 U421 ( .A1(n396), .A2(KEYINPUT44), .ZN(n395) );
  NAND2_X1 U422 ( .A1(n757), .A2(n534), .ZN(n535) );
  NAND2_X1 U423 ( .A1(n699), .A2(n406), .ZN(n405) );
  INV_X1 U424 ( .A(KEYINPUT85), .ZN(n406) );
  AND2_X1 U425 ( .A1(n616), .A2(KEYINPUT85), .ZN(n408) );
  INV_X1 U426 ( .A(n527), .ZN(n420) );
  XNOR2_X1 U427 ( .A(n526), .B(n418), .ZN(n417) );
  XNOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT90), .ZN(n418) );
  XOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n526) );
  XNOR2_X1 U430 ( .A(G134), .B(KEYINPUT101), .ZN(n510) );
  XNOR2_X1 U431 ( .A(n386), .B(n385), .ZN(n502) );
  XNOR2_X1 U432 ( .A(KEYINPUT98), .B(KEYINPUT12), .ZN(n386) );
  XNOR2_X1 U433 ( .A(G113), .B(G143), .ZN(n385) );
  XOR2_X1 U434 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n499) );
  XNOR2_X1 U435 ( .A(n530), .B(G131), .ZN(n498) );
  NAND2_X1 U436 ( .A1(n376), .A2(n374), .ZN(n373) );
  AND2_X1 U437 ( .A1(n571), .A2(n375), .ZN(n374) );
  NAND2_X1 U438 ( .A1(n727), .A2(n360), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n584) );
  XNOR2_X1 U440 ( .A(n509), .B(G475), .ZN(n383) );
  OR2_X1 U441 ( .A1(n668), .A2(G902), .ZN(n384) );
  INV_X1 U442 ( .A(KEYINPUT6), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n441), .B(n440), .ZN(n469) );
  INV_X1 U444 ( .A(G140), .ZN(n440) );
  XNOR2_X1 U445 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n441) );
  XNOR2_X1 U446 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n462) );
  XNOR2_X1 U447 ( .A(n543), .B(n542), .ZN(n437) );
  NAND2_X1 U448 ( .A1(n640), .A2(n620), .ZN(n621) );
  BUF_X1 U449 ( .A(n633), .Z(n413) );
  AND2_X1 U450 ( .A1(n649), .A2(G210), .ZN(n427) );
  INV_X1 U451 ( .A(KEYINPUT83), .ZN(n449) );
  INV_X1 U452 ( .A(KEYINPUT82), .ZN(n645) );
  OR2_X1 U453 ( .A1(n360), .A2(n727), .ZN(n377) );
  NOR2_X1 U454 ( .A1(n712), .A2(n485), .ZN(n495) );
  INV_X1 U455 ( .A(G137), .ZN(n486) );
  NAND2_X1 U456 ( .A1(n647), .A2(n645), .ZN(n457) );
  XNOR2_X1 U457 ( .A(n419), .B(n416), .ZN(n534) );
  XNOR2_X1 U458 ( .A(n417), .B(n525), .ZN(n416) );
  XNOR2_X1 U459 ( .A(n400), .B(n401), .ZN(n532) );
  XNOR2_X1 U460 ( .A(n531), .B(n402), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n528), .B(KEYINPUT16), .ZN(n402) );
  NAND2_X1 U462 ( .A1(G234), .A2(G237), .ZN(n477) );
  OR2_X1 U463 ( .A1(G237), .A2(G902), .ZN(n538) );
  INV_X1 U464 ( .A(n495), .ZN(n434) );
  INV_X1 U465 ( .A(n532), .ZN(n757) );
  XNOR2_X1 U466 ( .A(G122), .B(KEYINPUT102), .ZN(n512) );
  XNOR2_X1 U467 ( .A(n508), .B(n507), .ZN(n668) );
  INV_X1 U468 ( .A(n506), .ZN(n507) );
  XNOR2_X1 U469 ( .A(n505), .B(n504), .ZN(n508) );
  XNOR2_X1 U470 ( .A(G110), .B(G107), .ZN(n544) );
  XNOR2_X1 U471 ( .A(G101), .B(G104), .ZN(n546) );
  NAND2_X1 U472 ( .A1(n358), .A2(KEYINPUT2), .ZN(n649) );
  AND2_X1 U473 ( .A1(n557), .A2(n413), .ZN(n399) );
  AND2_X1 U474 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U475 ( .A1(n573), .A2(n639), .ZN(n452) );
  NOR2_X1 U476 ( .A1(n373), .A2(n372), .ZN(n573) );
  XNOR2_X1 U477 ( .A(n468), .B(n467), .ZN(n471) );
  NAND2_X1 U478 ( .A1(n379), .A2(n612), .ZN(n613) );
  INV_X1 U479 ( .A(KEYINPUT40), .ZN(n581) );
  INV_X1 U480 ( .A(KEYINPUT115), .ZN(n435) );
  AND2_X1 U481 ( .A1(n460), .A2(n424), .ZN(n422) );
  AND2_X1 U482 ( .A1(n622), .A2(n424), .ZN(n423) );
  INV_X1 U483 ( .A(KEYINPUT56), .ZN(n414) );
  XNOR2_X1 U484 ( .A(n446), .B(n445), .ZN(G75) );
  INV_X1 U485 ( .A(KEYINPUT53), .ZN(n445) );
  NOR2_X1 U486 ( .A1(n743), .A2(n366), .ZN(n447) );
  XOR2_X1 U487 ( .A(KEYINPUT21), .B(n484), .Z(n359) );
  XOR2_X1 U488 ( .A(n570), .B(KEYINPUT111), .Z(n360) );
  NOR2_X1 U489 ( .A1(n501), .A2(n656), .ZN(n361) );
  AND2_X1 U490 ( .A1(G210), .A2(n538), .ZN(n362) );
  XOR2_X1 U491 ( .A(n621), .B(KEYINPUT22), .Z(n363) );
  INV_X1 U492 ( .A(n712), .ZN(n424) );
  AND2_X1 U493 ( .A1(n639), .A2(n392), .ZN(n364) );
  AND2_X1 U494 ( .A1(n617), .A2(n405), .ZN(n365) );
  INV_X1 U495 ( .A(G902), .ZN(n521) );
  OR2_X1 U496 ( .A1(n711), .A2(G953), .ZN(n366) );
  XNOR2_X1 U497 ( .A(n578), .B(KEYINPUT39), .ZN(n367) );
  NOR2_X1 U498 ( .A1(n647), .A2(n645), .ZN(n368) );
  XOR2_X1 U499 ( .A(n650), .B(n652), .Z(n369) );
  XOR2_X1 U500 ( .A(n668), .B(n667), .Z(n370) );
  INV_X1 U501 ( .A(G210), .ZN(n656) );
  NAND2_X1 U502 ( .A1(n427), .A2(n371), .ZN(n426) );
  NAND2_X2 U503 ( .A1(n454), .A2(n453), .ZN(n371) );
  NAND2_X1 U504 ( .A1(n371), .A2(n649), .ZN(n744) );
  NAND2_X1 U505 ( .A1(n439), .A2(n371), .ZN(n411) );
  NAND2_X1 U506 ( .A1(n438), .A2(n371), .ZN(n412) );
  AND2_X1 U507 ( .A1(n587), .A2(n360), .ZN(n372) );
  OR2_X1 U508 ( .A1(n587), .A2(n377), .ZN(n376) );
  XNOR2_X1 U509 ( .A(n429), .B(n428), .ZN(n410) );
  NAND2_X1 U510 ( .A1(n596), .A2(n540), .ZN(n421) );
  XNOR2_X1 U511 ( .A(n709), .B(n449), .ZN(n448) );
  NAND2_X1 U512 ( .A1(n448), .A2(n447), .ZN(n446) );
  NAND2_X1 U513 ( .A1(n410), .A2(n408), .ZN(n407) );
  XNOR2_X1 U514 ( .A(n426), .B(n659), .ZN(n425) );
  NAND2_X1 U515 ( .A1(n395), .A2(n378), .ZN(n393) );
  XNOR2_X2 U516 ( .A(n471), .B(n470), .ZN(n746) );
  INV_X1 U517 ( .A(n381), .ZN(n379) );
  XNOR2_X1 U518 ( .A(n381), .B(n380), .ZN(n541) );
  INV_X1 U519 ( .A(KEYINPUT114), .ZN(n380) );
  NAND2_X1 U520 ( .A1(n524), .A2(n523), .ZN(n381) );
  XNOR2_X1 U521 ( .A(n714), .B(n391), .ZN(n633) );
  NOR2_X1 U522 ( .A1(n636), .A2(n392), .ZN(n722) );
  INV_X1 U523 ( .A(n714), .ZN(n392) );
  XNOR2_X2 U524 ( .A(n450), .B(G472), .ZN(n714) );
  XNOR2_X2 U525 ( .A(n393), .B(n644), .ZN(n752) );
  NAND2_X1 U526 ( .A1(n443), .A2(n442), .ZN(n394) );
  NAND2_X1 U527 ( .A1(n632), .A2(n631), .ZN(n396) );
  AND2_X2 U528 ( .A1(n737), .A2(n640), .ZN(n565) );
  XNOR2_X2 U529 ( .A(n398), .B(KEYINPUT33), .ZN(n737) );
  XNOR2_X1 U530 ( .A(n530), .B(n529), .ZN(n401) );
  XNOR2_X1 U531 ( .A(n403), .B(n420), .ZN(n419) );
  NOR2_X2 U532 ( .A1(n409), .A2(n404), .ZN(n703) );
  NAND2_X1 U533 ( .A1(n407), .A2(n365), .ZN(n404) );
  NOR2_X1 U534 ( .A1(n410), .A2(KEYINPUT85), .ZN(n409) );
  XNOR2_X1 U535 ( .A(n411), .B(n370), .ZN(n670) );
  XNOR2_X1 U536 ( .A(n451), .B(n367), .ZN(n580) );
  NAND2_X1 U537 ( .A1(n425), .A2(n669), .ZN(n415) );
  XNOR2_X1 U538 ( .A(n412), .B(n369), .ZN(n653) );
  XNOR2_X1 U539 ( .A(n415), .B(n414), .ZN(G51) );
  XNOR2_X2 U540 ( .A(n421), .B(KEYINPUT87), .ZN(n559) );
  NAND2_X1 U541 ( .A1(n363), .A2(n422), .ZN(n625) );
  NAND2_X1 U542 ( .A1(n363), .A2(n423), .ZN(n623) );
  NAND2_X1 U543 ( .A1(n431), .A2(n430), .ZN(n429) );
  AND2_X1 U544 ( .A1(n611), .A2(n610), .ZN(n430) );
  XNOR2_X1 U545 ( .A(n594), .B(n432), .ZN(n431) );
  INV_X1 U546 ( .A(KEYINPUT46), .ZN(n432) );
  NAND2_X1 U547 ( .A1(n433), .A2(G221), .ZN(n468) );
  AND2_X1 U548 ( .A1(n433), .A2(G217), .ZN(n520) );
  NOR2_X1 U549 ( .A1(n587), .A2(n434), .ZN(n589) );
  XNOR2_X1 U550 ( .A(n595), .B(KEYINPUT86), .ZN(n611) );
  AND2_X1 U551 ( .A1(n649), .A2(G472), .ZN(n438) );
  OR2_X2 U552 ( .A1(n650), .A2(G902), .ZN(n450) );
  NAND2_X1 U553 ( .A1(n629), .A2(n628), .ZN(n442) );
  NOR2_X1 U554 ( .A1(n774), .A2(n773), .ZN(n443) );
  XNOR2_X2 U555 ( .A(n444), .B(n673), .ZN(n590) );
  OR2_X2 U556 ( .A1(n674), .A2(G902), .ZN(n444) );
  XNOR2_X1 U557 ( .A(n550), .B(n549), .ZN(n674) );
  NAND2_X1 U558 ( .A1(n599), .A2(n577), .ZN(n451) );
  NAND2_X1 U559 ( .A1(n701), .A2(n645), .ZN(n455) );
  OR2_X1 U560 ( .A1(n764), .A2(G952), .ZN(n669) );
  XOR2_X1 U561 ( .A(n648), .B(KEYINPUT65), .Z(n458) );
  NOR2_X1 U562 ( .A1(n605), .A2(n604), .ZN(n459) );
  NOR2_X1 U563 ( .A1(n413), .A2(n718), .ZN(n460) );
  NOR2_X1 U564 ( .A1(n774), .A2(n630), .ZN(n632) );
  XNOR2_X1 U565 ( .A(n493), .B(n361), .ZN(n494) );
  XNOR2_X1 U566 ( .A(n466), .B(KEYINPUT24), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n582), .B(n581), .ZN(n660) );
  BUF_X1 U568 ( .A(n660), .Z(n661) );
  INV_X2 U569 ( .A(KEYINPUT64), .ZN(n461) );
  XNOR2_X2 U570 ( .A(n461), .B(G953), .ZN(n764) );
  NAND2_X1 U571 ( .A1(n764), .A2(G234), .ZN(n463) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n465) );
  XNOR2_X1 U573 ( .A(G137), .B(G128), .ZN(n464) );
  XNOR2_X1 U574 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U575 ( .A(G119), .B(G110), .Z(n529) );
  XNOR2_X1 U576 ( .A(n506), .B(n529), .ZN(n470) );
  NOR2_X2 U577 ( .A1(n746), .A2(G902), .ZN(n476) );
  XOR2_X1 U578 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n474) );
  NAND2_X1 U579 ( .A1(n647), .A2(G234), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n472), .B(KEYINPUT20), .ZN(n483) );
  NAND2_X1 U581 ( .A1(n483), .A2(G217), .ZN(n473) );
  XNOR2_X1 U582 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X2 U583 ( .A(n476), .B(n475), .ZN(n553) );
  BUF_X2 U584 ( .A(n553), .Z(n712) );
  XNOR2_X1 U585 ( .A(n477), .B(KEYINPUT92), .ZN(n478) );
  XNOR2_X1 U586 ( .A(KEYINPUT14), .B(n478), .ZN(n479) );
  NAND2_X1 U587 ( .A1(G952), .A2(n479), .ZN(n742) );
  NOR2_X1 U588 ( .A1(G953), .A2(n742), .ZN(n563) );
  NAND2_X1 U589 ( .A1(n479), .A2(G902), .ZN(n561) );
  OR2_X1 U590 ( .A1(n561), .A2(n764), .ZN(n480) );
  NOR2_X1 U591 ( .A1(G900), .A2(n480), .ZN(n481) );
  OR2_X1 U592 ( .A1(n563), .A2(n481), .ZN(n482) );
  XNOR2_X1 U593 ( .A(n482), .B(KEYINPUT80), .ZN(n571) );
  NAND2_X1 U594 ( .A1(G221), .A2(n483), .ZN(n484) );
  NAND2_X1 U595 ( .A1(n571), .A2(n359), .ZN(n485) );
  XNOR2_X2 U596 ( .A(G143), .B(G128), .ZN(n516) );
  XNOR2_X1 U597 ( .A(G134), .B(G131), .ZN(n487) );
  XNOR2_X1 U598 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U599 ( .A(G119), .B(G116), .ZN(n490) );
  XNOR2_X1 U600 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n489) );
  XNOR2_X1 U601 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n531), .B(n491), .ZN(n493) );
  NOR2_X1 U603 ( .A1(G953), .A2(G237), .ZN(n492) );
  XNOR2_X1 U604 ( .A(n492), .B(KEYINPUT75), .ZN(n501) );
  XNOR2_X1 U605 ( .A(n550), .B(n494), .ZN(n650) );
  NAND2_X1 U606 ( .A1(n495), .A2(n633), .ZN(n497) );
  INV_X1 U607 ( .A(KEYINPUT110), .ZN(n496) );
  XNOR2_X1 U608 ( .A(n497), .B(n496), .ZN(n524) );
  XNOR2_X1 U609 ( .A(n499), .B(n498), .ZN(n505) );
  INV_X1 U610 ( .A(G214), .ZN(n500) );
  NOR2_X1 U611 ( .A1(n501), .A2(n500), .ZN(n503) );
  XNOR2_X1 U612 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U613 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n509) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n511) );
  XNOR2_X1 U615 ( .A(n511), .B(n510), .ZN(n515) );
  XOR2_X1 U616 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n513) );
  XNOR2_X1 U617 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U618 ( .A(n515), .B(n514), .Z(n518) );
  XNOR2_X1 U619 ( .A(n516), .B(n528), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U621 ( .A(n520), .B(n519), .ZN(n663) );
  NAND2_X1 U622 ( .A1(n663), .A2(n521), .ZN(n522) );
  INV_X1 U623 ( .A(G478), .ZN(n662) );
  XNOR2_X1 U624 ( .A(n522), .B(n662), .ZN(n583) );
  INV_X1 U625 ( .A(n583), .ZN(n579) );
  NAND2_X1 U626 ( .A1(G224), .A2(n764), .ZN(n525) );
  INV_X1 U627 ( .A(n534), .ZN(n533) );
  NAND2_X1 U628 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U629 ( .A1(n536), .A2(n535), .ZN(n658) );
  NAND2_X1 U630 ( .A1(n658), .A2(n647), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n538), .A2(G214), .ZN(n539) );
  INV_X1 U632 ( .A(n727), .ZN(n540) );
  NAND2_X1 U633 ( .A1(n541), .A2(n559), .ZN(n543) );
  INV_X1 U634 ( .A(KEYINPUT36), .ZN(n542) );
  NAND2_X1 U635 ( .A1(n764), .A2(G227), .ZN(n545) );
  XNOR2_X1 U636 ( .A(n545), .B(n544), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n546), .B(G140), .ZN(n547) );
  XNOR2_X1 U638 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X1 U639 ( .A(G469), .ZN(n673) );
  XNOR2_X2 U640 ( .A(n590), .B(KEYINPUT1), .ZN(n718) );
  INV_X1 U641 ( .A(n718), .ZN(n551) );
  XOR2_X1 U642 ( .A(G125), .B(KEYINPUT37), .Z(n552) );
  XNOR2_X1 U643 ( .A(n595), .B(n552), .ZN(G27) );
  NAND2_X1 U644 ( .A1(n553), .A2(n359), .ZN(n554) );
  XNOR2_X1 U645 ( .A(n554), .B(KEYINPUT68), .ZN(n717) );
  OR2_X2 U646 ( .A1(n717), .A2(n718), .ZN(n636) );
  INV_X1 U647 ( .A(n636), .ZN(n556) );
  INV_X1 U648 ( .A(KEYINPUT108), .ZN(n555) );
  NAND2_X1 U649 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U650 ( .A1(n636), .A2(KEYINPUT108), .ZN(n557) );
  INV_X1 U651 ( .A(G953), .ZN(n751) );
  NOR2_X1 U652 ( .A1(n751), .A2(G898), .ZN(n560) );
  XNOR2_X1 U653 ( .A(n560), .B(KEYINPUT93), .ZN(n758) );
  NOR2_X1 U654 ( .A1(n561), .A2(n758), .ZN(n562) );
  NOR2_X1 U655 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U656 ( .A(n565), .B(KEYINPUT34), .ZN(n567) );
  OR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n566), .B(KEYINPUT109), .ZN(n597) );
  NAND2_X1 U659 ( .A1(n567), .A2(n597), .ZN(n569) );
  INV_X1 U660 ( .A(KEYINPUT35), .ZN(n568) );
  XNOR2_X2 U661 ( .A(n569), .B(n568), .ZN(n627) );
  XNOR2_X1 U662 ( .A(n627), .B(G122), .ZN(G24) );
  XNOR2_X1 U663 ( .A(KEYINPUT112), .B(KEYINPUT30), .ZN(n570) );
  INV_X1 U664 ( .A(KEYINPUT76), .ZN(n574) );
  INV_X1 U665 ( .A(n596), .ZN(n614) );
  INV_X1 U666 ( .A(KEYINPUT74), .ZN(n575) );
  XNOR2_X1 U667 ( .A(n575), .B(KEYINPUT38), .ZN(n576) );
  XNOR2_X1 U668 ( .A(n614), .B(n576), .ZN(n728) );
  INV_X1 U669 ( .A(n728), .ZN(n577) );
  INV_X1 U670 ( .A(KEYINPUT72), .ZN(n578) );
  NAND2_X1 U671 ( .A1(n584), .A2(n579), .ZN(n682) );
  OR2_X1 U672 ( .A1(n580), .A2(n682), .ZN(n617) );
  XNOR2_X1 U673 ( .A(n617), .B(G134), .ZN(G36) );
  NOR2_X2 U674 ( .A1(n580), .A2(n680), .ZN(n582) );
  NAND2_X1 U675 ( .A1(n584), .A2(n583), .ZN(n618) );
  NOR2_X1 U676 ( .A1(n727), .A2(n728), .ZN(n585) );
  XNOR2_X1 U677 ( .A(n585), .B(KEYINPUT113), .ZN(n733) );
  NOR2_X1 U678 ( .A1(n618), .A2(n733), .ZN(n586) );
  XNOR2_X1 U679 ( .A(n586), .B(KEYINPUT41), .ZN(n726) );
  INV_X1 U680 ( .A(KEYINPUT28), .ZN(n588) );
  XNOR2_X1 U681 ( .A(n589), .B(n588), .ZN(n591) );
  NOR2_X1 U682 ( .A1(n726), .A2(n601), .ZN(n592) );
  XNOR2_X1 U683 ( .A(n592), .B(KEYINPUT42), .ZN(n775) );
  INV_X1 U684 ( .A(n775), .ZN(n593) );
  NAND2_X1 U685 ( .A1(n660), .A2(n593), .ZN(n594) );
  AND2_X1 U686 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U687 ( .A1(n599), .A2(n598), .ZN(n690) );
  AND2_X1 U688 ( .A1(n680), .A2(n682), .ZN(n732) );
  INV_X1 U689 ( .A(n732), .ZN(n605) );
  INV_X1 U690 ( .A(KEYINPUT79), .ZN(n602) );
  NAND2_X1 U691 ( .A1(KEYINPUT73), .A2(n691), .ZN(n604) );
  OR2_X1 U692 ( .A1(n690), .A2(n459), .ZN(n609) );
  NOR2_X1 U693 ( .A1(n732), .A2(KEYINPUT73), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n691), .A2(n606), .ZN(n607) );
  XNOR2_X1 U695 ( .A(n607), .B(KEYINPUT47), .ZN(n608) );
  NOR2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n610) );
  AND2_X1 U697 ( .A1(n718), .A2(n540), .ZN(n612) );
  XNOR2_X1 U698 ( .A(n613), .B(KEYINPUT43), .ZN(n615) );
  AND2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n699) );
  INV_X1 U700 ( .A(n699), .ZN(n616) );
  INV_X1 U701 ( .A(n618), .ZN(n730) );
  NAND2_X1 U702 ( .A1(n730), .A2(n359), .ZN(n619) );
  XNOR2_X1 U703 ( .A(n619), .B(KEYINPUT105), .ZN(n620) );
  AND2_X1 U704 ( .A1(n587), .A2(n718), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n623), .B(KEYINPUT107), .ZN(n773) );
  INV_X1 U706 ( .A(KEYINPUT32), .ZN(n624) );
  XNOR2_X1 U707 ( .A(n625), .B(n624), .ZN(n774) );
  INV_X1 U708 ( .A(n627), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n630), .A2(KEYINPUT67), .ZN(n629) );
  NOR2_X1 U710 ( .A1(KEYINPUT67), .A2(KEYINPUT44), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U712 ( .A1(n773), .A2(KEYINPUT67), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n718), .A2(n712), .ZN(n634) );
  NOR2_X1 U714 ( .A1(n634), .A2(n413), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n363), .A2(n635), .ZN(n679) );
  NAND2_X1 U716 ( .A1(n640), .A2(n722), .ZN(n638) );
  XOR2_X1 U717 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n637) );
  XNOR2_X1 U718 ( .A(n638), .B(n637), .ZN(n697) );
  AND2_X1 U719 ( .A1(n640), .A2(n364), .ZN(n683) );
  OR2_X1 U720 ( .A1(n697), .A2(n683), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n641), .A2(n605), .ZN(n642) );
  AND2_X1 U722 ( .A1(n679), .A2(n642), .ZN(n643) );
  XNOR2_X1 U723 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n644) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n646) );
  OR2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U726 ( .A(KEYINPUT88), .B(KEYINPUT116), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n651), .B(KEYINPUT62), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n669), .ZN(n655) );
  XOR2_X1 U729 ( .A(KEYINPUT89), .B(KEYINPUT63), .Z(n654) );
  XNOR2_X1 U730 ( .A(n655), .B(n654), .ZN(G57) );
  XOR2_X1 U731 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  INV_X1 U733 ( .A(n669), .ZN(n750) );
  XNOR2_X1 U734 ( .A(n661), .B(G131), .ZN(G33) );
  NOR2_X1 U735 ( .A1(n744), .A2(n662), .ZN(n665) );
  XOR2_X1 U736 ( .A(KEYINPUT123), .B(n663), .Z(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U738 ( .A1(n666), .A2(n750), .ZN(G63) );
  XOR2_X1 U739 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n667) );
  NAND2_X1 U740 ( .A1(n670), .A2(n669), .ZN(n672) );
  XOR2_X1 U741 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G60) );
  NOR2_X1 U743 ( .A1(n744), .A2(n673), .ZN(n677) );
  XOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n675) );
  XOR2_X1 U745 ( .A(n675), .B(n674), .Z(n676) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n678), .A2(n750), .ZN(G54) );
  XNOR2_X1 U748 ( .A(G101), .B(n679), .ZN(G3) );
  NAND2_X1 U749 ( .A1(n683), .A2(n523), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n681), .B(G104), .ZN(G6) );
  XOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n685) );
  INV_X1 U752 ( .A(n682), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n683), .A2(n696), .ZN(n684) );
  XNOR2_X1 U754 ( .A(n685), .B(n684), .ZN(n687) );
  XOR2_X1 U755 ( .A(G107), .B(KEYINPUT117), .Z(n686) );
  XNOR2_X1 U756 ( .A(n687), .B(n686), .ZN(G9) );
  XOR2_X1 U757 ( .A(G128), .B(KEYINPUT29), .Z(n689) );
  NAND2_X1 U758 ( .A1(n691), .A2(n696), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n689), .B(n688), .ZN(G30) );
  XOR2_X1 U760 ( .A(G143), .B(n690), .Z(G45) );
  NAND2_X1 U761 ( .A1(n691), .A2(n523), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n692), .B(KEYINPUT118), .ZN(n693) );
  XNOR2_X1 U763 ( .A(G146), .B(n693), .ZN(G48) );
  XOR2_X1 U764 ( .A(G113), .B(KEYINPUT119), .Z(n695) );
  NAND2_X1 U765 ( .A1(n697), .A2(n523), .ZN(n694) );
  XNOR2_X1 U766 ( .A(n695), .B(n694), .ZN(G15) );
  NAND2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U768 ( .A(n698), .B(G116), .ZN(G18) );
  XOR2_X1 U769 ( .A(G140), .B(n699), .Z(G42) );
  INV_X1 U770 ( .A(KEYINPUT81), .ZN(n700) );
  XNOR2_X1 U771 ( .A(n702), .B(KEYINPUT2), .ZN(n708) );
  BUF_X1 U772 ( .A(n703), .Z(n704) );
  INV_X1 U773 ( .A(n704), .ZN(n705) );
  NAND2_X1 U774 ( .A1(n705), .A2(n752), .ZN(n706) );
  NAND2_X1 U775 ( .A1(n706), .A2(KEYINPUT81), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  INV_X1 U777 ( .A(n737), .ZN(n710) );
  NOR2_X1 U778 ( .A1(n726), .A2(n710), .ZN(n711) );
  NOR2_X1 U779 ( .A1(n712), .A2(n359), .ZN(n713) );
  XOR2_X1 U780 ( .A(KEYINPUT49), .B(n713), .Z(n715) );
  NOR2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U782 ( .A(n716), .B(KEYINPUT120), .Z(n721) );
  NAND2_X1 U783 ( .A1(n717), .A2(n718), .ZN(n719) );
  XOR2_X1 U784 ( .A(KEYINPUT50), .B(n719), .Z(n720) );
  NOR2_X1 U785 ( .A1(n721), .A2(n720), .ZN(n723) );
  NOR2_X1 U786 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U787 ( .A(KEYINPUT51), .B(n724), .Z(n725) );
  NOR2_X1 U788 ( .A1(n726), .A2(n725), .ZN(n739) );
  NAND2_X1 U789 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U790 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U791 ( .A(n731), .B(KEYINPUT121), .ZN(n735) );
  NOR2_X1 U792 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U795 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U796 ( .A(n740), .B(KEYINPUT52), .ZN(n741) );
  NOR2_X1 U797 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U798 ( .A(n744), .ZN(n745) );
  NAND2_X1 U799 ( .A1(n745), .A2(G217), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U801 ( .A1(n750), .A2(n749), .ZN(G66) );
  NAND2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n756) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n753) );
  XNOR2_X1 U804 ( .A(KEYINPUT61), .B(n753), .ZN(n754) );
  NAND2_X1 U805 ( .A1(n754), .A2(G898), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n756), .A2(n755), .ZN(n762) );
  XNOR2_X1 U807 ( .A(n757), .B(KEYINPUT125), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n760), .B(KEYINPUT126), .ZN(n761) );
  XOR2_X1 U810 ( .A(n762), .B(n761), .Z(G69) );
  XNOR2_X1 U811 ( .A(n763), .B(n506), .ZN(n768) );
  XNOR2_X1 U812 ( .A(n704), .B(n768), .ZN(n766) );
  INV_X1 U813 ( .A(n764), .ZN(n765) );
  NOR2_X1 U814 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U815 ( .A(KEYINPUT127), .B(n767), .ZN(n772) );
  XNOR2_X1 U816 ( .A(n768), .B(G227), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(G900), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n770), .A2(G953), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n772), .A2(n771), .ZN(G72) );
  XOR2_X1 U820 ( .A(G110), .B(n773), .Z(G12) );
  XOR2_X1 U821 ( .A(G119), .B(n774), .Z(G21) );
  XOR2_X1 U822 ( .A(G137), .B(n775), .Z(G39) );
endmodule

