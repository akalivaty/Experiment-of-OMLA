//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n211), .B2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n210), .A2(KEYINPUT64), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(G20), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n201), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n225), .B(new_n232), .C1(new_n235), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G58), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NOR3_X1   g0054(.A1(new_n228), .A2(new_n209), .A3(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n234), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n208), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G50), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n255), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(G50), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n257), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G33), .A3(new_n233), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT71), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(KEYINPUT9), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  OAI211_X1 g0076(.A(G1), .B(G13), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G222), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G223), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n275), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n282), .B(new_n285), .C1(new_n219), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n277), .B1(new_n290), .B2(KEYINPUT66), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(KEYINPUT66), .B2(new_n290), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n234), .B1(G33), .B2(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n277), .A2(new_n295), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n296), .B1(G226), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n292), .A2(G190), .A3(new_n299), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n274), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n274), .A2(new_n301), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n270), .B1(new_n300), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G179), .B2(new_n300), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n233), .A2(G33), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n267), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n219), .A2(new_n233), .B1(new_n264), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n257), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT68), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n255), .B2(new_n257), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n318), .A2(G77), .A3(new_n259), .A4(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n317), .B(new_n321), .C1(G77), .C2(new_n261), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n289), .A2(new_n283), .ZN(new_n323));
  INV_X1    g0123(.A(G232), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT67), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT67), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n281), .A2(new_n326), .A3(G232), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n280), .A2(G107), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n289), .A2(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n214), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n293), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n296), .B1(G244), .B2(new_n298), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(KEYINPUT70), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n331), .B1(new_n325), .B2(new_n327), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n339), .B2(new_n277), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n338), .B1(new_n340), .B2(new_n308), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(G179), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n322), .B(new_n337), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n322), .B1(new_n340), .B2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n344), .A2(new_n345), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  AOI211_X1 g0147(.A(KEYINPUT69), .B(new_n322), .C1(new_n340), .C2(G200), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n343), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT12), .B1(new_n261), .B2(G68), .ZN(new_n350));
  OR3_X1    g0150(.A1(new_n261), .A2(KEYINPUT12), .A3(G68), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n233), .A2(G33), .A3(G77), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n263), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n350), .A2(new_n351), .B1(new_n354), .B2(KEYINPUT11), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n318), .A2(G68), .A3(new_n259), .A4(new_n320), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(new_n356), .C1(KEYINPUT11), .C2(new_n354), .ZN(new_n357));
  INV_X1    g0157(.A(new_n295), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(new_n277), .A3(G274), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n297), .B2(new_n214), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n324), .A2(G1698), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n362), .B1(G226), .B2(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G97), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n293), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n277), .B1(new_n363), .B2(new_n364), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT13), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT14), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n372), .A3(G169), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(G179), .A3(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n371), .B2(G169), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n357), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n371), .A2(new_n346), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n368), .B2(new_n370), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n378), .A2(new_n380), .A3(new_n357), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n311), .A2(new_n349), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n359), .B1(new_n297), .B2(new_n324), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G226), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G1698), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n388), .B1(G223), .B2(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n293), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n346), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(G200), .B2(new_n393), .ZN(new_n395));
  INV_X1    g0195(.A(new_n258), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n265), .A2(new_n259), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n396), .A2(new_n397), .B1(new_n261), .B2(new_n265), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G58), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n213), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n401), .A2(new_n201), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(G20), .B1(G159), .B2(new_n267), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT7), .B1(new_n280), .B2(new_n233), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n287), .A2(new_n209), .A3(new_n288), .ZN(new_n405));
  AND2_X1   g0205(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n406));
  NOR2_X1   g0206(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT16), .B(new_n403), .C1(new_n410), .C2(new_n213), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n257), .ZN(new_n412));
  INV_X1    g0212(.A(new_n403), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n408), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n280), .A2(new_n233), .A3(KEYINPUT7), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT73), .B1(new_n405), .B2(new_n408), .ZN(new_n417));
  OAI21_X1  g0217(.A(G68), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(KEYINPUT74), .B(G68), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT16), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n395), .B(new_n399), .C1(new_n412), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n418), .A2(new_n419), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n403), .A3(new_n421), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT16), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n412), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n430), .A2(KEYINPUT17), .A3(new_n399), .A4(new_n395), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT76), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n386), .A2(new_n392), .A3(G179), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT75), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n277), .B1(new_n389), .B2(new_n390), .ZN(new_n437));
  OAI21_X1  g0237(.A(G169), .B1(new_n385), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n436), .B1(new_n435), .B2(new_n438), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n434), .B(new_n441), .C1(new_n429), .C2(new_n398), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n399), .B1(new_n422), .B2(new_n412), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n434), .B1(new_n444), .B2(new_n441), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n433), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n429), .B2(new_n398), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT18), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(KEYINPUT76), .A3(new_n442), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n432), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n384), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  XOR2_X1   g0252(.A(KEYINPUT80), .B(KEYINPUT19), .Z(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n312), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n289), .A2(new_n233), .A3(G68), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G33), .A3(G97), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(new_n233), .B1(new_n215), .B2(new_n205), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n452), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n453), .A2(new_n364), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n462), .A2(new_n466), .B1(G87), .B2(new_n206), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(KEYINPUT81), .A3(new_n456), .A4(new_n455), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n461), .A2(new_n468), .A3(new_n257), .ZN(new_n469));
  INV_X1    g0269(.A(new_n313), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n261), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n208), .A2(G33), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n258), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n472), .C1(new_n215), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n220), .A2(G1698), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n289), .B(new_n476), .C1(G238), .C2(G1698), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n277), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n277), .A2(new_n482), .A3(G250), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n277), .A2(G274), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n379), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(G190), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n475), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n474), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n470), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n469), .A2(new_n492), .A3(new_n472), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT82), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n469), .A2(new_n495), .A3(new_n492), .A4(new_n472), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n486), .A2(G169), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n335), .B2(new_n486), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n490), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  INV_X1    g0301(.A(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n255), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n233), .B(new_n504), .C1(G33), .C2(new_n454), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n256), .A2(new_n234), .B1(G20), .B2(new_n502), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(KEYINPUT20), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT20), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n208), .B2(G33), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n318), .A2(new_n320), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT83), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n318), .A2(KEYINPUT83), .A3(new_n320), .A4(new_n510), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n289), .A2(G257), .A3(new_n283), .ZN(new_n516));
  INV_X1    g0316(.A(G303), .ZN(new_n517));
  OAI221_X1 g0317(.A(new_n516), .B1(new_n517), .B2(new_n289), .C1(new_n330), .C2(new_n222), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n293), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT5), .B(G41), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n481), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n484), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n293), .B1(new_n481), .B2(new_n520), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(G270), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n519), .A2(G179), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n501), .B1(new_n515), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n514), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n507), .A2(new_n508), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n503), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n519), .A2(G179), .A3(new_n524), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(KEYINPUT84), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n519), .A2(new_n524), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G169), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n529), .A2(KEYINPUT21), .A3(G169), .A4(new_n534), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(G200), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n515), .B(new_n538), .C1(new_n346), .C2(new_n534), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n532), .A2(new_n536), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n289), .A2(G244), .A3(new_n283), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT78), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n543), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n289), .A2(new_n545), .A3(G244), .A4(new_n283), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n544), .A2(new_n504), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n293), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n522), .B1(G257), .B2(new_n523), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n335), .A3(new_n550), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n521), .A2(new_n484), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n523), .A2(G257), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n293), .B2(new_n548), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n555), .B2(G169), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n261), .A2(G97), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n491), .B2(G97), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT6), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n560), .A2(new_n454), .A3(G107), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n466), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n267), .A2(G77), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT77), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n416), .A2(new_n417), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n565), .B(new_n567), .C1(new_n568), .C2(new_n221), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n559), .B1(new_n569), .B2(new_n257), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT79), .B1(new_n556), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n233), .B2(new_n563), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n416), .A2(new_n417), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n558), .B1(new_n574), .B2(new_n263), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n549), .A2(new_n550), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n308), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .A4(new_n551), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n555), .A2(G190), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n570), .B(new_n580), .C1(new_n379), .C2(new_n555), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n571), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n289), .A2(G257), .A3(G1698), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G294), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n323), .C2(new_n216), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(new_n293), .B1(new_n523), .B2(G264), .ZN(new_n586));
  AOI21_X1  g0386(.A(G169), .B1(new_n586), .B2(new_n552), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n586), .A2(new_n552), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n335), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n289), .A2(new_n233), .A3(G87), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n591), .B(KEYINPUT22), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT23), .A2(G107), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n466), .A2(KEYINPUT85), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n478), .A2(G20), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n221), .A2(G20), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(KEYINPUT23), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT85), .B1(new_n466), .B2(new_n593), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n590), .B1(new_n592), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n592), .A2(new_n600), .A3(new_n590), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n263), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n228), .A2(G1), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(G20), .A3(new_n221), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT25), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n491), .B2(G107), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n589), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n603), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n257), .B1(new_n611), .B2(new_n601), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n588), .A2(G190), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n586), .A2(new_n552), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n612), .A2(new_n613), .A3(new_n608), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n582), .A2(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n451), .A2(new_n500), .A3(new_n540), .A4(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n497), .A2(new_n499), .ZN(new_n620));
  INV_X1    g0420(.A(new_n490), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n571), .A2(new_n579), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g0423(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n627));
  OAI211_X1 g0427(.A(KEYINPUT86), .B(G200), .C1(new_n479), .C2(new_n485), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n488), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n475), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n497), .B2(new_n499), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n556), .A2(new_n570), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n625), .B1(new_n626), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n620), .ZN(new_n636));
  INV_X1    g0436(.A(new_n532), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n536), .A2(new_n537), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n610), .ZN(new_n640));
  INV_X1    g0440(.A(new_n616), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n582), .A2(new_n641), .A3(new_n631), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n636), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n451), .B1(new_n635), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n343), .A2(new_n381), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n432), .B1(new_n377), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n435), .A2(new_n438), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n429), .B2(new_n398), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT18), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n444), .A2(new_n434), .A3(new_n648), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n307), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n310), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n233), .A2(new_n605), .ZN(new_n658));
  OAI21_X1  g0458(.A(G213), .B1(new_n658), .B2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT88), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(new_n662), .A3(KEYINPUT27), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n659), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n657), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(KEYINPUT89), .A3(G343), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n529), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n540), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n639), .B2(new_n670), .ZN(new_n672));
  XOR2_X1   g0472(.A(KEYINPUT90), .B(G330), .Z(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n617), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n669), .B1(new_n604), .B2(new_n609), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n669), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n610), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n669), .B(KEYINPUT91), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n610), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n639), .A2(new_n669), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n230), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n205), .A2(new_n215), .A3(new_n502), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n690), .A2(new_n208), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n238), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT92), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  OR2_X1    g0495(.A1(new_n630), .A2(new_n475), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n620), .A2(KEYINPUT26), .A3(new_n696), .A4(new_n633), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT94), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n632), .A2(KEYINPUT94), .A3(KEYINPUT26), .A4(new_n633), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n623), .A2(new_n624), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n643), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n680), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n634), .A2(new_n626), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n623), .B2(new_n624), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n684), .B1(new_n706), .B2(new_n643), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n704), .B1(new_n707), .B2(KEYINPUT29), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n618), .A2(new_n500), .A3(new_n540), .A4(new_n683), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n549), .A2(new_n586), .A3(new_n486), .A4(new_n550), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT30), .B1(new_n711), .B2(new_n525), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n586), .A2(new_n486), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n530), .A2(new_n713), .A3(new_n714), .A4(new_n555), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n486), .A2(G179), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n577), .A2(new_n716), .A3(new_n534), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n712), .A2(new_n715), .B1(new_n717), .B2(new_n614), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n710), .B1(new_n718), .B2(new_n680), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n715), .A2(new_n712), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(new_n614), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n684), .A2(new_n724), .A3(KEYINPUT31), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n709), .A2(new_n720), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n674), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n708), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n695), .B1(new_n729), .B2(G1), .ZN(G364));
  NOR2_X1   g0530(.A1(new_n466), .A2(new_n228), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n208), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n690), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n676), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n674), .B2(new_n672), .ZN(new_n736));
  INV_X1    g0536(.A(new_n734), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n689), .A2(new_n280), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n738), .A2(G355), .B1(new_n502), .B2(new_n689), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n689), .A2(new_n289), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G45), .B2(new_n237), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n253), .A2(new_n480), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n308), .A2(KEYINPUT95), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n209), .B1(KEYINPUT95), .B2(new_n308), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n234), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n737), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n379), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G20), .A3(G190), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n466), .A2(new_n346), .A3(new_n755), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n280), .B1(new_n517), .B2(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n233), .A2(new_n335), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n346), .A3(new_n379), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n762), .A2(G326), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n761), .A2(G190), .A3(new_n379), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n759), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n233), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G329), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n346), .A2(G200), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n233), .B1(new_n335), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(G294), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n760), .A2(new_n773), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT97), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n779), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n766), .B(new_n776), .C1(new_n777), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n774), .A2(new_n454), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n289), .B1(new_n215), .B2(new_n756), .C1(new_n771), .C2(new_n219), .ZN(new_n786));
  INV_X1    g0586(.A(new_n757), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n785), .B(new_n786), .C1(G107), .C2(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G50), .A2(new_n762), .B1(new_n764), .B2(G68), .ZN(new_n789));
  INV_X1    g0589(.A(new_n783), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G58), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n767), .A2(G159), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT32), .Z(new_n793));
  NAND4_X1  g0593(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n784), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n753), .B(new_n754), .C1(new_n747), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n750), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n672), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n736), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  NAND2_X1  g0600(.A1(new_n669), .A2(new_n322), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n343), .B(new_n801), .C1(new_n347), .C2(new_n348), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n341), .A2(new_n342), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n803), .A2(new_n322), .A3(new_n337), .A4(new_n669), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n707), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n734), .B1(new_n806), .B2(new_n727), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n727), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n747), .A2(new_n748), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n734), .B1(G77), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n790), .A2(G294), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n762), .A2(G303), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n280), .B1(new_n756), .B2(new_n221), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n814), .B(new_n785), .C1(new_n764), .C2(G283), .ZN(new_n815));
  INV_X1    g0615(.A(new_n767), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n816), .A2(new_n769), .B1(new_n502), .B2(new_n771), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G87), .B2(new_n787), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n771), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n762), .A2(G137), .B1(G159), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  INV_X1    g0622(.A(new_n764), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT98), .B(G143), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n821), .B1(new_n822), .B2(new_n823), .C1(new_n783), .C2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  AOI22_X1  g0626(.A1(new_n775), .A2(G58), .B1(new_n767), .B2(G132), .ZN(new_n827));
  INV_X1    g0627(.A(new_n756), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n280), .B1(new_n828), .B2(G50), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(new_n213), .C2(new_n757), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n819), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n811), .B1(new_n831), .B2(new_n747), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n749), .B2(new_n805), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n808), .A2(new_n833), .ZN(G384));
  NOR2_X1   g0634(.A1(new_n731), .A2(new_n208), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT39), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n444), .A2(new_n664), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n837), .A2(new_n447), .A3(new_n838), .A4(new_n423), .ZN(new_n839));
  OAI21_X1  g0639(.A(G68), .B1(new_n404), .B2(new_n409), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT16), .B1(new_n840), .B2(new_n403), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n399), .B1(new_n412), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n648), .B2(new_n664), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n423), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n839), .B1(new_n844), .B2(new_n838), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n664), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n450), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(KEYINPUT38), .B(new_n845), .C1(new_n450), .C2(new_n846), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(KEYINPUT99), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT99), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n847), .A2(new_n852), .A3(new_n848), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n836), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n650), .A2(new_n425), .A3(new_n431), .A4(new_n651), .ZN(new_n855));
  INV_X1    g0655(.A(new_n837), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT100), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n837), .A2(new_n423), .A3(new_n649), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n857), .A2(new_n858), .B1(new_n839), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n855), .A2(KEYINPUT100), .A3(new_n856), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT39), .B1(new_n864), .B2(new_n850), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n371), .A2(G169), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT14), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n374), .A3(new_n373), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n357), .A3(new_n680), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n854), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n683), .B(new_n805), .C1(new_n635), .C2(new_n644), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n343), .A2(new_n669), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n669), .A2(new_n357), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n377), .A2(new_n382), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n357), .B(new_n669), .C1(new_n868), .C2(new_n381), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n851), .A2(new_n853), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n879), .A2(new_n880), .B1(new_n652), .B2(new_n664), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n704), .B(new_n451), .C1(new_n707), .C2(KEYINPUT29), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n655), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT101), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n883), .B(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n878), .A2(new_n805), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(new_n719), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n888), .B(new_n889), .C1(new_n709), .C2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n850), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n863), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(KEYINPUT103), .B(new_n892), .C1(new_n863), .C2(new_n893), .ZN(new_n897));
  AOI211_X1 g0697(.A(KEYINPUT102), .B(new_n889), .C1(new_n709), .C2(new_n891), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n709), .A2(new_n891), .ZN(new_n900));
  INV_X1    g0700(.A(new_n889), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n851), .A2(new_n903), .A3(new_n853), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n896), .A2(new_n897), .B1(new_n904), .B2(new_n888), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n451), .A2(new_n900), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n673), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n835), .B1(new_n887), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n887), .B2(new_n909), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n564), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n564), .A2(KEYINPUT35), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(G116), .A3(new_n235), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n237), .A2(new_n219), .A3(new_n401), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n213), .A2(G50), .ZN(new_n917));
  OAI211_X1 g0717(.A(G1), .B(new_n228), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n911), .A2(new_n915), .A3(new_n918), .ZN(G367));
  INV_X1    g0719(.A(new_n622), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(new_n581), .C1(new_n570), .C2(new_n683), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n684), .A2(new_n633), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n924), .B2(new_n610), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n683), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n686), .A2(new_n677), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT42), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n924), .A2(KEYINPUT42), .A3(new_n927), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n475), .A2(new_n669), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n632), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n620), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT104), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n935), .B1(new_n930), .B2(new_n937), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n682), .A2(new_n924), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n687), .A2(new_n923), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT45), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n687), .A2(new_n923), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n676), .A3(new_n681), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n682), .A3(new_n948), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n927), .B1(new_n681), .B2(new_n686), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n675), .B2(KEYINPUT105), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n675), .A2(KEYINPUT105), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n729), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n690), .B(KEYINPUT41), .Z(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n944), .B1(new_n960), .B2(new_n733), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n689), .A2(new_n246), .A3(new_n289), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n751), .B1(new_n230), .B2(new_n313), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n734), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n775), .A2(G68), .ZN(new_n965));
  INV_X1    g0765(.A(G137), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n965), .B1(new_n202), .B2(new_n771), .C1(new_n966), .C2(new_n816), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n757), .A2(new_n219), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n280), .B(new_n968), .C1(G58), .C2(new_n828), .ZN(new_n969));
  INV_X1    g0769(.A(new_n762), .ZN(new_n970));
  INV_X1    g0770(.A(G159), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n969), .B1(new_n970), .B2(new_n824), .C1(new_n971), .C2(new_n823), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n967), .B(new_n972), .C1(G150), .C2(new_n790), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n502), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT46), .B1(new_n756), .B2(new_n502), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n289), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(G294), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n976), .B1(new_n970), .B2(new_n769), .C1(new_n977), .C2(new_n823), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n783), .A2(new_n517), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n787), .A2(G97), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n758), .B2(new_n771), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n816), .A2(new_n982), .B1(new_n221), .B2(new_n774), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n978), .A2(new_n979), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT47), .Z(new_n986));
  AOI21_X1  g0786(.A(new_n964), .B1(new_n986), .B2(new_n747), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n933), .B2(new_n797), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n961), .A2(new_n988), .ZN(G387));
  AOI22_X1  g0789(.A1(new_n738), .A2(new_n691), .B1(new_n221), .B2(new_n689), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n243), .A2(new_n480), .ZN(new_n991));
  AOI211_X1 g0791(.A(G45), .B(new_n691), .C1(G68), .C2(G77), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n265), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT50), .B1(new_n265), .B2(new_n202), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n740), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n990), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n750), .B(new_n747), .C1(new_n997), .C2(KEYINPUT106), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(KEYINPUT106), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n737), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n681), .B2(new_n797), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n280), .B1(new_n828), .B2(G77), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n980), .B(new_n1002), .C1(new_n816), .C2(new_n822), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT107), .Z(new_n1004));
  AOI22_X1  g0804(.A1(new_n820), .A2(G68), .B1(new_n775), .B2(new_n470), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n823), .B2(new_n264), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G159), .B2(new_n762), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1004), .B(new_n1007), .C1(new_n202), .C2(new_n783), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n289), .B1(new_n767), .B2(G326), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n774), .A2(new_n758), .B1(new_n977), .B2(new_n756), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n764), .A2(G311), .B1(G303), .B2(new_n820), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n777), .B2(new_n970), .C1(new_n783), .C2(new_n982), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT48), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1009), .B1(new_n502), .B2(new_n757), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1008), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1001), .B1(new_n747), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT108), .Z(new_n1021));
  INV_X1    g0821(.A(new_n956), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n729), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n690), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1022), .A2(new_n729), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1021), .B1(new_n732), .B2(new_n956), .C1(new_n1024), .C2(new_n1025), .ZN(G393));
  NAND3_X1  g0826(.A1(new_n950), .A2(new_n733), .A3(new_n951), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n740), .A2(new_n250), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n751), .B1(new_n230), .B2(new_n454), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n734), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n289), .B1(new_n213), .B2(new_n756), .C1(new_n757), .C2(new_n215), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n775), .A2(G77), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n264), .B2(new_n771), .C1(new_n816), .C2(new_n824), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(G50), .C2(new_n764), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n790), .A2(G159), .B1(G150), .B2(new_n762), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT51), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT109), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n783), .A2(new_n769), .B1(new_n982), .B2(new_n970), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT52), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n289), .B1(new_n828), .B2(G283), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n221), .B2(new_n757), .C1(new_n816), .C2(new_n777), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT110), .Z(new_n1046));
  NAND2_X1  g0846(.A1(new_n764), .A2(G303), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n820), .A2(G294), .B1(new_n775), .B2(G116), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1041), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1030), .B1(new_n1051), .B2(new_n747), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n923), .B2(new_n797), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1027), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT111), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n952), .A2(new_n1023), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n952), .A2(new_n1023), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n1057), .A3(new_n690), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT112), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1055), .A2(KEYINPUT112), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(new_n805), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n669), .B(new_n1064), .C1(new_n702), .C2(new_n643), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(new_n872), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n726), .A2(new_n674), .A3(new_n805), .A4(new_n878), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n878), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n900), .A2(G330), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n1064), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1066), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n727), .B2(new_n1064), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1069), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n901), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n874), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n451), .A2(new_n1073), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n884), .A2(new_n655), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n865), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1068), .B1(new_n871), .B2(new_n873), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n869), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n878), .B1(new_n1065), .B2(new_n872), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n864), .A2(new_n850), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n869), .B(KEYINPUT113), .Z(new_n1090));
  AND2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1083), .A2(new_n1087), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n1074), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n854), .A2(new_n865), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1067), .C1(new_n1095), .C2(new_n1086), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1080), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n884), .A2(new_n655), .A3(new_n1078), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1076), .B2(new_n1071), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1096), .B(new_n1100), .C1(new_n1092), .C2(new_n1074), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n690), .A3(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1032), .B1(new_n454), .B2(new_n771), .C1(new_n977), .C2(new_n816), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n280), .B1(new_n756), .B2(new_n215), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n787), .B2(G68), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n970), .B2(new_n758), .C1(new_n221), .C2(new_n823), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(G116), .C2(new_n790), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n762), .A2(G128), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n828), .A2(G150), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT53), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n280), .B1(new_n1109), .B2(KEYINPUT53), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT54), .B(G143), .Z(new_n1113));
  AOI22_X1  g0913(.A1(new_n820), .A2(new_n1113), .B1(new_n775), .B2(G159), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G125), .A2(new_n767), .B1(new_n787), .B2(G50), .ZN(new_n1115));
  INV_X1    g0915(.A(G132), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1115), .C1(new_n783), .C2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1112), .B(new_n1117), .C1(G137), .C2(new_n764), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n747), .B1(new_n1107), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n734), .B1(new_n265), .B2(new_n810), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT114), .Z(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1083), .B2(new_n748), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n733), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1102), .A2(new_n1125), .ZN(G378));
  NAND2_X1  g0926(.A1(new_n1101), .A2(new_n1079), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n896), .A2(new_n897), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n904), .A2(new_n888), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(G330), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n665), .A2(new_n270), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n311), .B(new_n1131), .Z(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n905), .A2(G330), .A3(new_n1134), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT118), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n870), .B2(new_n881), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n880), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(new_n1084), .B1(new_n653), .B2(new_n665), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1081), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT118), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1138), .A2(KEYINPUT119), .A3(new_n1140), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1134), .B1(new_n905), .B2(G330), .ZN(new_n1146));
  AND4_X1   g0946(.A1(G330), .A2(new_n1128), .A3(new_n1129), .A4(new_n1134), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1136), .A2(new_n1137), .A3(new_n882), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT119), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1127), .B(new_n1145), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n690), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1155), .B1(new_n1101), .B2(new_n1079), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1138), .A2(new_n883), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1151), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1157), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n733), .B(new_n1145), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n734), .B1(G50), .B2(new_n810), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n820), .A2(G137), .B1(new_n828), .B2(new_n1113), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n823), .B2(new_n1116), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n762), .A2(G125), .B1(G150), .B2(new_n775), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT115), .Z(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(G128), .C2(new_n790), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT59), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT116), .B(G124), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n275), .B(new_n276), .C1(new_n816), .C2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G159), .B2(new_n787), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n762), .A2(G116), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n280), .A2(new_n276), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n828), .B2(G77), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n965), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n757), .A2(new_n400), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n771), .A2(new_n313), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G283), .C2(new_n767), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n221), .B2(new_n783), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1180), .B(new_n1184), .C1(G97), .C2(new_n764), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1178), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1176), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1164), .B1(new_n1189), .B2(new_n747), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1134), .B2(new_n749), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT117), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1163), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1162), .A2(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1068), .A2(new_n748), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n734), .B1(G68), .B2(new_n810), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n289), .B(new_n968), .C1(G97), .C2(new_n828), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n502), .B2(new_n823), .C1(new_n977), .C2(new_n970), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n775), .A2(new_n470), .B1(new_n767), .B2(G303), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n221), .B2(new_n771), .C1(new_n783), .C2(new_n758), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G132), .A2(new_n762), .B1(new_n764), .B2(new_n1113), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n289), .B1(new_n756), .B2(new_n971), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1206), .B(new_n1181), .C1(G128), .C2(new_n767), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(new_n966), .C2(new_n783), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n771), .A2(new_n822), .B1(new_n774), .B2(new_n202), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT121), .Z(new_n1210));
  OAI22_X1  g1010(.A1(new_n1202), .A2(new_n1204), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1200), .B1(new_n1211), .B2(new_n747), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1077), .A2(new_n733), .B1(new_n1199), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1100), .A2(new_n958), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1099), .A2(new_n1076), .A3(new_n1071), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(G381));
  AND2_X1   g1018(.A1(new_n961), .A2(new_n988), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1217), .A3(new_n1220), .ZN(new_n1221));
  OR4_X1    g1021(.A1(G390), .A2(G375), .A3(G378), .A4(new_n1221), .ZN(G407));
  NAND2_X1  g1022(.A1(new_n666), .A2(G213), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT122), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1197), .A2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(new_n1225), .C2(new_n1227), .ZN(G409));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1062), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT112), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1219), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1061), .A2(G387), .A3(new_n1062), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT125), .B1(G390), .B2(new_n1219), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(G393), .B(new_n799), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1232), .A2(KEYINPUT125), .A3(new_n1233), .A4(new_n1236), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1162), .A2(G378), .A3(new_n1193), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1160), .A2(new_n733), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1191), .B(new_n1243), .C1(new_n1154), .C2(new_n958), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1226), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1080), .A2(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1216), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1099), .A2(KEYINPUT60), .A3(new_n1071), .A4(new_n1076), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n690), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(G384), .A3(new_n1213), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1250), .B1(new_n1247), .B2(new_n1216), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1214), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(KEYINPUT123), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT123), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT62), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1246), .A2(new_n1225), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT123), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G384), .B1(new_n1252), .B2(new_n1213), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1255), .A2(new_n1254), .A3(new_n1214), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1257), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1246), .A2(new_n1223), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1224), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(KEYINPUT126), .A3(new_n1261), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1264), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  INV_X1    g1076(.A(G2897), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1258), .A2(new_n1259), .B1(new_n1277), .B2(new_n1223), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(G2897), .A3(new_n1224), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1223), .A2(new_n1277), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(new_n1268), .B2(new_n1257), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1279), .A2(new_n1277), .A3(new_n1225), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT124), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1276), .B1(new_n1288), .B2(new_n1273), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1241), .B1(new_n1275), .B2(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1238), .A2(new_n1276), .A3(new_n1239), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1270), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1246), .A2(new_n1223), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1283), .A3(new_n1287), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1273), .A2(KEYINPUT63), .A3(new_n1269), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1292), .A2(new_n1294), .A3(new_n1296), .A4(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1229), .B1(new_n1291), .B2(new_n1299), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n1224), .B(new_n1260), .C1(new_n1242), .C2(new_n1245), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(KEYINPUT126), .A2(new_n1301), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1289), .B1(new_n1302), .B2(new_n1264), .ZN(new_n1303));
  OAI211_X1 g1103(.A(KEYINPUT127), .B(new_n1298), .C1(new_n1303), .C2(new_n1241), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(G405));
  NAND2_X1  g1105(.A1(new_n1194), .A2(G378), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1227), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1280), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1227), .A2(new_n1269), .A3(new_n1306), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1308), .A2(new_n1240), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1240), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


