//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n189), .A3(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G122), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n188), .A2(KEYINPUT13), .A3(new_n191), .ZN(new_n196));
  OAI21_X1  g010(.A(G134), .B1(new_n188), .B2(KEYINPUT13), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n192), .B(new_n195), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G122), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G116), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n194), .B1(new_n200), .B2(KEYINPUT14), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n201), .B(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(new_n192), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n189), .B1(new_n188), .B2(new_n191), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT9), .B(G234), .ZN(new_n207));
  INV_X1    g021(.A(G217), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n207), .A2(new_n208), .A3(G953), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n198), .A2(new_n205), .A3(new_n209), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT69), .B(G902), .Z(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G478), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n215), .A2(new_n221), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n222), .A2(KEYINPUT89), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT89), .B1(new_n222), .B2(new_n223), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(G237), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(G214), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n187), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT67), .A2(G237), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT67), .A2(G237), .ZN(new_n233));
  AOI21_X1  g047(.A(G953), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G143), .A3(G214), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n231), .A2(new_n239), .A3(new_n235), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G125), .ZN(new_n242));
  OR3_X1    g056(.A1(new_n242), .A2(KEYINPUT16), .A3(G140), .ZN(new_n243));
  XOR2_X1   g057(.A(G125), .B(G140), .Z(new_n244));
  INV_X1    g058(.A(KEYINPUT16), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n249));
  OAI211_X1 g063(.A(G146), .B(new_n243), .C1(new_n244), .C2(new_n245), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(KEYINPUT71), .A3(new_n247), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n239), .B1(new_n231), .B2(new_n235), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT17), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n241), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G113), .B(G122), .ZN(new_n257));
  INV_X1    g071(.A(G104), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT18), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n231), .B(new_n235), .C1(new_n260), .C2(new_n239), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n244), .A2(G146), .ZN(new_n262));
  XNOR2_X1  g076(.A(G125), .B(G140), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n247), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n261), .B(new_n265), .C1(new_n237), .C2(new_n260), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n256), .A2(new_n259), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n259), .B1(new_n256), .B2(new_n266), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n227), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G475), .ZN(new_n270));
  INV_X1    g084(.A(G952), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n271), .A2(KEYINPUT90), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(KEYINPUT90), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n229), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(G234), .B2(G237), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n229), .B(new_n214), .C1(G234), .C2(G237), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT21), .B(G898), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n278), .B(KEYINPUT91), .Z(new_n279));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n263), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n263), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n250), .B1(new_n284), .B2(G146), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT87), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n250), .B(new_n287), .C1(new_n284), .C2(G146), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n240), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n254), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n266), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n259), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n256), .A2(new_n259), .A3(new_n266), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G475), .A2(G902), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n280), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  AOI211_X1 g113(.A(KEYINPUT20), .B(new_n299), .C1(new_n294), .C2(new_n295), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n270), .B(new_n279), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n226), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n207), .B2(G902), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n247), .A2(G143), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n187), .B2(G146), .ZN(new_n307));
  AND2_X1   g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NOR2_X1   g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G143), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G146), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n187), .B2(G146), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n307), .A2(new_n310), .B1(new_n313), .B2(new_n308), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n194), .A3(G104), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n258), .A2(KEYINPUT74), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G104), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n320), .A3(G107), .ZN(new_n321));
  AOI21_X1  g135(.A(G107), .B1(new_n318), .B2(new_n320), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n317), .B(new_n321), .C1(new_n322), .C2(new_n316), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G101), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT74), .B(G104), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n325), .B2(G107), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n317), .A4(new_n321), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n315), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT4), .B1(new_n323), .B2(G101), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n314), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n194), .A2(G104), .ZN(new_n332));
  OAI21_X1  g146(.A(G101), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n317), .B1(new_n322), .B2(new_n316), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n327), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT75), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n338));
  OAI21_X1  g152(.A(G128), .B1(new_n312), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n307), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n311), .A2(KEYINPUT64), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G143), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(G146), .ZN(new_n344));
  INV_X1    g158(.A(new_n312), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n328), .A2(new_n349), .A3(new_n333), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n313), .B1(G128), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n347), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n328), .B(new_n333), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT65), .ZN(new_n358));
  INV_X1    g172(.A(G137), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT65), .A2(G137), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT11), .A2(G134), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT11), .A2(G134), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT11), .A2(G134), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(G137), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n363), .A2(new_n239), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n239), .B1(new_n363), .B2(new_n366), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n331), .A2(new_n351), .A3(new_n357), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n366), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G131), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n363), .A2(new_n366), .A3(new_n239), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT12), .B1(new_n374), .B2(KEYINPUT76), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n336), .A2(new_n340), .A3(new_n347), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n369), .B(new_n375), .C1(new_n355), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n375), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n355), .A2(new_n376), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(new_n374), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n370), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G140), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n229), .A2(G227), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n331), .A2(new_n351), .A3(new_n357), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n374), .ZN(new_n387));
  INV_X1    g201(.A(new_n384), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n370), .A3(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n385), .A2(KEYINPUT77), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT77), .B1(new_n385), .B2(new_n389), .ZN(new_n391));
  INV_X1    g205(.A(G469), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n377), .A2(new_n380), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n370), .A2(new_n388), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n388), .B1(new_n387), .B2(new_n370), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n392), .B(new_n214), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(G469), .A2(G902), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n304), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n400), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n385), .A2(new_n389), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n385), .A2(KEYINPUT77), .A3(new_n389), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(G469), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(KEYINPUT78), .A3(new_n304), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n303), .B1(new_n403), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n344), .A2(new_n345), .A3(new_n308), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n341), .A2(new_n343), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n305), .B1(new_n414), .B2(new_n247), .ZN(new_n415));
  INV_X1    g229(.A(new_n310), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n242), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n242), .B2(new_n348), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT83), .B(G224), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n229), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n419), .B(new_n421), .Z(new_n422));
  INV_X1    g236(.A(G119), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G116), .ZN(new_n424));
  INV_X1    g238(.A(G116), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G119), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT2), .B(G113), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n428), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n329), .B2(new_n330), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT5), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n434), .B(G113), .C1(KEYINPUT5), .C2(new_n424), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n435), .A2(new_n429), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n337), .A2(new_n433), .A3(new_n350), .A4(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n337), .A2(new_n350), .A3(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT80), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G122), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n438), .A2(KEYINPUT6), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n432), .A3(new_n437), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT6), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n441), .B(KEYINPUT81), .Z(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n446), .B1(new_n443), .B2(new_n447), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n422), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n421), .A2(KEYINPUT7), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n336), .A2(new_n436), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n441), .B(KEYINPUT8), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n336), .B2(new_n436), .ZN(new_n455));
  OAI22_X1  g269(.A1(new_n419), .A2(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n419), .A2(new_n452), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n419), .A2(KEYINPUT84), .A3(new_n452), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n451), .A2(new_n463), .A3(new_n465), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n468), .ZN(new_n469));
  AOI211_X1 g283(.A(KEYINPUT85), .B(new_n465), .C1(new_n451), .C2(new_n463), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G214), .B1(G237), .B2(G902), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n473), .B(KEYINPUT79), .Z(new_n474));
  NOR2_X1   g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n412), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G110), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G119), .B(G128), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT23), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n423), .B2(G128), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n482), .B(new_n483), .C1(G119), .C2(new_n190), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n479), .A2(new_n480), .B1(G110), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n251), .A2(new_n485), .A3(new_n252), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n479), .A2(new_n480), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n484), .A2(G110), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n250), .B(new_n264), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT22), .B(G137), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n490), .B(new_n494), .Z(new_n495));
  AOI21_X1  g309(.A(new_n208), .B1(new_n214), .B2(G234), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(KEYINPUT25), .A3(new_n214), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n490), .B(new_n494), .ZN(new_n501));
  INV_X1    g315(.A(new_n214), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n496), .B1(new_n503), .B2(KEYINPUT73), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n498), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G472), .A2(G902), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT66), .B1(new_n369), .B2(new_n417), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n314), .A2(new_n374), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n360), .A2(new_n189), .A3(new_n361), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n239), .B1(G134), .B2(G137), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n348), .A2(new_n373), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n508), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n314), .A2(new_n374), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n516), .A2(new_n508), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n431), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n234), .A2(G210), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT27), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n521), .B(KEYINPUT27), .ZN(new_n526));
  INV_X1    g340(.A(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n373), .A2(new_n515), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n340), .B2(new_n347), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n509), .B2(new_n511), .ZN(new_n532));
  INV_X1    g346(.A(new_n431), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n520), .A2(KEYINPUT68), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT68), .B1(new_n520), .B2(new_n534), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI211_X1 g352(.A(new_n431), .B(new_n531), .C1(new_n509), .C2(new_n511), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT28), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n531), .B1(new_n374), .B2(new_n314), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n533), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT28), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n540), .B(new_n544), .C1(new_n533), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n529), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n369), .A2(new_n417), .A3(KEYINPUT66), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n510), .B1(new_n314), .B2(new_n374), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n533), .B(new_n516), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n525), .A2(new_n528), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n516), .A2(new_n508), .A3(new_n518), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n532), .B2(new_n508), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n431), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n507), .B1(new_n538), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT32), .ZN(new_n558));
  INV_X1    g372(.A(new_n507), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n516), .B1(new_n547), .B2(new_n548), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n519), .B1(new_n560), .B2(KEYINPUT30), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n534), .B1(new_n561), .B2(new_n533), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT68), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n520), .A2(KEYINPUT68), .A3(new_n534), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT31), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n545), .A2(new_n529), .B1(new_n554), .B2(new_n537), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n559), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n558), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n545), .A2(new_n529), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n539), .B1(new_n553), .B2(new_n431), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n550), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n572), .A2(KEYINPUT29), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n532), .A2(new_n533), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT28), .B1(new_n576), .B2(new_n539), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n544), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n550), .A2(KEYINPUT29), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n214), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G472), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n506), .B1(new_n571), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n476), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  AOI21_X1  g398(.A(new_n502), .B1(new_n566), .B2(new_n567), .ZN(new_n585));
  INV_X1    g399(.A(G472), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n587), .A2(new_n506), .A3(new_n568), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT78), .B1(new_n410), .B2(new_n304), .ZN(new_n589));
  INV_X1    g403(.A(new_n304), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n402), .B(new_n590), .C1(new_n404), .C2(new_n409), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n588), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT92), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n403), .A2(new_n411), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n588), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n270), .B1(new_n298), .B2(new_n300), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT93), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n599), .A2(KEYINPUT93), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n213), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n211), .A2(KEYINPUT93), .A3(new_n599), .A4(new_n212), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(G478), .A3(new_n214), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n215), .A2(new_n216), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n598), .A2(new_n607), .A3(new_n279), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n465), .B1(new_n451), .B2(new_n463), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n451), .A2(new_n463), .A3(new_n465), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n608), .B(new_n473), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n597), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n473), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n224), .A2(new_n225), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n301), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n617), .B(new_n618), .C1(new_n610), .C2(new_n609), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n597), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT94), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT35), .B(G107), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NOR2_X1   g438(.A1(new_n587), .A2(new_n568), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n494), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n490), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n497), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n504), .B2(new_n505), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n476), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  AOI21_X1  g450(.A(new_n631), .B1(new_n571), .B2(new_n581), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n594), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT96), .B(G900), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n276), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n275), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n270), .B(new_n642), .C1(new_n298), .C2(new_n300), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n617), .B(new_n644), .C1(new_n610), .C2(new_n609), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n190), .ZN(G30));
  XNOR2_X1  g461(.A(new_n642), .B(KEYINPUT39), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n594), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT40), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n529), .B1(new_n576), .B2(new_n539), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n564), .A2(new_n565), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(G902), .B1(new_n652), .B2(KEYINPUT97), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(KEYINPUT97), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n571), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT98), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n472), .B(KEYINPUT38), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n631), .A2(new_n598), .A3(new_n617), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n414), .ZN(G45));
  AND3_X1   g476(.A1(new_n598), .A2(new_n607), .A3(new_n642), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(new_n473), .C1(new_n609), .C2(new_n610), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n247), .ZN(G48));
  INV_X1    g480(.A(new_n506), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n568), .A2(new_n569), .ZN(new_n668));
  AOI211_X1 g482(.A(KEYINPUT32), .B(new_n559), .C1(new_n566), .C2(new_n567), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n581), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n387), .A2(new_n370), .ZN(new_n671));
  OAI22_X1  g485(.A1(new_n671), .A2(new_n388), .B1(new_n394), .B2(new_n395), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n214), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G469), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n304), .A3(new_n398), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n612), .A2(new_n667), .A3(new_n670), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G15));
  NAND4_X1  g493(.A1(new_n620), .A2(new_n670), .A3(new_n667), .A4(new_n676), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  OAI21_X1  g495(.A(new_n473), .B1(new_n610), .B2(new_n609), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n675), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n670), .A3(new_n302), .A4(new_n630), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n578), .A2(new_n529), .B1(new_n554), .B2(new_n537), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n566), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n688), .B2(new_n507), .ZN(new_n689));
  AOI211_X1 g503(.A(KEYINPUT99), .B(new_n559), .C1(new_n566), .C2(new_n687), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n214), .B1(new_n538), .B2(new_n556), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(G472), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT100), .B1(new_n585), .B2(new_n586), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n691), .A2(new_n667), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n617), .B(new_n598), .C1(new_n610), .C2(new_n609), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n279), .A3(new_n676), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n199), .ZN(G24));
  NAND2_X1  g515(.A1(new_n694), .A2(new_n695), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n689), .A2(new_n690), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n630), .A3(new_n663), .A4(new_n683), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  NOR2_X1   g520(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n616), .B1(new_n469), .B2(new_n471), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n385), .A2(G469), .A3(new_n389), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n398), .A2(new_n399), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT101), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n398), .A2(new_n712), .A3(new_n399), .A4(new_n709), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n590), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n708), .A2(new_n667), .A3(new_n670), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n663), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n707), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n472), .A2(new_n473), .A3(new_n714), .ZN(new_n718));
  INV_X1    g532(.A(new_n707), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n582), .A3(new_n663), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  NOR3_X1   g536(.A1(new_n643), .A2(new_n224), .A3(new_n225), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n718), .A2(new_n582), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n405), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT103), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n726), .B1(new_n390), .B2(new_n391), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(G469), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n399), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n398), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n590), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n648), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n605), .A2(new_n606), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n598), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT43), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n626), .A2(new_n630), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n708), .B(KEYINPUT104), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n359), .ZN(G39));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n736), .B2(new_n590), .ZN(new_n750));
  OAI211_X1 g564(.A(KEYINPUT47), .B(new_n304), .C1(new_n734), .C2(new_n735), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n708), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n753), .A2(new_n667), .A3(new_n670), .A4(new_n716), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  NAND2_X1  g570(.A1(new_n674), .A2(new_n398), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT49), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT49), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n506), .A2(new_n474), .A3(new_n590), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n740), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n657), .A2(new_n658), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n658), .A2(new_n616), .A3(new_n676), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT110), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n741), .A2(new_n275), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n667), .A3(new_n704), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n766), .B1(KEYINPUT111), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n763), .A2(KEYINPUT110), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT50), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(KEYINPUT50), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n764), .A2(new_n768), .A3(new_n773), .A4(new_n769), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n674), .A2(new_n590), .A3(new_n398), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n750), .A2(new_n751), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n766), .A2(new_n745), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT113), .A4(new_n776), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n753), .A2(new_n675), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n765), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n784), .A2(new_n631), .A3(new_n703), .A4(new_n702), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n667), .A2(new_n657), .A3(new_n275), .A4(new_n783), .ZN(new_n786));
  INV_X1    g600(.A(new_n598), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n739), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n775), .A2(new_n782), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n777), .A2(new_n780), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n772), .A2(new_n796), .A3(new_n774), .A4(new_n790), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n793), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n786), .A2(new_n598), .A3(new_n607), .ZN(new_n799));
  INV_X1    g613(.A(new_n582), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n784), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n766), .A2(new_n682), .A3(new_n675), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n799), .A2(new_n803), .A3(new_n274), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n795), .A2(new_n798), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n684), .B1(new_n696), .B2(new_n699), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n677), .A2(new_n680), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n721), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n610), .A2(new_n609), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n470), .B1(new_n812), .B2(KEYINPUT85), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT105), .ZN(new_n814));
  INV_X1    g628(.A(new_n474), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n222), .A2(new_n223), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n787), .A2(new_n279), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n469), .A2(new_n471), .A3(new_n817), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT105), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n593), .A3(new_n596), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n813), .A2(new_n815), .A3(new_n608), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n593), .A2(new_n596), .A3(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n475), .B(new_n412), .C1(new_n632), .C2(new_n582), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n811), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n645), .ZN(new_n828));
  INV_X1    g642(.A(new_n664), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n637), .B(new_n594), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n630), .B1(new_n641), .B2(new_n640), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n656), .A2(new_n698), .A3(new_n714), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n705), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n830), .A2(new_n705), .A3(new_n835), .A4(new_n832), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n718), .A2(new_n630), .A3(new_n663), .A4(new_n704), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n643), .A2(new_n816), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n637), .A2(new_n594), .A3(new_n708), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n724), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT106), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n838), .A2(new_n724), .A3(KEYINPUT106), .A4(new_n840), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n827), .A2(new_n837), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT108), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT53), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT108), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n827), .A2(new_n837), .A3(new_n845), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(KEYINPUT108), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n807), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT109), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n834), .A2(KEYINPUT107), .A3(new_n836), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(new_n849), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n846), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n849), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n837), .A3(new_n827), .A4(new_n845), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n854), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n852), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n834), .A2(new_n836), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n843), .B2(new_n844), .ZN(new_n866));
  INV_X1    g680(.A(new_n852), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n827), .A3(new_n850), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT54), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n807), .B1(new_n858), .B2(new_n860), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT109), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n806), .B1(new_n863), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n762), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT115), .B(new_n762), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(G75));
  NAND2_X1  g692(.A1(new_n864), .A2(new_n868), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n214), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n466), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n449), .A2(new_n450), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n422), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT55), .Z(new_n885));
  AND3_X1   g699(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n881), .B2(new_n882), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n229), .A2(G952), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G51));
  OAI21_X1  g703(.A(KEYINPUT116), .B1(new_n879), .B2(new_n807), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n864), .A2(new_n868), .A3(new_n891), .A4(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n854), .A3(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n399), .B(KEYINPUT57), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n672), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n730), .B(KEYINPUT117), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n880), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n888), .B1(new_n896), .B2(new_n898), .ZN(G54));
  NAND3_X1  g713(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n900));
  INV_X1    g714(.A(new_n296), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n888), .ZN(G60));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n863), .A2(new_n871), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n604), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n906), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n888), .B1(new_n893), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT118), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(G63));
  XNOR2_X1  g731(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n208), .A2(new_n227), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n501), .B1(new_n879), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n864), .A2(new_n868), .A3(new_n628), .A4(new_n920), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n922), .B(new_n923), .C1(G952), .C2(new_n229), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n924), .B(new_n925), .Z(G66));
  INV_X1    g740(.A(new_n277), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n229), .B1(new_n927), .B2(new_n420), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n810), .A2(new_n822), .A3(new_n824), .A4(new_n825), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n229), .ZN(new_n930));
  INV_X1    g744(.A(G898), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n883), .B1(new_n931), .B2(G953), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n930), .B(new_n932), .ZN(G69));
  AOI21_X1  g747(.A(new_n229), .B1(G227), .B2(G900), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n284), .B(KEYINPUT121), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n553), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n787), .A2(new_n816), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n787), .B2(new_n739), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n649), .A2(new_n582), .A3(new_n708), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n738), .B2(new_n746), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(KEYINPUT123), .B(new_n939), .C1(new_n738), .C2(new_n746), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n830), .A2(new_n705), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n650), .B2(new_n660), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n947), .A2(KEYINPUT62), .B1(new_n752), .B2(new_n754), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT122), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n946), .A2(KEYINPUT122), .A3(new_n949), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n944), .B(new_n948), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n936), .B1(new_n952), .B2(new_n229), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(G900), .A2(G953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n800), .A2(new_n697), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n737), .A2(new_n648), .A3(new_n957), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT125), .Z(new_n959));
  INV_X1    g773(.A(new_n724), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n747), .A2(new_n960), .A3(new_n945), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n959), .A2(new_n721), .A3(new_n755), .A4(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n936), .B(new_n956), .C1(new_n962), .C2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n953), .B2(KEYINPUT124), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n934), .B1(new_n955), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n966));
  INV_X1    g780(.A(new_n934), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n966), .A2(new_n967), .A3(new_n954), .A4(new_n963), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  NOR2_X1   g785(.A1(new_n574), .A2(KEYINPUT126), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n574), .A2(KEYINPUT126), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n564), .A3(new_n565), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n861), .B(new_n971), .C1(new_n972), .C2(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT127), .Z(new_n976));
  OAI21_X1  g790(.A(new_n971), .B1(new_n952), .B2(new_n929), .ZN(new_n977));
  INV_X1    g791(.A(new_n573), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n550), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n971), .B1(new_n962), .B2(new_n929), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n550), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n888), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n976), .A2(new_n979), .A3(new_n982), .ZN(G57));
endmodule


