

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584;

  XOR2_X1 U325 ( .A(n310), .B(n309), .Z(n556) );
  INV_X1 U326 ( .A(KEYINPUT48), .ZN(n398) );
  XNOR2_X1 U327 ( .A(n399), .B(n398), .ZN(n532) );
  INV_X1 U328 ( .A(G190GAT), .ZN(n450) );
  XNOR2_X1 U329 ( .A(n450), .B(KEYINPUT58), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n294) );
  XNOR2_X1 U332 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n310) );
  XOR2_X1 U334 ( .A(G29GAT), .B(G43GAT), .Z(n296) );
  XNOR2_X1 U335 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U336 ( .A(n296), .B(n295), .ZN(n338) );
  XNOR2_X1 U337 ( .A(G99GAT), .B(G85GAT), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n297), .B(KEYINPUT75), .ZN(n363) );
  XNOR2_X1 U339 ( .A(n338), .B(n363), .ZN(n302) );
  XOR2_X1 U340 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n299) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U343 ( .A(n300), .B(KEYINPUT78), .Z(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .Z(n404) );
  XOR2_X1 U346 ( .A(n404), .B(G92GAT), .Z(n304) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n421) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(n421), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n308) );
  XNOR2_X1 U351 ( .A(G134GAT), .B(G218GAT), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U353 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n312) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT87), .ZN(n311) );
  XNOR2_X1 U355 ( .A(n312), .B(n311), .ZN(n429) );
  XOR2_X1 U356 ( .A(G85GAT), .B(n429), .Z(n314) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U359 ( .A(G29GAT), .B(n315), .ZN(n332) );
  XOR2_X1 U360 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n317) );
  XNOR2_X1 U361 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U363 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n319) );
  XNOR2_X1 U364 ( .A(G1GAT), .B(G57GAT), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U367 ( .A(G162GAT), .B(G155GAT), .Z(n323) );
  XNOR2_X1 U368 ( .A(G120GAT), .B(G148GAT), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U370 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U371 ( .A(n326), .B(KEYINPUT90), .Z(n330) );
  XOR2_X1 U372 ( .A(G127GAT), .B(KEYINPUT0), .Z(n328) );
  XNOR2_X1 U373 ( .A(G113GAT), .B(G134GAT), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n328), .B(n327), .ZN(n436) );
  XNOR2_X1 U375 ( .A(n436), .B(KEYINPUT91), .ZN(n329) );
  XNOR2_X1 U376 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U377 ( .A(n332), .B(n331), .ZN(n519) );
  XOR2_X1 U378 ( .A(G197GAT), .B(G22GAT), .Z(n334) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(G141GAT), .ZN(n333) );
  XNOR2_X1 U380 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U381 ( .A(n335), .B(G36GAT), .Z(n337) );
  XOR2_X1 U382 ( .A(G15GAT), .B(G1GAT), .Z(n383) );
  XNOR2_X1 U383 ( .A(n383), .B(G50GAT), .ZN(n336) );
  XNOR2_X1 U384 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U385 ( .A(G169GAT), .B(G8GAT), .Z(n407) );
  XOR2_X1 U386 ( .A(n338), .B(n407), .Z(n340) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U388 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U389 ( .A(n342), .B(n341), .Z(n350) );
  XOR2_X1 U390 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n344) );
  XNOR2_X1 U391 ( .A(KEYINPUT69), .B(KEYINPUT72), .ZN(n343) );
  XNOR2_X1 U392 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U393 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n346) );
  XNOR2_X1 U394 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U396 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U397 ( .A(n350), .B(n349), .ZN(n570) );
  XOR2_X1 U398 ( .A(G57GAT), .B(KEYINPUT13), .Z(n370) );
  XOR2_X1 U399 ( .A(G64GAT), .B(G92GAT), .Z(n352) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(G204GAT), .ZN(n351) );
  XNOR2_X1 U401 ( .A(n352), .B(n351), .ZN(n406) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U403 ( .A(n406), .B(n435), .ZN(n354) );
  AND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U406 ( .A(n370), .B(n355), .Z(n357) );
  XNOR2_X1 U407 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U409 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n359) );
  XNOR2_X1 U410 ( .A(KEYINPUT31), .B(KEYINPUT76), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U412 ( .A(n361), .B(n360), .Z(n365) );
  XNOR2_X1 U413 ( .A(G106GAT), .B(G78GAT), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n362), .B(G148GAT), .ZN(n428) );
  XNOR2_X1 U415 ( .A(n428), .B(n363), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n575) );
  XOR2_X1 U417 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n366) );
  XNOR2_X1 U418 ( .A(n575), .B(n366), .ZN(n559) );
  NOR2_X1 U419 ( .A1(n570), .A2(n559), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n367), .B(KEYINPUT46), .ZN(n389) );
  XOR2_X1 U421 ( .A(G78GAT), .B(G127GAT), .Z(n369) );
  XNOR2_X1 U422 ( .A(G183GAT), .B(G71GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U424 ( .A(n371), .B(n370), .Z(n373) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(G211GAT), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n387) );
  XOR2_X1 U427 ( .A(G22GAT), .B(G155GAT), .Z(n418) );
  XOR2_X1 U428 ( .A(KEYINPUT80), .B(n418), .Z(n375) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U431 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n377) );
  XNOR2_X1 U432 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U434 ( .A(n379), .B(n378), .Z(n385) );
  XOR2_X1 U435 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n381) );
  XNOR2_X1 U436 ( .A(G64GAT), .B(KEYINPUT84), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U440 ( .A(n387), .B(n386), .Z(n579) );
  NAND2_X1 U441 ( .A1(n556), .A2(n579), .ZN(n388) );
  NOR2_X1 U442 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n390), .B(KEYINPUT47), .ZN(n397) );
  XNOR2_X1 U444 ( .A(KEYINPUT36), .B(n556), .ZN(n582) );
  NOR2_X1 U445 ( .A1(n579), .A2(n582), .ZN(n391) );
  XNOR2_X1 U446 ( .A(KEYINPUT45), .B(n391), .ZN(n392) );
  NAND2_X1 U447 ( .A1(n392), .A2(n575), .ZN(n394) );
  INV_X1 U448 ( .A(KEYINPUT116), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  NAND2_X1 U450 ( .A1(n395), .A2(n570), .ZN(n396) );
  NAND2_X1 U451 ( .A1(n397), .A2(n396), .ZN(n399) );
  XOR2_X1 U452 ( .A(G211GAT), .B(KEYINPUT21), .Z(n401) );
  XNOR2_X1 U453 ( .A(G197GAT), .B(G218GAT), .ZN(n400) );
  XNOR2_X1 U454 ( .A(n401), .B(n400), .ZN(n420) );
  XOR2_X1 U455 ( .A(KEYINPUT94), .B(n420), .Z(n403) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U458 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U459 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U460 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U461 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n411) );
  XNOR2_X1 U462 ( .A(KEYINPUT86), .B(G183GAT), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U464 ( .A(KEYINPUT17), .B(n412), .Z(n446) );
  INV_X1 U465 ( .A(n446), .ZN(n413) );
  XOR2_X1 U466 ( .A(n414), .B(n413), .Z(n521) );
  INV_X1 U467 ( .A(n521), .ZN(n494) );
  XNOR2_X1 U468 ( .A(n494), .B(KEYINPUT122), .ZN(n415) );
  NOR2_X1 U469 ( .A1(n532), .A2(n415), .ZN(n416) );
  XOR2_X1 U470 ( .A(KEYINPUT54), .B(n416), .Z(n417) );
  NOR2_X1 U471 ( .A1(n519), .A2(n417), .ZN(n569) );
  XNOR2_X1 U472 ( .A(n418), .B(KEYINPUT24), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n419), .B(G204GAT), .ZN(n433) );
  XOR2_X1 U474 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U477 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n425) );
  XNOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U480 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n433), .B(n432), .ZN(n462) );
  NAND2_X1 U484 ( .A1(n569), .A2(n462), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n434), .B(KEYINPUT55), .ZN(n449) );
  XOR2_X1 U486 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U489 ( .A(G176GAT), .B(KEYINPUT85), .Z(n440) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U492 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U493 ( .A(G190GAT), .B(G99GAT), .Z(n444) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G15GAT), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U497 ( .A(n448), .B(n447), .ZN(n533) );
  NAND2_X1 U498 ( .A1(n449), .A2(n533), .ZN(n564) );
  NOR2_X1 U499 ( .A1(n556), .A2(n564), .ZN(n452) );
  INV_X1 U500 ( .A(n570), .ZN(n504) );
  NAND2_X1 U501 ( .A1(n575), .A2(n504), .ZN(n486) );
  INV_X1 U502 ( .A(n519), .ZN(n489) );
  NAND2_X1 U503 ( .A1(n533), .A2(n521), .ZN(n453) );
  NAND2_X1 U504 ( .A1(n462), .A2(n453), .ZN(n454) );
  XOR2_X1 U505 ( .A(KEYINPUT25), .B(n454), .Z(n458) );
  XOR2_X1 U506 ( .A(n494), .B(KEYINPUT27), .Z(n461) );
  NOR2_X1 U507 ( .A1(n533), .A2(n462), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT26), .B(n455), .Z(n456) );
  XNOR2_X1 U509 ( .A(KEYINPUT95), .B(n456), .ZN(n568) );
  NAND2_X1 U510 ( .A1(n461), .A2(n568), .ZN(n457) );
  NAND2_X1 U511 ( .A1(n458), .A2(n457), .ZN(n459) );
  NAND2_X1 U512 ( .A1(n489), .A2(n459), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT96), .ZN(n466) );
  NAND2_X1 U514 ( .A1(n519), .A2(n461), .ZN(n531) );
  NOR2_X1 U515 ( .A1(n533), .A2(n531), .ZN(n464) );
  XNOR2_X1 U516 ( .A(KEYINPUT66), .B(KEYINPUT28), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n463), .B(n462), .ZN(n535) );
  NAND2_X1 U518 ( .A1(n464), .A2(n535), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n482) );
  INV_X1 U520 ( .A(n579), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n556), .A2(n467), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT16), .B(n468), .Z(n469) );
  NAND2_X1 U523 ( .A1(n482), .A2(n469), .ZN(n470) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(n470), .Z(n506) );
  NOR2_X1 U525 ( .A1(n486), .A2(n506), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n471), .B(KEYINPUT98), .ZN(n479) );
  NAND2_X1 U527 ( .A1(n479), .A2(n519), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT34), .ZN(n473) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  XOR2_X1 U530 ( .A(G8GAT), .B(KEYINPUT99), .Z(n475) );
  NAND2_X1 U531 ( .A1(n479), .A2(n521), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n477) );
  NAND2_X1 U534 ( .A1(n533), .A2(n479), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(n478), .ZN(G1326GAT) );
  XOR2_X1 U537 ( .A(G22GAT), .B(KEYINPUT101), .Z(n481) );
  INV_X1 U538 ( .A(n535), .ZN(n526) );
  NAND2_X1 U539 ( .A1(n526), .A2(n479), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(G1327GAT) );
  NAND2_X1 U541 ( .A1(n579), .A2(n482), .ZN(n483) );
  NOR2_X1 U542 ( .A1(n582), .A2(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n518) );
  NOR2_X1 U545 ( .A1(n518), .A2(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT103), .B(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n502) );
  NOR2_X1 U548 ( .A1(n489), .A2(n502), .ZN(n493) );
  XOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n491) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n494), .A2(n502), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT106), .B(n495), .Z(n496) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n498) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(KEYINPUT108), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n501) );
  INV_X1 U559 ( .A(n533), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n502), .A2(n499), .ZN(n500) );
  XOR2_X1 U561 ( .A(n501), .B(n500), .Z(G1330GAT) );
  NOR2_X1 U562 ( .A1(n502), .A2(n535), .ZN(n503) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  NOR2_X1 U564 ( .A1(n559), .A2(n504), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT109), .ZN(n517) );
  NOR2_X1 U566 ( .A1(n506), .A2(n517), .ZN(n514) );
  NAND2_X1 U567 ( .A1(n514), .A2(n519), .ZN(n509) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT110), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(G64GAT), .B(KEYINPUT111), .Z(n511) );
  NAND2_X1 U572 ( .A1(n514), .A2(n521), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n514), .A2(n533), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U578 ( .A1(n514), .A2(n526), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n518), .A2(n517), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n519), .A2(n527), .ZN(n520) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  XOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT113), .Z(n523) );
  NAND2_X1 U584 ( .A1(n527), .A2(n521), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n527), .A2(n533), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n524), .B(KEYINPUT114), .ZN(n525) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n529) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n548) );
  NAND2_X1 U594 ( .A1(n533), .A2(n548), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n534), .B(KEYINPUT117), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X1 U597 ( .A1(n570), .A2(n543), .ZN(n537) );
  XOR2_X1 U598 ( .A(n537), .B(KEYINPUT118), .Z(n538) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n559), .A2(n543), .ZN(n540) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n579), .A2(n543), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(n541), .Z(n542) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  NOR2_X1 U606 ( .A1(n543), .A2(n556), .ZN(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n545) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT120), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n568), .ZN(n555) );
  NOR2_X1 U612 ( .A1(n570), .A2(n555), .ZN(n549) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U614 ( .A1(n555), .A2(n559), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n579), .A2(n555), .ZN(n554) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n554), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n570), .A2(n564), .ZN(n558) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n558), .Z(G1348GAT) );
  NOR2_X1 U625 ( .A1(n564), .A2(n559), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U630 ( .A1(n579), .A2(n564), .ZN(n565) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n581) );
  NOR2_X1 U636 ( .A1(n570), .A2(n581), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n581), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

