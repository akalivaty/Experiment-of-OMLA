

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U324 ( .A(n367), .B(n366), .ZN(n370) );
  XNOR2_X1 U325 ( .A(n398), .B(KEYINPUT47), .ZN(n399) );
  XNOR2_X1 U326 ( .A(n400), .B(n399), .ZN(n405) );
  XNOR2_X1 U327 ( .A(n365), .B(KEYINPUT68), .ZN(n366) );
  XNOR2_X1 U328 ( .A(n421), .B(n420), .ZN(n447) );
  XNOR2_X1 U329 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U330 ( .A(KEYINPUT36), .B(n546), .ZN(n584) );
  XNOR2_X1 U331 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U332 ( .A(n456), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT64), .B(G190GAT), .Z(n293) );
  XNOR2_X1 U335 ( .A(G15GAT), .B(G99GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U337 ( .A(n294), .B(G134GAT), .Z(n296) );
  XOR2_X1 U338 ( .A(G120GAT), .B(G71GAT), .Z(n355) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(n355), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n302) );
  XOR2_X1 U341 ( .A(G127GAT), .B(KEYINPUT0), .Z(n298) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n438) );
  XOR2_X1 U344 ( .A(G169GAT), .B(n438), .Z(n300) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U347 ( .A(n302), .B(n301), .Z(n312) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(G183GAT), .Z(n304) );
  XNOR2_X1 U349 ( .A(KEYINPUT17), .B(KEYINPUT84), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n305), .B(KEYINPUT18), .Z(n307) );
  XNOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT85), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n419) );
  XOR2_X1 U354 ( .A(G176GAT), .B(KEYINPUT81), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n419), .B(n310), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n533) );
  XOR2_X1 U359 ( .A(G50GAT), .B(G162GAT), .Z(n390) );
  XOR2_X1 U360 ( .A(G155GAT), .B(KEYINPUT2), .Z(n314) );
  XNOR2_X1 U361 ( .A(KEYINPUT87), .B(KEYINPUT3), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n434) );
  XOR2_X1 U363 ( .A(G211GAT), .B(KEYINPUT21), .Z(n316) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(G218GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n415) );
  XNOR2_X1 U366 ( .A(n434), .B(n415), .ZN(n321) );
  XOR2_X1 U367 ( .A(G78GAT), .B(G148GAT), .Z(n318) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n349) );
  XNOR2_X1 U370 ( .A(n349), .B(KEYINPUT86), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n319), .B(KEYINPUT22), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U373 ( .A(n322), .B(KEYINPUT24), .Z(n324) );
  XOR2_X1 U374 ( .A(G141GAT), .B(G22GAT), .Z(n361) );
  XNOR2_X1 U375 ( .A(n361), .B(KEYINPUT23), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U377 ( .A(n390), .B(n325), .Z(n327) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n470) );
  XOR2_X1 U380 ( .A(G64GAT), .B(G71GAT), .Z(n329) );
  XNOR2_X1 U381 ( .A(G183GAT), .B(G127GAT), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U383 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n331) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n344) );
  XOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT13), .Z(n352) );
  XOR2_X1 U388 ( .A(G78GAT), .B(G211GAT), .Z(n335) );
  XNOR2_X1 U389 ( .A(G22GAT), .B(G155GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U391 ( .A(n352), .B(n336), .Z(n338) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U394 ( .A(n339), .B(KEYINPUT78), .Z(n342) );
  XNOR2_X1 U395 ( .A(G15GAT), .B(G1GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n340), .B(KEYINPUT70), .ZN(n368) );
  XNOR2_X1 U397 ( .A(n368), .B(KEYINPUT77), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n579) );
  XOR2_X1 U400 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n346) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n347), .B(KEYINPUT33), .ZN(n351) );
  XNOR2_X1 U404 ( .A(G99GAT), .B(G85GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n348), .B(KEYINPUT71), .ZN(n379) );
  XNOR2_X1 U406 ( .A(n349), .B(n379), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n357) );
  XNOR2_X1 U409 ( .A(G176GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n354), .B(G64GAT), .ZN(n414) );
  XNOR2_X1 U411 ( .A(n355), .B(n414), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n479) );
  XOR2_X1 U413 ( .A(n479), .B(KEYINPUT41), .Z(n538) );
  XOR2_X1 U414 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n359) );
  XNOR2_X1 U415 ( .A(G197GAT), .B(G113GAT), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n364) );
  XOR2_X1 U417 ( .A(G36GAT), .B(G50GAT), .Z(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U419 ( .A(G169GAT), .B(G8GAT), .Z(n410) );
  XNOR2_X1 U420 ( .A(n362), .B(n410), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n367) );
  AND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XOR2_X1 U423 ( .A(n368), .B(KEYINPUT30), .Z(n369) );
  XOR2_X1 U424 ( .A(n370), .B(n369), .Z(n374) );
  XOR2_X1 U425 ( .A(KEYINPUT7), .B(KEYINPUT69), .Z(n372) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(G29GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U428 ( .A(KEYINPUT8), .B(n373), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n374), .B(n377), .ZN(n536) );
  NOR2_X1 U430 ( .A1(n538), .A2(n536), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n375), .B(KEYINPUT46), .ZN(n376) );
  NOR2_X1 U432 ( .A1(n579), .A2(n376), .ZN(n397) );
  INV_X1 U433 ( .A(n377), .ZN(n396) );
  INV_X1 U434 ( .A(KEYINPUT73), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n381) );
  NAND2_X1 U436 ( .A1(G232GAT), .A2(G233GAT), .ZN(n380) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n383) );
  XNOR2_X1 U438 ( .A(G36GAT), .B(G190GAT), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT76), .ZN(n407) );
  XNOR2_X1 U440 ( .A(n383), .B(n407), .ZN(n394) );
  XOR2_X1 U441 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n385) );
  XNOR2_X1 U442 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U444 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n387) );
  XNOR2_X1 U445 ( .A(G218GAT), .B(G106GAT), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n392) );
  XOR2_X1 U448 ( .A(G134GAT), .B(KEYINPUT75), .Z(n437) );
  XNOR2_X1 U449 ( .A(n390), .B(n437), .ZN(n391) );
  XOR2_X1 U450 ( .A(n396), .B(n395), .Z(n559) );
  INV_X1 U451 ( .A(n559), .ZN(n546) );
  NAND2_X1 U452 ( .A1(n397), .A2(n546), .ZN(n400) );
  XOR2_X1 U453 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n398) );
  INV_X1 U454 ( .A(n579), .ZN(n542) );
  NOR2_X1 U455 ( .A1(n584), .A2(n542), .ZN(n401) );
  XNOR2_X1 U456 ( .A(KEYINPUT45), .B(n401), .ZN(n402) );
  NAND2_X1 U457 ( .A1(n402), .A2(n479), .ZN(n403) );
  INV_X1 U458 ( .A(n536), .ZN(n569) );
  NOR2_X1 U459 ( .A1(n403), .A2(n569), .ZN(n404) );
  NOR2_X1 U460 ( .A1(n405), .A2(n404), .ZN(n406) );
  XOR2_X1 U461 ( .A(KEYINPUT48), .B(n406), .Z(n531) );
  XOR2_X1 U462 ( .A(n407), .B(KEYINPUT95), .Z(n409) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n410), .B(G204GAT), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n411), .B(KEYINPUT96), .ZN(n412) );
  XOR2_X1 U467 ( .A(n413), .B(n412), .Z(n417) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U470 ( .A(n419), .B(n418), .Z(n462) );
  NAND2_X1 U471 ( .A1(n531), .A2(n462), .ZN(n421) );
  XOR2_X1 U472 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n420) );
  XOR2_X1 U473 ( .A(G57GAT), .B(KEYINPUT5), .Z(n423) );
  XNOR2_X1 U474 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U476 ( .A(G85GAT), .B(G148GAT), .Z(n425) );
  XNOR2_X1 U477 ( .A(G141GAT), .B(G120GAT), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n446) );
  XOR2_X1 U480 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n429) );
  XNOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U483 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n431) );
  XNOR2_X1 U484 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U486 ( .A(n433), .B(n432), .Z(n444) );
  XOR2_X1 U487 ( .A(n434), .B(KEYINPUT1), .Z(n436) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n442) );
  XOR2_X1 U490 ( .A(n437), .B(G162GAT), .Z(n440) );
  XNOR2_X1 U491 ( .A(G29GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n446), .B(n445), .ZN(n519) );
  NAND2_X1 U496 ( .A1(n447), .A2(n519), .ZN(n567) );
  NOR2_X1 U497 ( .A1(n470), .A2(n567), .ZN(n448) );
  XNOR2_X1 U498 ( .A(KEYINPUT55), .B(n448), .ZN(n449) );
  NOR2_X1 U499 ( .A1(n533), .A2(n449), .ZN(n451) );
  INV_X1 U500 ( .A(KEYINPUT119), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n451), .B(n450), .ZN(n564) );
  INV_X1 U502 ( .A(n538), .ZN(n553) );
  NAND2_X1 U503 ( .A1(n564), .A2(n553), .ZN(n455) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT121), .Z(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  NAND2_X1 U508 ( .A1(n564), .A2(n559), .ZN(n458) );
  XOR2_X1 U509 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n456) );
  INV_X1 U510 ( .A(n519), .ZN(n468) );
  INV_X1 U511 ( .A(n462), .ZN(n522) );
  NOR2_X1 U512 ( .A1(n533), .A2(n522), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n470), .A2(n459), .ZN(n460) );
  XOR2_X1 U514 ( .A(n460), .B(KEYINPUT25), .Z(n461) );
  XNOR2_X1 U515 ( .A(KEYINPUT98), .B(n461), .ZN(n466) );
  XOR2_X1 U516 ( .A(n462), .B(KEYINPUT27), .Z(n472) );
  XOR2_X1 U517 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n464) );
  NAND2_X1 U518 ( .A1(n470), .A2(n533), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n568) );
  NOR2_X1 U520 ( .A1(n472), .A2(n568), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT99), .B(n469), .Z(n475) );
  XNOR2_X1 U524 ( .A(n470), .B(KEYINPUT66), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n471), .B(KEYINPUT28), .ZN(n489) );
  NOR2_X1 U526 ( .A1(n519), .A2(n472), .ZN(n530) );
  NAND2_X1 U527 ( .A1(n530), .A2(n533), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n489), .A2(n473), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n475), .A2(n474), .ZN(n492) );
  XOR2_X1 U530 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n477) );
  NAND2_X1 U531 ( .A1(n579), .A2(n546), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n477), .B(n476), .ZN(n478) );
  NOR2_X1 U533 ( .A1(n492), .A2(n478), .ZN(n507) );
  INV_X1 U534 ( .A(n479), .ZN(n575) );
  NOR2_X1 U535 ( .A1(n575), .A2(n536), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n480), .B(KEYINPUT72), .ZN(n496) );
  NAND2_X1 U537 ( .A1(n507), .A2(n496), .ZN(n490) );
  NOR2_X1 U538 ( .A1(n519), .A2(n490), .ZN(n481) );
  XOR2_X1 U539 ( .A(KEYINPUT34), .B(n481), .Z(n482) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n522), .A2(n490), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT100), .B(n483), .Z(n484) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n484), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n490), .A2(n533), .ZN(n488) );
  XOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n486) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT102), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  INV_X1 U549 ( .A(n489), .ZN(n534) );
  NOR2_X1 U550 ( .A1(n534), .A2(n490), .ZN(n491) );
  XOR2_X1 U551 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n495) );
  NOR2_X1 U554 ( .A1(n584), .A2(n492), .ZN(n493) );
  NAND2_X1 U555 ( .A1(n493), .A2(n542), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n518) );
  NAND2_X1 U557 ( .A1(n496), .A2(n518), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(KEYINPUT38), .ZN(n504) );
  NOR2_X1 U559 ( .A1(n519), .A2(n504), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n504), .A2(n522), .ZN(n500) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(n500), .Z(n501) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  NOR2_X1 U564 ( .A1(n533), .A2(n504), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(n502), .Z(n503) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U567 ( .A1(n504), .A2(n534), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  NOR2_X1 U570 ( .A1(n569), .A2(n538), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n517), .A2(n507), .ZN(n513) );
  NOR2_X1 U572 ( .A1(n519), .A2(n513), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n510), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n522), .A2(n513), .ZN(n511) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n533), .A2(n513), .ZN(n512) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n534), .A2(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n526) );
  NOR2_X1 U585 ( .A1(n519), .A2(n526), .ZN(n520) );
  XOR2_X1 U586 ( .A(G85GAT), .B(n520), .Z(n521) );
  XNOR2_X1 U587 ( .A(KEYINPUT108), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n526), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n533), .A2(n526), .ZN(n525) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n534), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U596 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT113), .B(n532), .Z(n550) );
  NOR2_X1 U599 ( .A1(n533), .A2(n550), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n545) );
  NOR2_X1 U601 ( .A1(n536), .A2(n545), .ZN(n537) );
  XOR2_X1 U602 ( .A(G113GAT), .B(n537), .Z(G1340GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n545), .ZN(n540) );
  XNOR2_X1 U604 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n542), .A2(n545), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U611 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n549), .Z(G1343GAT) );
  NOR2_X1 U614 ( .A1(n550), .A2(n568), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n551), .B(KEYINPUT116), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n560), .A2(n569), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U619 ( .A1(n560), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  XOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT117), .Z(n558) );
  NAND2_X1 U623 ( .A1(n579), .A2(n560), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n569), .A2(n564), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n579), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G183GAT), .B(n566), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n571) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n582) );
  NAND2_X1 U635 ( .A1(n582), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(n572), .B(KEYINPUT124), .Z(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  INV_X1 U647 ( .A(n582), .ZN(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

