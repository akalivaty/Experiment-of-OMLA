

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595;

  XNOR2_X1 U325 ( .A(n439), .B(n438), .ZN(n577) );
  NOR2_X1 U326 ( .A1(n483), .A2(n482), .ZN(n497) );
  XNOR2_X1 U327 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U328 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U329 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U330 ( .A(KEYINPUT113), .ZN(n434) );
  XOR2_X1 U331 ( .A(G29GAT), .B(G36GAT), .Z(n293) );
  XOR2_X1 U332 ( .A(n480), .B(n479), .Z(n294) );
  XNOR2_X1 U333 ( .A(n450), .B(n410), .ZN(n411) );
  INV_X1 U334 ( .A(KEYINPUT32), .ZN(n416) );
  INV_X1 U335 ( .A(n455), .ZN(n456) );
  INV_X1 U336 ( .A(KEYINPUT66), .ZN(n397) );
  XNOR2_X1 U337 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U338 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U339 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U340 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U341 ( .A(KEYINPUT36), .B(n491), .Z(n591) );
  XNOR2_X1 U342 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U343 ( .A(n465), .B(KEYINPUT122), .ZN(n571) );
  XOR2_X1 U344 ( .A(n463), .B(n462), .Z(n541) );
  XNOR2_X1 U345 ( .A(n488), .B(n487), .ZN(n516) );
  XNOR2_X1 U346 ( .A(n492), .B(G190GAT), .ZN(n493) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U348 ( .A(n494), .B(n493), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n442) );
  XOR2_X1 U351 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n296) );
  XNOR2_X1 U352 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U354 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n298) );
  XOR2_X1 U355 ( .A(G50GAT), .B(G162GAT), .Z(n396) );
  XOR2_X1 U356 ( .A(G22GAT), .B(G155GAT), .Z(n372) );
  XNOR2_X1 U357 ( .A(n396), .B(n372), .ZN(n297) );
  XNOR2_X1 U358 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U359 ( .A(n300), .B(n299), .Z(n302) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n309) );
  INV_X1 U362 ( .A(G148GAT), .ZN(n303) );
  NAND2_X1 U363 ( .A1(n303), .A2(G78GAT), .ZN(n306) );
  INV_X1 U364 ( .A(G78GAT), .ZN(n304) );
  NAND2_X1 U365 ( .A1(n304), .A2(G148GAT), .ZN(n305) );
  NAND2_X1 U366 ( .A1(n306), .A2(n305), .ZN(n308) );
  XNOR2_X1 U367 ( .A(G106GAT), .B(G204GAT), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n409) );
  XOR2_X1 U369 ( .A(n309), .B(n409), .Z(n316) );
  XNOR2_X1 U370 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n310), .B(KEYINPUT90), .ZN(n311) );
  XOR2_X1 U372 ( .A(n311), .B(KEYINPUT89), .Z(n313) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(G218GAT), .ZN(n312) );
  XOR2_X1 U374 ( .A(n313), .B(n312), .Z(n351) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n314), .B(KEYINPUT2), .ZN(n326) );
  XOR2_X1 U377 ( .A(n351), .B(n326), .Z(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n476) );
  XOR2_X1 U379 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n318) );
  XNOR2_X1 U380 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n330) );
  XOR2_X1 U382 ( .A(G57GAT), .B(G120GAT), .Z(n320) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(G127GAT), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U385 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n322) );
  XNOR2_X1 U386 ( .A(KEYINPUT95), .B(KEYINPUT97), .ZN(n321) );
  XNOR2_X1 U387 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U388 ( .A(n324), .B(n323), .Z(n328) );
  XNOR2_X1 U389 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n325), .B(KEYINPUT80), .ZN(n453) );
  XNOR2_X1 U391 ( .A(n453), .B(n326), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n338) );
  NAND2_X1 U394 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XOR2_X1 U395 ( .A(G85GAT), .B(G155GAT), .Z(n332) );
  XNOR2_X1 U396 ( .A(G148GAT), .B(G162GAT), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U398 ( .A(G29GAT), .B(G134GAT), .Z(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U401 ( .A(n338), .B(n337), .Z(n576) );
  AND2_X1 U402 ( .A1(n476), .A2(n576), .ZN(n440) );
  XOR2_X1 U403 ( .A(G183GAT), .B(KEYINPUT87), .Z(n340) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U406 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n342) );
  XNOR2_X1 U407 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U409 ( .A(n344), .B(n343), .Z(n463) );
  XOR2_X1 U410 ( .A(G92GAT), .B(G64GAT), .Z(n415) );
  XOR2_X1 U411 ( .A(G204GAT), .B(G176GAT), .Z(n346) );
  XNOR2_X1 U412 ( .A(G36GAT), .B(G8GAT), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U414 ( .A(n415), .B(n347), .Z(n349) );
  NAND2_X1 U415 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n463), .B(n350), .ZN(n353) );
  INV_X1 U418 ( .A(n351), .ZN(n352) );
  XOR2_X1 U419 ( .A(n353), .B(n352), .Z(n512) );
  XNOR2_X1 U420 ( .A(G1GAT), .B(KEYINPUT72), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n354), .B(G8GAT), .ZN(n384) );
  XOR2_X1 U422 ( .A(G50GAT), .B(n384), .Z(n356) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U425 ( .A(n357), .B(G43GAT), .Z(n365) );
  XOR2_X1 U426 ( .A(G113GAT), .B(G141GAT), .Z(n359) );
  XNOR2_X1 U427 ( .A(G197GAT), .B(G22GAT), .ZN(n358) );
  XNOR2_X1 U428 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U429 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n361) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(G15GAT), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U434 ( .A(n366), .B(KEYINPUT29), .Z(n369) );
  XNOR2_X1 U435 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n293), .B(n367), .ZN(n393) );
  XNOR2_X1 U437 ( .A(n393), .B(KEYINPUT30), .ZN(n368) );
  XOR2_X1 U438 ( .A(n369), .B(n368), .Z(n470) );
  INV_X1 U439 ( .A(n470), .ZN(n580) );
  XOR2_X1 U440 ( .A(KEYINPUT69), .B(KEYINPUT45), .Z(n404) );
  XOR2_X1 U441 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U444 ( .A(n372), .B(G78GAT), .Z(n374) );
  XOR2_X1 U445 ( .A(G15GAT), .B(G127GAT), .Z(n455) );
  XNOR2_X1 U446 ( .A(n455), .B(G211GAT), .ZN(n373) );
  XNOR2_X1 U447 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U448 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U449 ( .A1(G231GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U450 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U451 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n380) );
  XNOR2_X1 U452 ( .A(G183GAT), .B(G64GAT), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U454 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U455 ( .A(G71GAT), .B(G57GAT), .ZN(n383) );
  XNOR2_X1 U456 ( .A(n383), .B(KEYINPUT13), .ZN(n408) );
  XNOR2_X1 U457 ( .A(n384), .B(n408), .ZN(n385) );
  XNOR2_X1 U458 ( .A(n386), .B(n385), .ZN(n589) );
  XOR2_X1 U459 ( .A(G92GAT), .B(KEYINPUT9), .Z(n388) );
  NAND2_X1 U460 ( .A1(G232GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U461 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U462 ( .A(G106GAT), .B(n389), .Z(n402) );
  XOR2_X1 U463 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n391) );
  XNOR2_X1 U464 ( .A(G190GAT), .B(KEYINPUT68), .ZN(n390) );
  XNOR2_X1 U465 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U466 ( .A(G99GAT), .B(G85GAT), .Z(n407) );
  XOR2_X1 U467 ( .A(n392), .B(n407), .Z(n395) );
  XOR2_X1 U468 ( .A(G43GAT), .B(G134GAT), .Z(n454) );
  XNOR2_X1 U469 ( .A(n393), .B(n454), .ZN(n394) );
  XNOR2_X1 U470 ( .A(n395), .B(n394), .ZN(n400) );
  XNOR2_X1 U471 ( .A(G218GAT), .B(n396), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n402), .B(n401), .ZN(n491) );
  NAND2_X1 U473 ( .A1(n589), .A2(n591), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n422) );
  XOR2_X1 U475 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n406) );
  XNOR2_X1 U476 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n421) );
  XOR2_X1 U478 ( .A(n408), .B(n407), .Z(n414) );
  XNOR2_X1 U479 ( .A(n409), .B(KEYINPUT76), .ZN(n412) );
  XOR2_X1 U480 ( .A(G176GAT), .B(G120GAT), .Z(n450) );
  AND2_X1 U481 ( .A1(G230GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U482 ( .A(n414), .B(n413), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n415), .B(KEYINPUT75), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n426) );
  NOR2_X1 U485 ( .A1(n422), .A2(n426), .ZN(n423) );
  XOR2_X1 U486 ( .A(KEYINPUT112), .B(n423), .Z(n424) );
  NOR2_X1 U487 ( .A1(n580), .A2(n424), .ZN(n433) );
  XNOR2_X1 U488 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n425) );
  XOR2_X1 U489 ( .A(n426), .B(n425), .Z(n570) );
  INV_X1 U490 ( .A(n570), .ZN(n545) );
  NAND2_X1 U491 ( .A1(n545), .A2(n580), .ZN(n428) );
  XOR2_X1 U492 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U494 ( .A(n589), .B(KEYINPUT110), .Z(n549) );
  INV_X1 U495 ( .A(n491), .ZN(n567) );
  AND2_X1 U496 ( .A1(n549), .A2(n491), .ZN(n429) );
  AND2_X1 U497 ( .A1(n430), .A2(n429), .ZN(n431) );
  XOR2_X1 U498 ( .A(n431), .B(KEYINPUT47), .Z(n432) );
  NOR2_X1 U499 ( .A1(n433), .A2(n432), .ZN(n437) );
  XOR2_X1 U500 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n435) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n556) );
  NAND2_X1 U502 ( .A1(n512), .A2(n556), .ZN(n439) );
  XNOR2_X1 U503 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n438) );
  NAND2_X1 U504 ( .A1(n440), .A2(n577), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n443), .B(KEYINPUT120), .ZN(n464) );
  XOR2_X1 U507 ( .A(KEYINPUT67), .B(KEYINPUT81), .Z(n445) );
  NAND2_X1 U508 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U510 ( .A(KEYINPUT20), .B(n446), .ZN(n461) );
  XOR2_X1 U511 ( .A(KEYINPUT82), .B(KEYINPUT85), .Z(n448) );
  XNOR2_X1 U512 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U514 ( .A(n449), .B(G71GAT), .Z(n452) );
  XNOR2_X1 U515 ( .A(n450), .B(G99GAT), .ZN(n451) );
  XNOR2_X1 U516 ( .A(n452), .B(n451), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n454), .B(n453), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U519 ( .A(n541), .ZN(n503) );
  NAND2_X1 U520 ( .A1(n464), .A2(n503), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n571), .A2(n470), .ZN(n467) );
  INV_X1 U522 ( .A(G169GAT), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n467), .B(n466), .ZN(G1348GAT) );
  NOR2_X1 U524 ( .A1(n549), .A2(n571), .ZN(n469) );
  INV_X1 U525 ( .A(G183GAT), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(G1350GAT) );
  XOR2_X1 U527 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n488) );
  NOR2_X1 U528 ( .A1(n470), .A2(n426), .ZN(n498) );
  XNOR2_X1 U529 ( .A(n476), .B(KEYINPUT28), .ZN(n537) );
  INV_X1 U530 ( .A(n537), .ZN(n515) );
  INV_X1 U531 ( .A(n512), .ZN(n532) );
  XNOR2_X1 U532 ( .A(KEYINPUT27), .B(n532), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n515), .A2(n474), .ZN(n471) );
  INV_X1 U534 ( .A(n576), .ZN(n509) );
  NAND2_X1 U535 ( .A1(n471), .A2(n509), .ZN(n540) );
  XOR2_X1 U536 ( .A(KEYINPUT88), .B(n541), .Z(n472) );
  NOR2_X1 U537 ( .A1(n540), .A2(n472), .ZN(n483) );
  NOR2_X1 U538 ( .A1(n476), .A2(n503), .ZN(n473) );
  XOR2_X1 U539 ( .A(KEYINPUT26), .B(n473), .Z(n578) );
  NOR2_X1 U540 ( .A1(n578), .A2(n474), .ZN(n557) );
  NAND2_X1 U541 ( .A1(n503), .A2(n512), .ZN(n475) );
  XNOR2_X1 U542 ( .A(KEYINPUT98), .B(n475), .ZN(n477) );
  NAND2_X1 U543 ( .A1(n477), .A2(n476), .ZN(n480) );
  XNOR2_X1 U544 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n478) );
  XNOR2_X1 U545 ( .A(n478), .B(KEYINPUT25), .ZN(n479) );
  NOR2_X1 U546 ( .A1(n557), .A2(n294), .ZN(n481) );
  NOR2_X1 U547 ( .A1(n481), .A2(n509), .ZN(n482) );
  NOR2_X1 U548 ( .A1(n589), .A2(n497), .ZN(n484) );
  XOR2_X1 U549 ( .A(KEYINPUT103), .B(n484), .Z(n485) );
  NAND2_X1 U550 ( .A1(n591), .A2(n485), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n486), .B(KEYINPUT37), .ZN(n530) );
  NAND2_X1 U552 ( .A1(n498), .A2(n530), .ZN(n487) );
  NAND2_X1 U553 ( .A1(n503), .A2(n516), .ZN(n490) );
  NOR2_X1 U554 ( .A1(n571), .A2(n491), .ZN(n494) );
  INV_X1 U555 ( .A(KEYINPUT58), .ZN(n492) );
  NAND2_X1 U556 ( .A1(n589), .A2(n491), .ZN(n495) );
  XNOR2_X1 U557 ( .A(KEYINPUT16), .B(n495), .ZN(n496) );
  NOR2_X1 U558 ( .A1(n497), .A2(n496), .ZN(n519) );
  NAND2_X1 U559 ( .A1(n519), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT101), .ZN(n507) );
  NAND2_X1 U561 ( .A1(n509), .A2(n507), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U564 ( .A1(n512), .A2(n507), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U567 ( .A1(n507), .A2(n503), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G15GAT), .B(n506), .ZN(G1326GAT) );
  NAND2_X1 U570 ( .A1(n507), .A2(n515), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .Z(n511) );
  NAND2_X1 U573 ( .A1(n516), .A2(n509), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  XOR2_X1 U575 ( .A(G36GAT), .B(KEYINPUT105), .Z(n514) );
  NAND2_X1 U576 ( .A1(n516), .A2(n512), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1329GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n517), .B(KEYINPUT106), .ZN(n518) );
  XNOR2_X1 U580 ( .A(G50GAT), .B(n518), .ZN(G1331GAT) );
  NOR2_X1 U581 ( .A1(n580), .A2(n570), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n529), .A2(n519), .ZN(n525) );
  NOR2_X1 U583 ( .A1(n576), .A2(n525), .ZN(n521) );
  XNOR2_X1 U584 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n522), .ZN(G1332GAT) );
  NOR2_X1 U587 ( .A1(n532), .A2(n525), .ZN(n523) );
  XOR2_X1 U588 ( .A(G64GAT), .B(n523), .Z(G1333GAT) );
  NOR2_X1 U589 ( .A1(n541), .A2(n525), .ZN(n524) );
  XOR2_X1 U590 ( .A(G71GAT), .B(n524), .Z(G1334GAT) );
  NOR2_X1 U591 ( .A1(n537), .A2(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G78GAT), .B(n528), .ZN(G1335GAT) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U596 ( .A1(n576), .A2(n536), .ZN(n531) );
  XOR2_X1 U597 ( .A(G85GAT), .B(n531), .Z(G1336GAT) );
  NOR2_X1 U598 ( .A1(n532), .A2(n536), .ZN(n533) );
  XOR2_X1 U599 ( .A(G92GAT), .B(n533), .Z(G1337GAT) );
  NOR2_X1 U600 ( .A1(n541), .A2(n536), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1338GAT) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U604 ( .A(KEYINPUT44), .B(n538), .Z(n539) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n556), .A2(n542), .ZN(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT114), .B(n543), .ZN(n548) );
  INV_X1 U609 ( .A(n548), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n553), .A2(n580), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U613 ( .A1(n553), .A2(n545), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  XNOR2_X1 U615 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U620 ( .A1(n567), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n576), .A2(n558), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n568), .A2(n580), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT116), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n562) );
  NAND2_X1 U628 ( .A1(n568), .A2(n545), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT117), .Z(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n589), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(KEYINPUT118), .ZN(n566) );
  XNOR2_X1 U634 ( .A(G155GAT), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n573) );
  XNOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n579) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n592) );
  AND2_X1 U644 ( .A1(n580), .A2(n592), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n582) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(KEYINPUT124), .B(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U651 ( .A1(n592), .A2(n426), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G204GAT), .B(n588), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n592), .A2(n589), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n594) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

