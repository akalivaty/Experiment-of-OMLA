//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT67), .Z(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n215), .A2(G50), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OR3_X1    g0020(.A1(new_n206), .A2(KEYINPUT65), .A3(G13), .ZN(new_n221));
  OAI21_X1  g0021(.A(KEYINPUT65), .B1(new_n206), .B2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT0), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n225), .B2(new_n224), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n214), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n232), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G97), .B(G107), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  OR2_X1    g0044(.A1(KEYINPUT8), .A2(G58), .ZN(new_n245));
  NAND2_X1  g0045(.A1(KEYINPUT8), .A2(G58), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n248), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(KEYINPUT15), .B(G87), .Z(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n259), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G77), .ZN(new_n266));
  INV_X1    g0066(.A(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G13), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n260), .B(new_n266), .C1(G77), .C2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT69), .B1(new_n270), .B2(new_n258), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n218), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT70), .ZN(new_n278));
  INV_X1    g0078(.A(new_n276), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n271), .B2(new_n274), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n278), .A2(G244), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  AOI211_X1 g0084(.A(new_n284), .B(new_n276), .C1(new_n271), .C2(new_n274), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n270), .A2(new_n258), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G232), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(G238), .A3(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G107), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(new_n290), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n289), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n296), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n287), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n269), .B1(new_n299), .B2(G200), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n287), .A2(G190), .A3(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT72), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n287), .A2(new_n308), .A3(new_n298), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n269), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT73), .Z(new_n312));
  NAND3_X1  g0112(.A1(new_n278), .A2(G238), .A3(new_n282), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n290), .A2(G232), .A3(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n290), .A2(G226), .A3(new_n291), .ZN(new_n315));
  INV_X1    g0115(.A(G97), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n314), .B(new_n315), .C1(new_n251), .C2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n285), .B1(new_n317), .B2(new_n288), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n313), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n313), .B2(new_n318), .ZN(new_n322));
  OAI21_X1  g0122(.A(G169), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT14), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT14), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n325), .B(G169), .C1(new_n321), .C2(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(new_n322), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G179), .A3(new_n320), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G13), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n263), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G68), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT12), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n252), .A2(G77), .B1(G20), .B2(new_n332), .ZN(new_n335));
  INV_X1    g0135(.A(G50), .ZN(new_n336));
  INV_X1    g0136(.A(new_n249), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n334), .B(new_n339), .C1(new_n332), .C2(new_n264), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT11), .B1(new_n338), .B2(new_n259), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n329), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n327), .A2(G190), .A3(new_n320), .ZN(new_n346));
  OAI21_X1  g0146(.A(G200), .B1(new_n321), .B2(new_n322), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n346), .A2(new_n347), .A3(new_n342), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G20), .ZN(new_n350));
  INV_X1    g0150(.A(new_n201), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n202), .ZN(new_n352));
  INV_X1    g0152(.A(G150), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n247), .A2(new_n253), .B1(new_n353), .B2(new_n337), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n259), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n268), .A2(G50), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n265), .B2(G50), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n278), .A2(G226), .A3(new_n282), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n290), .A2(G223), .A3(G1698), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(new_n290), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n285), .B1(new_n364), .B2(new_n288), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(G179), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n359), .B(new_n367), .C1(new_n306), .C2(new_n366), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n358), .B(KEYINPUT9), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(G200), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n366), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n370), .B2(KEYINPUT74), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n374), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n312), .A2(new_n349), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G33), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n379), .A2(new_n381), .A3(G226), .A4(G1698), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT80), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n290), .A2(new_n384), .A3(G226), .A4(G1698), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n290), .A2(G223), .A3(new_n291), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n383), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n288), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n284), .B1(new_n271), .B2(new_n274), .ZN(new_n390));
  AOI22_X1  g0190(.A1(G232), .A2(new_n280), .B1(new_n390), .B2(new_n279), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G169), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n308), .B2(new_n392), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n249), .ZN(new_n397));
  AOI21_X1  g0197(.A(G20), .B1(new_n379), .B2(new_n381), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n401));
  NOR2_X1   g0201(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n403), .A2(new_n290), .A3(G20), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT16), .B(new_n397), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n259), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT76), .B1(new_n398), .B2(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n409), .C1(new_n290), .C2(G20), .ZN(new_n410));
  OR3_X1    g0210(.A1(new_n380), .A2(KEYINPUT77), .A3(G33), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n381), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n399), .A2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n407), .A2(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n397), .B1(new_n415), .B2(new_n332), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n406), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n247), .A2(new_n267), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT78), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n259), .B(new_n331), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n421), .A2(new_n423), .B1(new_n331), .B2(new_n247), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT79), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n405), .A2(new_n259), .ZN(new_n427));
  INV_X1    g0227(.A(new_n397), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n413), .A2(new_n414), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n380), .A2(G33), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n350), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n408), .B1(new_n432), .B2(new_n409), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n398), .A2(KEYINPUT76), .A3(new_n403), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n428), .B1(new_n435), .B2(G68), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n427), .B1(new_n436), .B2(KEYINPUT16), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n424), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n395), .B1(new_n426), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n418), .A2(new_n425), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT81), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n389), .A2(G190), .A3(new_n391), .ZN(new_n446));
  INV_X1    g0246(.A(G200), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n389), .B2(new_n391), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT17), .A4(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n437), .A3(new_n445), .A4(new_n424), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n450), .B(new_n453), .C1(new_n440), .C2(new_n441), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n443), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n378), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT25), .B1(new_n268), .B2(G107), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT25), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n331), .A2(new_n460), .A3(new_n294), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n262), .A2(G33), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n268), .A2(new_n261), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n459), .B(new_n461), .C1(new_n463), .C2(new_n294), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT94), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n350), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n294), .A2(KEYINPUT23), .A3(G20), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n468), .A2(new_n469), .B1(new_n252), .B2(G116), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT92), .B(KEYINPUT22), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n290), .A2(new_n472), .A3(new_n350), .A4(G87), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT93), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n379), .A2(new_n381), .A3(new_n350), .A4(G87), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n473), .A2(new_n474), .B1(KEYINPUT22), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g0276(.A(KEYINPUT92), .B(KEYINPUT22), .Z(new_n477));
  OR3_X1    g0277(.A1(new_n475), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n471), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n259), .B1(new_n479), .B2(KEYINPUT24), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n473), .A2(new_n474), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n470), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n466), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n379), .A2(new_n381), .A3(G250), .A4(new_n291), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT95), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT95), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n290), .A2(new_n491), .A3(G250), .A4(new_n291), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G294), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n379), .A2(new_n381), .A3(G257), .A4(G1698), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT96), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n494), .A2(new_n493), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT96), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(new_n492), .A4(new_n490), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n288), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  INV_X1    g0301(.A(G41), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT5), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(KEYINPUT84), .B2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(G45), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G1), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n390), .A2(new_n279), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n262), .A2(G45), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n501), .A2(new_n502), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(new_n503), .B1(new_n271), .B2(new_n274), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G264), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n500), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n306), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n500), .A2(new_n308), .A3(new_n510), .A4(new_n515), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n488), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n379), .A2(new_n381), .A3(G257), .A4(new_n291), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n379), .A2(new_n381), .A3(G264), .A4(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(new_n290), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n288), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n275), .A2(G270), .A3(new_n508), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n510), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT90), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT90), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n524), .A2(new_n510), .A3(new_n528), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n350), .C1(G33), .C2(new_n316), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n259), .C1(new_n350), .C2(G116), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n268), .A2(G116), .ZN(new_n536));
  INV_X1    g0336(.A(new_n463), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(G116), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n306), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n530), .B(new_n539), .C1(KEYINPUT91), .C2(KEYINPUT21), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n533), .B(KEYINPUT20), .ZN(new_n541));
  INV_X1    g0341(.A(new_n536), .ZN(new_n542));
  INV_X1    g0342(.A(G116), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n463), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n545), .A2(new_n308), .A3(new_n526), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n285), .A2(new_n509), .B1(new_n514), .B2(G270), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n528), .B1(new_n547), .B2(new_n524), .ZN(new_n548));
  INV_X1    g0348(.A(new_n529), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n539), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n519), .A2(new_n540), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n268), .A2(G97), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n463), .B2(new_n316), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n242), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n294), .A2(G97), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(G20), .B1(G77), .B2(new_n249), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n415), .B2(new_n294), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n556), .B1(new_n562), .B2(new_n259), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n258), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n272), .B1(new_n218), .B2(new_n273), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n508), .B(G257), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT85), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n275), .A2(KEYINPUT85), .A3(G257), .A4(new_n508), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n569), .B1(new_n285), .B2(new_n509), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n379), .A2(new_n381), .A3(G244), .A4(new_n291), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT4), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n290), .A2(new_n573), .A3(G244), .A4(new_n291), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n379), .A2(new_n381), .A3(G250), .A4(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n531), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(KEYINPUT83), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n288), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT83), .B1(new_n575), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n570), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G169), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n575), .A2(new_n578), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n288), .A3(new_n579), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G179), .A3(new_n570), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n563), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n556), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n559), .A2(new_n557), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n557), .B2(new_n242), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n592), .A2(new_n350), .B1(new_n363), .B2(new_n337), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n435), .B2(G107), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n590), .B1(new_n594), .B2(new_n261), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n563), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n582), .A2(new_n447), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n570), .B(new_n371), .C1(new_n580), .C2(new_n581), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n589), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n516), .A2(G200), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n261), .B1(new_n485), .B2(new_n486), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n486), .B2(new_n485), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n500), .A2(G190), .A3(new_n510), .A4(new_n515), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n604), .A2(new_n606), .A3(new_n466), .A4(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n527), .A2(G190), .A3(new_n529), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n545), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n447), .B1(new_n527), .B2(new_n529), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n613));
  OR2_X1    g0413(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n614));
  AND2_X1   g0414(.A1(G33), .A2(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n613), .B1(new_n617), .B2(new_n350), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n379), .A2(new_n381), .A3(new_n350), .A4(G68), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n350), .A2(G33), .A3(G97), .ZN(new_n620));
  INV_X1    g0420(.A(new_n616), .ZN(new_n621));
  NOR2_X1   g0421(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n259), .B1(new_n618), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n255), .A2(new_n331), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT89), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(KEYINPUT89), .A3(new_n626), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n628), .A2(new_n629), .B1(new_n254), .B2(new_n537), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n379), .A2(new_n381), .A3(G244), .A4(G1698), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n379), .A2(new_n381), .A3(G238), .A4(new_n291), .ZN(new_n632));
  NAND2_X1  g0432(.A1(G33), .A2(G116), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT87), .B1(new_n506), .B2(G1), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n262), .A3(G45), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n635), .A2(new_n637), .A3(G250), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n634), .A2(new_n288), .B1(new_n275), .B2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(G274), .B(new_n507), .C1(new_n564), .C2(new_n565), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(KEYINPUT86), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT86), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n390), .B2(new_n507), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n306), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n639), .B(new_n308), .C1(new_n641), .C2(new_n643), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n639), .B(G190), .C1(new_n641), .C2(new_n643), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n537), .A2(G87), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n625), .A2(KEYINPUT89), .A3(new_n626), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n627), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n644), .A2(G200), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n630), .A2(new_n647), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n612), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n553), .A2(new_n603), .A3(new_n608), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n458), .A2(new_n656), .ZN(G372));
  NAND2_X1  g0457(.A1(new_n437), .A2(new_n424), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n394), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n441), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(KEYINPUT18), .A3(new_n394), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n310), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n345), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n453), .A2(new_n450), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(new_n348), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n375), .A2(new_n376), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n368), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n646), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n640), .A2(KEYINPUT86), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n390), .A2(new_n642), .A3(new_n507), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(G169), .B1(new_n673), .B2(new_n639), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n650), .A2(new_n627), .B1(new_n255), .B2(new_n463), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI211_X1 g0477(.A(KEYINPUT97), .B(new_n447), .C1(new_n673), .C2(new_n639), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT97), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n644), .B2(G200), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n651), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n681), .A2(new_n682), .B1(new_n676), .B2(new_n675), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n562), .A2(new_n259), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n597), .B1(new_n684), .B2(new_n590), .ZN(new_n685));
  AOI211_X1 g0485(.A(KEYINPUT82), .B(new_n556), .C1(new_n562), .C2(new_n259), .ZN(new_n686));
  INV_X1    g0486(.A(new_n601), .ZN(new_n687));
  AOI21_X1  g0487(.A(G200), .B1(new_n587), .B2(new_n570), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n583), .A2(new_n588), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n595), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n683), .A2(new_n689), .A3(new_n691), .A4(new_n608), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n677), .B1(new_n692), .B2(new_n553), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT26), .B1(new_n691), .B2(new_n654), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n685), .A2(new_n686), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n683), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n694), .B1(new_n696), .B2(KEYINPUT26), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n669), .B1(new_n458), .B2(new_n698), .ZN(G369));
  NOR2_X1   g0499(.A1(new_n330), .A2(G20), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n262), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g0504(.A(KEYINPUT98), .B(G343), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n519), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n552), .A2(new_n540), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n707), .ZN(new_n710));
  AND4_X1   g0510(.A1(new_n466), .A2(new_n604), .A3(new_n606), .A4(new_n607), .ZN(new_n711));
  INV_X1    g0511(.A(new_n707), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n606), .B2(new_n466), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n519), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n708), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n545), .A2(new_n712), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT99), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT99), .ZN(new_n720));
  INV_X1    g0520(.A(new_n611), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n545), .A3(new_n609), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n709), .A2(new_n722), .A3(new_n717), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  INV_X1    g0525(.A(new_n708), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n714), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n715), .B1(new_n725), .B2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n223), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n613), .A2(new_n543), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n730), .A2(new_n262), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n217), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(new_n730), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT28), .Z(new_n735));
  INV_X1    g0535(.A(KEYINPUT100), .ZN(new_n736));
  INV_X1    g0536(.A(new_n644), .ZN(new_n737));
  AND4_X1   g0537(.A1(G179), .A2(new_n524), .A3(new_n510), .A4(new_n525), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(new_n515), .A4(new_n500), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n736), .B1(new_n739), .B2(new_n582), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n736), .B(new_n742), .C1(new_n739), .C2(new_n582), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n737), .A2(G179), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n516), .A3(new_n530), .A4(new_n582), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT31), .B1(new_n656), .B2(new_n707), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n707), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G330), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT101), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT101), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n682), .A2(new_n652), .B1(new_n675), .B2(new_n676), .ZN(new_n755));
  AND4_X1   g0555(.A1(new_n691), .A2(new_n689), .A3(new_n755), .A4(new_n722), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(new_n553), .A3(new_n608), .A4(new_n712), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(KEYINPUT31), .B1(new_n707), .B2(new_n746), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n754), .B(G330), .C1(new_n758), .C2(new_n748), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n696), .A2(KEYINPUT26), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n755), .A2(new_n589), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(KEYINPUT26), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n712), .B1(new_n764), .B2(new_n693), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n765), .A2(KEYINPUT29), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT29), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n698), .A2(new_n707), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n735), .B1(new_n771), .B2(G1), .ZN(G364));
  INV_X1    g0572(.A(new_n730), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n262), .B1(new_n700), .B2(G45), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n724), .B2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n724), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n258), .B1(G20), .B2(new_n306), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n350), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n447), .A2(G179), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G283), .A2(new_n784), .B1(new_n787), .B2(G329), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT104), .Z(new_n789));
  NOR2_X1   g0589(.A1(new_n308), .A2(new_n447), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n781), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n350), .A2(new_n371), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n782), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n792), .A2(new_n793), .B1(new_n796), .B2(G303), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n781), .A2(G179), .A3(new_n447), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n350), .A2(new_n308), .A3(new_n371), .A4(G200), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(G311), .B1(new_n800), .B2(G322), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n379), .A2(new_n381), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n794), .A2(new_n790), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n371), .A2(G179), .A3(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n350), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n805), .B1(G294), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n789), .A2(new_n797), .A3(new_n801), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n796), .A2(G87), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n332), .B2(new_n791), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G77), .B2(new_n799), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n783), .A2(new_n294), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n290), .B1(new_n803), .B2(new_n336), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G58), .C2(new_n800), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n808), .A2(G97), .ZN(new_n817));
  INV_X1    g0617(.A(G159), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n786), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT32), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n813), .A2(new_n816), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n780), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n330), .A2(new_n251), .A3(KEYINPUT103), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT103), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(G13), .B2(G33), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G20), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n779), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n729), .A2(new_n802), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(G355), .B1(new_n543), .B2(new_n729), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n240), .A2(G45), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n729), .A2(new_n290), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n506), .B2(new_n733), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n832), .B1(new_n835), .B2(KEYINPUT102), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n835), .A2(KEYINPUT102), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n775), .B(new_n822), .C1(new_n829), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n828), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n724), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n778), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NOR2_X1   g0643(.A1(new_n826), .A2(new_n779), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT105), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n791), .A2(new_n353), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n803), .A2(new_n848), .B1(new_n798), .B2(new_n818), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(G143), .C2(new_n800), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n290), .B1(new_n795), .B2(new_n336), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n783), .A2(new_n332), .B1(new_n786), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(G58), .C2(new_n808), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(G311), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n798), .A2(new_n543), .B1(new_n786), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n784), .A2(G87), .ZN(new_n860));
  INV_X1    g0660(.A(new_n803), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n859), .B(new_n860), .C1(G303), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n802), .B1(new_n795), .B2(new_n294), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT106), .Z(new_n864));
  AOI22_X1  g0664(.A1(G283), .A2(new_n792), .B1(new_n800), .B2(G294), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n817), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n857), .A2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n776), .B1(G77), .B2(new_n846), .C1(new_n867), .C2(new_n780), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n269), .A2(new_n707), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n663), .B1(new_n305), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n310), .A2(new_n707), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n868), .B1(new_n873), .B2(new_n826), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n761), .A2(new_n873), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n753), .B2(new_n759), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n768), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n776), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n768), .A3(new_n877), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(G384));
  NOR2_X1   g0682(.A1(new_n700), .A2(new_n262), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n397), .B1(new_n400), .B2(new_n404), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n885), .A2(new_n417), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n424), .B1(new_n886), .B2(new_n406), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT108), .ZN(new_n888));
  INV_X1    g0688(.A(new_n704), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT108), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(new_n424), .C1(new_n886), .C2(new_n406), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n426), .A2(new_n439), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n441), .B1(new_n893), .B2(new_n394), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n665), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n892), .B1(new_n895), .B2(new_n442), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n444), .A2(new_n449), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n440), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n704), .B1(new_n426), .B2(new_n439), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n888), .A2(new_n394), .A3(new_n891), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n892), .A2(new_n903), .A3(new_n897), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n900), .A2(new_n902), .B1(new_n904), .B2(KEYINPUT37), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n884), .B1(new_n896), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n892), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n443), .B2(new_n454), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n893), .A2(new_n394), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n902), .A2(new_n909), .A3(new_n898), .A4(new_n897), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(KEYINPUT109), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n342), .A2(new_n712), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n915), .B(new_n348), .C1(new_n329), .C2(new_n343), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n344), .A2(new_n712), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n872), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n689), .A2(new_n755), .A3(new_n691), .A4(new_n722), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n519), .A2(new_n552), .A3(new_n540), .ZN(new_n920));
  NOR4_X1   g0720(.A1(new_n919), .A2(new_n920), .A3(new_n711), .A4(new_n707), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT31), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n750), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT112), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n746), .A2(new_n925), .A3(KEYINPUT31), .A4(new_n707), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n918), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT109), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n908), .A2(new_n912), .A3(new_n929), .A4(KEYINPUT38), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n914), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n932), .B(new_n918), .C1(new_n923), .C2(new_n927), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT111), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n913), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n908), .A2(new_n912), .A3(KEYINPUT111), .A4(KEYINPUT38), .ZN(new_n936));
  INV_X1    g0736(.A(new_n662), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n901), .B1(new_n937), .B2(new_n665), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n897), .A2(new_n659), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT37), .B1(new_n939), .B2(new_n901), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n910), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT110), .B(KEYINPUT38), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n935), .A2(new_n936), .A3(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n931), .A2(new_n932), .B1(new_n933), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n923), .A2(new_n927), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n457), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n931), .A2(new_n932), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n933), .A2(new_n945), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(G330), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n752), .B1(new_n923), .B2(new_n927), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n457), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n948), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n344), .A2(new_n707), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT39), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n935), .A2(new_n944), .A3(new_n961), .A4(new_n936), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n914), .A2(new_n930), .ZN(new_n964));
  INV_X1    g0764(.A(new_n870), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n712), .B(new_n965), .C1(new_n693), .C2(new_n697), .ZN(new_n966));
  INV_X1    g0766(.A(new_n871), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n916), .A2(new_n917), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n964), .A2(new_n971), .B1(new_n662), .B2(new_n889), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n963), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n669), .B1(new_n769), .B2(new_n458), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n883), .B1(new_n957), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n957), .B2(new_n975), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n219), .A2(new_n543), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n560), .B2(KEYINPUT35), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n978), .B1(new_n980), .B2(KEYINPUT107), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(KEYINPUT107), .B2(new_n980), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT36), .Z(new_n983));
  INV_X1    g0783(.A(G58), .ZN(new_n984));
  OAI21_X1  g0784(.A(G77), .B1(new_n984), .B2(new_n332), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n217), .A2(new_n985), .B1(new_n332), .B2(new_n201), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(G1), .A3(new_n330), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n977), .A2(new_n983), .A3(new_n987), .ZN(G367));
  AOI22_X1  g0788(.A1(G58), .A2(new_n796), .B1(new_n787), .B2(G137), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n290), .C1(new_n363), .C2(new_n783), .ZN(new_n990));
  INV_X1    g0790(.A(new_n800), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n991), .A2(new_n353), .B1(new_n351), .B2(new_n798), .ZN(new_n992));
  INV_X1    g0792(.A(G143), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n803), .A2(new_n993), .B1(new_n791), .B2(new_n818), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n807), .A2(new_n332), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n990), .A2(new_n992), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n861), .A2(G311), .B1(new_n787), .B2(G317), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n316), .B2(new_n783), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n796), .A2(KEYINPUT46), .A3(G116), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n795), .B2(new_n543), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(new_n294), .C2(new_n807), .ZN(new_n1002));
  INV_X1    g0802(.A(G283), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n802), .B1(new_n798), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(G294), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n991), .A2(new_n522), .B1(new_n791), .B2(new_n1005), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n998), .A2(new_n1002), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n996), .A2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT47), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(KEYINPUT47), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(new_n779), .A3(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n829), .B1(new_n223), .B2(new_n255), .C1(new_n236), .C2(new_n834), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT115), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n776), .A3(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT116), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n649), .B1(new_n650), .B2(new_n627), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n707), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n683), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n677), .B2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1015), .B1(new_n840), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n774), .B(KEYINPUT114), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n603), .B1(new_n599), .B2(new_n712), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n695), .A2(new_n690), .A3(new_n707), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(KEYINPUT113), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n715), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(KEYINPUT113), .C2(new_n1025), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT113), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(KEYINPUT44), .C1(new_n715), .C2(new_n1024), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT45), .B1(new_n715), .B2(new_n1024), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1028), .B(new_n1030), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n725), .A2(new_n727), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n727), .B(new_n710), .Z(new_n1039));
  XNOR2_X1  g0839(.A(new_n725), .B(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n771), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n730), .B(KEYINPUT41), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1021), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n727), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n710), .ZN(new_n1045));
  OR3_X1    g0845(.A1(new_n1045), .A2(KEYINPUT42), .A3(new_n1022), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n519), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n712), .B1(new_n1047), .B2(new_n589), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT42), .B1(new_n1045), .B2(new_n1022), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1035), .A2(new_n1024), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1020), .B1(new_n1043), .B2(new_n1060), .ZN(G387));
  NOR2_X1   g0861(.A1(new_n770), .A2(new_n1040), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n770), .A2(new_n1040), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n730), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n802), .B1(new_n786), .B2(new_n804), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n808), .A2(G283), .B1(new_n796), .B2(G294), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT117), .B(G322), .Z(new_n1068));
  AOI22_X1  g0868(.A1(new_n861), .A2(new_n1068), .B1(new_n792), .B2(G311), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n799), .A2(G303), .B1(new_n800), .B2(G317), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1067), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT49), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1066), .B(new_n1075), .C1(G116), .C2(new_n784), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n248), .A2(new_n792), .B1(new_n787), .B2(G150), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n290), .C1(new_n316), .C2(new_n783), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n795), .A2(new_n363), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G159), .B2(new_n861), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n336), .B2(new_n991), .C1(new_n332), .C2(new_n798), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1078), .B(new_n1081), .C1(new_n254), .C2(new_n808), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n779), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n834), .B1(new_n232), .B2(G45), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n731), .B2(new_n830), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT50), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n248), .B2(new_n336), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n247), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n506), .B1(new_n332), .B2(new_n363), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n731), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1085), .A2(new_n1090), .B1(G107), .B2(new_n223), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n775), .B1(new_n1091), .B2(new_n829), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1083), .B(new_n1092), .C1(new_n1044), .C2(new_n840), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1021), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1065), .B(new_n1093), .C1(new_n1040), .C2(new_n1094), .ZN(G393));
  INV_X1    g0895(.A(new_n1038), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n773), .B1(new_n1096), .B2(new_n1062), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1063), .A2(new_n1038), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1021), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n829), .B1(new_n316), .B2(new_n223), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n834), .A2(new_n243), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n776), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n861), .A2(G317), .B1(new_n800), .B2(G311), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n799), .A2(G294), .B1(new_n787), .B2(new_n1068), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G303), .A2(new_n792), .B1(new_n796), .B2(G283), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n290), .B(new_n814), .C1(G116), .C2(new_n808), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n861), .A2(G150), .B1(new_n800), .B2(G159), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT51), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n795), .A2(new_n332), .B1(new_n786), .B2(new_n993), .ZN(new_n1112));
  OR4_X1    g0912(.A1(new_n802), .A2(new_n1111), .A3(new_n860), .A4(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n351), .A2(new_n791), .B1(new_n798), .B2(new_n247), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT119), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1114), .A2(new_n1115), .B1(G77), .B2(new_n808), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1115), .B2(new_n1114), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT120), .Z(new_n1118));
  OAI21_X1  g0918(.A(new_n1109), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1103), .B1(new_n1119), .B2(new_n779), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1024), .B2(new_n840), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1099), .A2(new_n1100), .A3(new_n1121), .ZN(G390));
  NAND2_X1  g0922(.A1(new_n971), .A2(new_n959), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n960), .A2(new_n1123), .A3(new_n962), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n967), .B1(new_n765), .B2(new_n870), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n970), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n945), .A3(new_n959), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n918), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n953), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n760), .A2(new_n1129), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1132), .A2(KEYINPUT121), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n954), .B(new_n669), .C1(new_n769), .C2(new_n458), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1130), .B1(new_n876), .B2(new_n970), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n968), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1125), .B1(new_n760), .B2(new_n1129), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n872), .B1(new_n953), .B2(KEYINPUT122), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT122), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1141), .B(new_n752), .C1(new_n923), .C2(new_n927), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n969), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1136), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1130), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT121), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1135), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1124), .A2(new_n1134), .A3(new_n1127), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1151));
  AOI211_X1 g0951(.A(KEYINPUT121), .B(new_n1130), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1137), .A2(new_n968), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1151), .A2(new_n1152), .B1(new_n1153), .B2(new_n1136), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1149), .A2(new_n730), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n960), .A2(new_n826), .A3(new_n962), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n776), .B1(new_n846), .B2(new_n248), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n795), .A2(new_n353), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT53), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n784), .A2(new_n201), .B1(new_n800), .B2(G132), .ZN(new_n1161));
  INV_X1    g0961(.A(G125), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1161), .C1(new_n1162), .C2(new_n786), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT54), .B(G143), .Z(new_n1164));
  AOI22_X1  g0964(.A1(new_n799), .A2(new_n1164), .B1(new_n792), .B2(G137), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n802), .B1(new_n861), .B2(G128), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(new_n818), .C2(new_n807), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n799), .A2(G97), .B1(new_n800), .B2(G116), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n294), .B2(new_n791), .C1(new_n1005), .C2(new_n786), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n861), .A2(G283), .B1(new_n784), .B2(G68), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n808), .A2(G77), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1170), .A2(new_n802), .A3(new_n811), .A4(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1163), .A2(new_n1167), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1158), .B1(new_n1173), .B2(new_n779), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1156), .A2(new_n1021), .B1(new_n1157), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1155), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1136), .B1(new_n1156), .B2(new_n1145), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n358), .A2(new_n889), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n377), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n377), .A2(new_n1179), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n951), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n946), .A2(G330), .A3(new_n1186), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1188), .A2(new_n973), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n973), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1177), .B1(new_n1178), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1136), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1194), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1194), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n973), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n951), .A2(new_n1187), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1186), .B1(new_n946), .B2(G330), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1188), .A2(new_n1189), .A3(new_n973), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1199), .A2(KEYINPUT57), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1193), .A2(new_n1206), .A3(new_n730), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1187), .A2(new_n826), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n826), .A2(new_n779), .A3(new_n201), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n800), .A2(G128), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n854), .B2(new_n791), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G137), .A2(new_n799), .B1(new_n796), .B2(new_n1164), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1162), .B2(new_n803), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(G150), .C2(new_n808), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n784), .A2(G159), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n802), .A2(new_n502), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n336), .C1(G33), .C2(G41), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n254), .A2(new_n799), .B1(new_n784), .B2(G58), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n294), .B2(new_n991), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n791), .A2(new_n316), .B1(new_n786), .B2(new_n1003), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1224), .A2(new_n1079), .A3(new_n1221), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n995), .B1(G116), .B2(new_n861), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT123), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT58), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1229), .A2(KEYINPUT58), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1220), .A2(new_n1222), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n775), .B(new_n1209), .C1(new_n1232), .C2(new_n779), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1208), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1205), .B2(new_n1021), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1207), .A2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1153), .A2(new_n1136), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1198), .A2(new_n1042), .A3(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT124), .Z(new_n1239));
  OAI21_X1  g1039(.A(new_n776), .B1(new_n846), .B2(G68), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G97), .A2(new_n796), .B1(new_n800), .B2(G283), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n543), .B2(new_n791), .C1(new_n522), .C2(new_n786), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G294), .A2(new_n861), .B1(new_n799), .B2(G107), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n290), .B1(new_n784), .B2(G77), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n255), .C2(new_n807), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n792), .A2(new_n1164), .B1(new_n796), .B2(G159), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n799), .A2(G150), .B1(new_n787), .B2(G128), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n861), .A2(G132), .B1(new_n800), .B2(G137), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n802), .B1(new_n784), .B2(G58), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n336), .C2(new_n807), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1242), .A2(new_n1245), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1240), .B1(new_n1252), .B2(new_n779), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n970), .B2(new_n827), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1153), .B2(new_n1094), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1239), .A2(new_n1256), .ZN(G381));
  NOR2_X1   g1057(.A1(G375), .A2(G378), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1100), .A2(new_n1121), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n1020), .C1(new_n1043), .C2(new_n1060), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1261), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1256), .A3(new_n1239), .A4(new_n1262), .ZN(G407));
  NAND2_X1  g1063(.A1(new_n1258), .A2(new_n706), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(G213), .A3(new_n1264), .ZN(G409));
  XNOR2_X1  g1065(.A(G393), .B(new_n842), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G390), .A2(G387), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1261), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1268), .B1(new_n1261), .B2(new_n1269), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1267), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1261), .A2(new_n1269), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT126), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1261), .A2(new_n1269), .A3(new_n1268), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1266), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n706), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1235), .A2(new_n1155), .A3(new_n1175), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1149), .A2(new_n1194), .B1(new_n1204), .B2(new_n1203), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1042), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1280), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1235), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n773), .B1(new_n1282), .B2(KEYINPUT57), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1193), .ZN(new_n1287));
  INV_X1    g1087(.A(G378), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1284), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1237), .B1(new_n1145), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n1136), .ZN(new_n1293));
  AND4_X1   g1093(.A1(new_n1290), .A2(new_n1292), .A3(new_n730), .A4(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT60), .B1(new_n1153), .B2(new_n1136), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n773), .B1(new_n1295), .B2(new_n1237), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1290), .B1(new_n1296), .B2(new_n1293), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1256), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n881), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1292), .A2(new_n730), .A3(new_n1293), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT125), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1296), .A2(new_n1290), .A3(new_n1293), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(G384), .A3(new_n1256), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1278), .B1(new_n1289), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G384), .B1(new_n1303), .B2(new_n1256), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n881), .B(new_n1255), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1235), .A2(new_n1155), .A3(new_n1175), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1042), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1178), .A2(new_n1311), .A3(new_n1192), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1279), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(G375), .B2(G378), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1309), .A2(new_n1314), .A3(KEYINPUT62), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1306), .A2(KEYINPUT127), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1317), .B(new_n1278), .C1(new_n1289), .C2(new_n1305), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1280), .A2(G2897), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1321), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1299), .A2(new_n1304), .A3(new_n1320), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n1289), .A3(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1318), .A2(new_n1319), .A3(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1277), .B1(new_n1316), .B2(new_n1325), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1289), .A2(new_n1305), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1277), .B1(KEYINPUT63), .B2(new_n1327), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1327), .A2(KEYINPUT63), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1319), .A4(new_n1324), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1326), .A2(new_n1330), .ZN(G405));
  NOR2_X1   g1131(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1332));
  OR3_X1    g1132(.A1(new_n1309), .A2(new_n1332), .A3(new_n1258), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1277), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1309), .B1(new_n1332), .B2(new_n1258), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1334), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(G402));
endmodule


