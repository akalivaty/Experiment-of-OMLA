

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U550 ( .A1(n521), .A2(G2105), .ZN(n870) );
  NAND2_X1 U551 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XNOR2_X1 U552 ( .A(n536), .B(KEYINPUT89), .ZN(G164) );
  BUF_X1 U553 ( .A(n757), .Z(n540) );
  AND2_X2 U554 ( .A1(n766), .A2(n679), .ZN(n705) );
  NOR2_X2 U555 ( .A1(n529), .A2(n528), .ZN(G160) );
  NAND2_X1 U556 ( .A1(n783), .A2(n782), .ZN(n516) );
  OR2_X1 U557 ( .A1(n779), .A2(n778), .ZN(n517) );
  AND2_X1 U558 ( .A1(n705), .A2(G1996), .ZN(n680) );
  XNOR2_X1 U559 ( .A(KEYINPUT26), .B(n680), .ZN(n681) );
  NOR2_X1 U560 ( .A1(n962), .A2(n684), .ZN(n690) );
  AND2_X1 U561 ( .A1(n726), .A2(n725), .ZN(n727) );
  INV_X1 U562 ( .A(n705), .ZN(n728) );
  NAND2_X1 U563 ( .A1(G8), .A2(n728), .ZN(n781) );
  NOR2_X1 U564 ( .A1(G651), .A2(n646), .ZN(n642) );
  OR2_X1 U565 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X2 U566 ( .A(G2104), .B(KEYINPUT65), .ZN(n521) );
  NOR2_X4 U567 ( .A1(G2105), .A2(n521), .ZN(n867) );
  NAND2_X1 U568 ( .A1(n867), .A2(G101), .ZN(n520) );
  XNOR2_X1 U569 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n518) );
  XNOR2_X1 U570 ( .A(n518), .B(KEYINPUT66), .ZN(n519) );
  XNOR2_X1 U571 ( .A(n520), .B(n519), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n870), .A2(G125), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n524), .Z(n757) );
  NAND2_X1 U576 ( .A1(n757), .A2(G137), .ZN(n527) );
  XOR2_X2 U577 ( .A(KEYINPUT68), .B(n525), .Z(n871) );
  NAND2_X1 U578 ( .A1(G113), .A2(n871), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G126), .A2(n870), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G102), .A2(n867), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U583 ( .A1(n757), .A2(G138), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n871), .A2(G114), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n870), .A2(G123), .ZN(n537) );
  XNOR2_X1 U587 ( .A(n537), .B(KEYINPUT18), .ZN(n539) );
  NAND2_X1 U588 ( .A1(G99), .A2(n867), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n544) );
  NAND2_X1 U590 ( .A1(n540), .A2(G135), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G111), .A2(n871), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U593 ( .A1(n544), .A2(n543), .ZN(n923) );
  XNOR2_X1 U594 ( .A(n923), .B(G2096), .ZN(n545) );
  XNOR2_X1 U595 ( .A(n545), .B(KEYINPUT81), .ZN(n546) );
  OR2_X1 U596 ( .A1(G2100), .A2(n546), .ZN(G156) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  INV_X1 U599 ( .A(G651), .ZN(n550) );
  NOR2_X1 U600 ( .A1(n646), .A2(n550), .ZN(n636) );
  NAND2_X1 U601 ( .A1(G75), .A2(n636), .ZN(n549) );
  NOR2_X1 U602 ( .A1(G543), .A2(G651), .ZN(n547) );
  XNOR2_X1 U603 ( .A(n547), .B(KEYINPUT64), .ZN(n633) );
  NAND2_X1 U604 ( .A1(G88), .A2(n633), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G50), .A2(n642), .ZN(n554) );
  NOR2_X1 U607 ( .A1(G543), .A2(n550), .ZN(n552) );
  XNOR2_X1 U608 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n552), .B(n551), .ZN(n649) );
  NAND2_X1 U610 ( .A1(G62), .A2(n649), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U612 ( .A1(n556), .A2(n555), .ZN(G166) );
  NAND2_X1 U613 ( .A1(G52), .A2(n642), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G64), .A2(n649), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G77), .A2(n636), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G90), .A2(n633), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U620 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U621 ( .A1(G94), .A2(G452), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n564), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n819) );
  NAND2_X1 U626 ( .A1(n819), .A2(G567), .ZN(n566) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U628 ( .A1(G81), .A2(n633), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G68), .A2(n636), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(n570), .ZN(n577) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n572) );
  NAND2_X1 U634 ( .A1(G56), .A2(n649), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n572), .B(n571), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G43), .A2(n642), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT77), .B(n573), .ZN(n574) );
  NOR2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n962) );
  INV_X1 U640 ( .A(G860), .ZN(n610) );
  OR2_X1 U641 ( .A1(n962), .A2(n610), .ZN(G153) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U644 ( .A1(G79), .A2(n636), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G92), .A2(n633), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G54), .A2(n642), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G66), .A2(n649), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT15), .B(n584), .Z(n892) );
  INV_X1 U652 ( .A(n892), .ZN(n972) );
  INV_X1 U653 ( .A(G868), .ZN(n662) );
  NAND2_X1 U654 ( .A1(n972), .A2(n662), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(G284) );
  XNOR2_X1 U656 ( .A(KEYINPUT7), .B(KEYINPUT80), .ZN(n599) );
  NAND2_X1 U657 ( .A1(G89), .A2(n633), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT4), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G76), .A2(n636), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT5), .ZN(n597) );
  XNOR2_X1 U662 ( .A(KEYINPUT6), .B(KEYINPUT79), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n642), .A2(G51), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT78), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G63), .A2(n649), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n595), .B(n594), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n599), .B(n598), .ZN(G168) );
  XOR2_X1 U670 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U671 ( .A1(n636), .A2(G78), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT72), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G91), .A2(n633), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U675 ( .A(KEYINPUT73), .B(n603), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n642), .A2(G53), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G65), .A2(n649), .ZN(n604) );
  AND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(G299) );
  NAND2_X1 U680 ( .A1(G868), .A2(G286), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G299), .A2(n662), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U683 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n611), .A2(n892), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n962), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G868), .A2(n892), .ZN(n613) );
  NOR2_X1 U688 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G80), .A2(n636), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G67), .A2(n649), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G93), .A2(n633), .ZN(n618) );
  XNOR2_X1 U694 ( .A(KEYINPUT83), .B(n618), .ZN(n619) );
  NOR2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n642), .A2(G55), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n663) );
  NAND2_X1 U698 ( .A1(G559), .A2(n892), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT82), .ZN(n659) );
  XNOR2_X1 U700 ( .A(n659), .B(n962), .ZN(n624) );
  NOR2_X1 U701 ( .A1(G860), .A2(n624), .ZN(n625) );
  XOR2_X1 U702 ( .A(n663), .B(n625), .Z(G145) );
  NAND2_X1 U703 ( .A1(G72), .A2(n636), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G85), .A2(n633), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G60), .A2(n649), .ZN(n628) );
  XOR2_X1 U707 ( .A(KEYINPUT70), .B(n628), .Z(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n642), .A2(G47), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U711 ( .A1(n649), .A2(G61), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G86), .A2(n633), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n636), .A2(G73), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n637), .Z(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(G48), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U719 ( .A1(G49), .A2(n642), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT84), .B(n645), .Z(n648) );
  NAND2_X1 U723 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n650) );
  NOR2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n651), .B(KEYINPUT85), .ZN(G288) );
  INV_X1 U727 ( .A(G299), .ZN(n699) );
  XNOR2_X1 U728 ( .A(n699), .B(n962), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U730 ( .A(G290), .B(G166), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n656) );
  XOR2_X1 U732 ( .A(G305), .B(G288), .Z(n654) );
  XNOR2_X1 U733 ( .A(n663), .B(n654), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n658), .B(n657), .ZN(n889) );
  XNOR2_X1 U736 ( .A(n889), .B(n659), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n660), .A2(G868), .ZN(n661) );
  XOR2_X1 U738 ( .A(KEYINPUT87), .B(n661), .Z(n665) );
  NAND2_X1 U739 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n666) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U745 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XOR2_X1 U746 ( .A(KEYINPUT74), .B(G57), .Z(G237) );
  XNOR2_X1 U747 ( .A(KEYINPUT88), .B(G44), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U749 ( .A(KEYINPUT75), .B(G132), .ZN(G219) );
  NAND2_X1 U750 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U751 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G69), .A2(n672), .ZN(n824) );
  NAND2_X1 U753 ( .A1(n824), .A2(G567), .ZN(n677) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U756 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G96), .A2(n675), .ZN(n823) );
  NAND2_X1 U758 ( .A1(n823), .A2(G2106), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n677), .A2(n676), .ZN(n826) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U761 ( .A1(n826), .A2(n678), .ZN(n822) );
  NAND2_X1 U762 ( .A1(n822), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n766) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n765) );
  INV_X1 U766 ( .A(n765), .ZN(n679) );
  NAND2_X1 U767 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U768 ( .A(n681), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n728), .A2(G1341), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n892), .A2(n690), .ZN(n689) );
  NAND2_X1 U772 ( .A1(n728), .A2(G1348), .ZN(n685) );
  XNOR2_X1 U773 ( .A(n685), .B(KEYINPUT96), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n705), .A2(G2067), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U776 ( .A1(n689), .A2(n688), .ZN(n692) );
  OR2_X1 U777 ( .A1(n690), .A2(n892), .ZN(n691) );
  NAND2_X1 U778 ( .A1(n692), .A2(n691), .ZN(n697) );
  NAND2_X1 U779 ( .A1(n705), .A2(G2072), .ZN(n693) );
  XNOR2_X1 U780 ( .A(n693), .B(KEYINPUT27), .ZN(n695) );
  INV_X1 U781 ( .A(G1956), .ZN(n990) );
  NOR2_X1 U782 ( .A1(n990), .A2(n705), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n699), .A2(n698), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n703) );
  NOR2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U787 ( .A(KEYINPUT28), .B(KEYINPUT95), .ZN(n700) );
  XNOR2_X1 U788 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U790 ( .A(n704), .B(KEYINPUT29), .ZN(n710) );
  NAND2_X1 U791 ( .A1(n728), .A2(G1961), .ZN(n707) );
  XOR2_X1 U792 ( .A(KEYINPUT25), .B(G2078), .Z(n941) );
  NAND2_X1 U793 ( .A1(n705), .A2(n941), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U795 ( .A(n708), .B(KEYINPUT94), .Z(n715) );
  AND2_X1 U796 ( .A1(G171), .A2(n715), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n720) );
  NOR2_X1 U798 ( .A1(G1966), .A2(n781), .ZN(n724) );
  NOR2_X1 U799 ( .A1(G2084), .A2(n728), .ZN(n722) );
  INV_X1 U800 ( .A(n722), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n711), .A2(G8), .ZN(n712) );
  OR2_X1 U802 ( .A1(n724), .A2(n712), .ZN(n713) );
  XNOR2_X1 U803 ( .A(KEYINPUT30), .B(n713), .ZN(n714) );
  NOR2_X1 U804 ( .A1(G168), .A2(n714), .ZN(n717) );
  NOR2_X1 U805 ( .A1(G171), .A2(n715), .ZN(n716) );
  NOR2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U807 ( .A(n718), .B(KEYINPUT31), .ZN(n719) );
  NOR2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U809 ( .A(n721), .B(KEYINPUT97), .ZN(n732) );
  XNOR2_X1 U810 ( .A(n732), .B(KEYINPUT98), .ZN(n726) );
  AND2_X1 U811 ( .A1(n722), .A2(G8), .ZN(n723) );
  NOR2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U813 ( .A(n727), .B(KEYINPUT99), .ZN(n738) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n781), .ZN(n730) );
  NOR2_X1 U815 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U817 ( .A1(G303), .A2(n731), .ZN(n734) );
  NAND2_X1 U818 ( .A1(n732), .A2(G286), .ZN(n733) );
  NAND2_X1 U819 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n735), .A2(G8), .ZN(n736) );
  XNOR2_X1 U821 ( .A(KEYINPUT32), .B(n736), .ZN(n737) );
  NAND2_X1 U822 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U823 ( .A(n739), .B(KEYINPUT100), .ZN(n773) );
  NOR2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NOR2_X1 U825 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U826 ( .A1(n744), .A2(n740), .ZN(n981) );
  NAND2_X1 U827 ( .A1(n773), .A2(n981), .ZN(n741) );
  NAND2_X1 U828 ( .A1(n980), .A2(n741), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n781), .A2(n742), .ZN(n743) );
  NOR2_X1 U830 ( .A1(KEYINPUT33), .A2(n743), .ZN(n747) );
  NAND2_X1 U831 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n745), .A2(n781), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n771) );
  XOR2_X1 U834 ( .A(G1981), .B(G305), .Z(n967) );
  NAND2_X1 U835 ( .A1(n540), .A2(G141), .ZN(n749) );
  NAND2_X1 U836 ( .A1(G117), .A2(n871), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n867), .A2(G105), .ZN(n750) );
  XOR2_X1 U839 ( .A(KEYINPUT38), .B(n750), .Z(n751) );
  NOR2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n870), .A2(G129), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n881) );
  AND2_X1 U843 ( .A1(n881), .A2(G1996), .ZN(n764) );
  NAND2_X1 U844 ( .A1(n870), .A2(G119), .ZN(n756) );
  NAND2_X1 U845 ( .A1(G107), .A2(n871), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n762) );
  NAND2_X1 U847 ( .A1(G131), .A2(n757), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G95), .A2(n867), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U850 ( .A(KEYINPUT93), .B(n760), .Z(n761) );
  OR2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n878) );
  AND2_X1 U852 ( .A1(n878), .A2(G1991), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n921) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n813) );
  INV_X1 U855 ( .A(n813), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n921), .A2(n767), .ZN(n806) );
  XNOR2_X1 U857 ( .A(G1986), .B(G290), .ZN(n964) );
  NAND2_X1 U858 ( .A1(n964), .A2(n813), .ZN(n768) );
  XOR2_X1 U859 ( .A(KEYINPUT90), .B(n768), .Z(n769) );
  NOR2_X1 U860 ( .A1(n806), .A2(n769), .ZN(n772) );
  AND2_X1 U861 ( .A1(n967), .A2(n772), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n787) );
  INV_X1 U863 ( .A(n772), .ZN(n785) );
  INV_X1 U864 ( .A(n773), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G166), .A2(G8), .ZN(n774) );
  NOR2_X1 U866 ( .A1(G2090), .A2(n774), .ZN(n777) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U868 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  NOR2_X1 U869 ( .A1(n781), .A2(n776), .ZN(n780) );
  OR2_X1 U870 ( .A1(n777), .A2(n780), .ZN(n778) );
  INV_X1 U871 ( .A(n780), .ZN(n783) );
  INV_X1 U872 ( .A(n781), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n517), .A2(n516), .ZN(n784) );
  OR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n800) );
  XNOR2_X1 U876 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  NAND2_X1 U877 ( .A1(G116), .A2(n871), .ZN(n788) );
  XOR2_X1 U878 ( .A(KEYINPUT91), .B(n788), .Z(n790) );
  NAND2_X1 U879 ( .A1(n870), .A2(G128), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U881 ( .A(KEYINPUT35), .B(n791), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n867), .A2(G104), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n540), .A2(G140), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U885 ( .A(KEYINPUT34), .B(n794), .Z(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U887 ( .A(KEYINPUT36), .B(n797), .Z(n885) );
  NOR2_X1 U888 ( .A1(n801), .A2(n885), .ZN(n928) );
  NAND2_X1 U889 ( .A1(n928), .A2(n813), .ZN(n798) );
  XOR2_X1 U890 ( .A(KEYINPUT92), .B(n798), .Z(n810) );
  INV_X1 U891 ( .A(n810), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n817) );
  AND2_X1 U893 ( .A1(n801), .A2(n885), .ZN(n935) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n881), .ZN(n802) );
  XOR2_X1 U895 ( .A(KEYINPUT101), .B(n802), .Z(n918) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U897 ( .A1(n878), .A2(G1991), .ZN(n803) );
  XNOR2_X1 U898 ( .A(n803), .B(KEYINPUT102), .ZN(n922) );
  NOR2_X1 U899 ( .A1(n804), .A2(n922), .ZN(n805) );
  NOR2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n918), .A2(n807), .ZN(n808) );
  XOR2_X1 U902 ( .A(KEYINPUT39), .B(n808), .Z(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n935), .A2(n811), .ZN(n812) );
  XNOR2_X1 U905 ( .A(KEYINPUT103), .B(n812), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U907 ( .A(n815), .B(KEYINPUT104), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U909 ( .A(KEYINPUT40), .B(n818), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(G188) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G108), .ZN(G238) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U922 ( .A(G261), .ZN(G325) );
  INV_X1 U923 ( .A(n826), .ZN(G319) );
  XOR2_X1 U924 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n828) );
  XNOR2_X1 U925 ( .A(KEYINPUT42), .B(G2678), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U927 ( .A(KEYINPUT106), .B(G2072), .Z(n830) );
  XNOR2_X1 U928 ( .A(G2067), .B(G2090), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U930 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U931 ( .A(G2096), .B(G2100), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n836) );
  XOR2_X1 U933 ( .A(G2084), .B(G2078), .Z(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1981), .B(G1966), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1991), .B(G1996), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n848) );
  XOR2_X1 U938 ( .A(KEYINPUT41), .B(KEYINPUT109), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1986), .B(KEYINPUT108), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(G1976), .B(G1971), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1961), .B(G1956), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U945 ( .A(G2474), .B(KEYINPUT110), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U948 ( .A1(n870), .A2(G124), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U950 ( .A1(G100), .A2(n867), .ZN(n850) );
  NAND2_X1 U951 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n540), .A2(G136), .ZN(n853) );
  NAND2_X1 U953 ( .A1(G112), .A2(n871), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U955 ( .A1(n855), .A2(n854), .ZN(G162) );
  XOR2_X1 U956 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n857) );
  XNOR2_X1 U957 ( .A(KEYINPUT112), .B(KEYINPUT111), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n866) );
  NAND2_X1 U959 ( .A1(n870), .A2(G130), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G118), .A2(n871), .ZN(n858) );
  NAND2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G142), .A2(n540), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G106), .A2(n867), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U965 ( .A(n862), .B(KEYINPUT45), .Z(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U967 ( .A(n866), .B(n865), .Z(n877) );
  NAND2_X1 U968 ( .A1(G139), .A2(n540), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G103), .A2(n867), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U971 ( .A1(n870), .A2(G127), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G115), .A2(n871), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n912) );
  XOR2_X1 U976 ( .A(n877), .B(n912), .Z(n880) );
  XOR2_X1 U977 ( .A(n878), .B(n923), .Z(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n887) );
  XNOR2_X1 U979 ( .A(G162), .B(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U982 ( .A(n885), .B(n884), .Z(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U984 ( .A1(G37), .A2(n888), .ZN(G395) );
  XOR2_X1 U985 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n891) );
  XNOR2_X1 U986 ( .A(G171), .B(n889), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n894) );
  XOR2_X1 U988 ( .A(G286), .B(n892), .Z(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2451), .B(G2430), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2438), .B(G2443), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n903) );
  XOR2_X1 U994 ( .A(G2435), .B(G2454), .Z(n899) );
  XNOR2_X1 U995 ( .A(G1341), .B(G1348), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U997 ( .A(G2446), .B(G2427), .Z(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(n903), .B(n902), .Z(n904) );
  NAND2_X1 U1000 ( .A1(G14), .A2(n904), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n905) );
  XOR2_X1 U1003 ( .A(KEYINPUT49), .B(n905), .Z(n906) );
  XNOR2_X1 U1004 ( .A(n906), .B(KEYINPUT115), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(n911), .ZN(G401) );
  XOR2_X1 U1010 ( .A(G2072), .B(n912), .Z(n914) );
  XOR2_X1 U1011 ( .A(G164), .B(G2078), .Z(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT50), .B(n915), .ZN(n933) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT118), .B(n916), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1017 ( .A(KEYINPUT51), .B(n919), .Z(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n931) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(KEYINPUT116), .B(n924), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(KEYINPUT117), .B(n929), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n936), .ZN(n937) );
  INV_X1 U1029 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n957), .ZN(n938) );
  NAND2_X1 U1031 ( .A1(n938), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1032 ( .A(G2090), .B(G35), .ZN(n952) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(G1996), .B(G32), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(n941), .B(G27), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT119), .B(n946), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n947), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G25), .B(G1991), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT53), .B(n950), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1046 ( .A(G2084), .B(G34), .Z(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(n953), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(n957), .B(n956), .ZN(n959) );
  INV_X1 U1050 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n960), .ZN(n1018) );
  XNOR2_X1 U1053 ( .A(G16), .B(KEYINPUT56), .ZN(n988) );
  XOR2_X1 U1054 ( .A(G1341), .B(KEYINPUT124), .Z(n961) );
  XNOR2_X1 U1055 ( .A(n962), .B(n961), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G1956), .B(G299), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n979) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G168), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n969), .B(KEYINPUT121), .ZN(n970) );
  XOR2_X1 U1063 ( .A(n971), .B(n970), .Z(n977) );
  XNOR2_X1 U1064 ( .A(G301), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n972), .B(G1348), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(KEYINPUT122), .B(n975), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n986) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n983) );
  AND2_X1 U1071 ( .A1(G303), .A2(G1971), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1073 ( .A(KEYINPUT123), .B(n984), .Z(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n1016) );
  INV_X1 U1076 ( .A(G16), .ZN(n1014) );
  XNOR2_X1 U1077 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n1012) );
  XNOR2_X1 U1078 ( .A(KEYINPUT125), .B(G1961), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n989), .B(G5), .ZN(n1010) );
  XOR2_X1 U1080 ( .A(G1966), .B(G21), .Z(n1000) );
  XNOR2_X1 U1081 ( .A(G20), .B(n990), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1086 ( .A(KEYINPUT59), .B(G1348), .Z(n995) );
  XNOR2_X1 U1087 ( .A(G4), .B(n995), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(KEYINPUT60), .B(n998), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(G1986), .B(KEYINPUT126), .Z(n1003) );
  XNOR2_X1 U1095 ( .A(G24), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

