

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U547 ( .A(n674), .B(KEYINPUT32), .ZN(n699) );
  XOR2_X1 U548 ( .A(n666), .B(KEYINPUT96), .Z(n643) );
  XOR2_X1 U549 ( .A(n654), .B(KEYINPUT29), .Z(n512) );
  NOR2_X1 U550 ( .A1(n706), .A2(n693), .ZN(n513) );
  AND2_X1 U551 ( .A1(n692), .A2(n513), .ZN(n696) );
  NOR2_X1 U552 ( .A1(G164), .A2(G1384), .ZN(n601) );
  NOR2_X2 U553 ( .A1(G2105), .A2(n516), .ZN(n863) );
  NOR2_X1 U554 ( .A1(n572), .A2(G651), .ZN(n783) );
  AND2_X1 U555 ( .A1(n522), .A2(n521), .ZN(G164) );
  NOR2_X1 U556 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XOR2_X2 U557 ( .A(KEYINPUT17), .B(n514), .Z(n862) );
  NAND2_X1 U558 ( .A1(G138), .A2(n862), .ZN(n515) );
  XNOR2_X1 U559 ( .A(n515), .B(KEYINPUT90), .ZN(n522) );
  AND2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n867) );
  AND2_X1 U561 ( .A1(n867), .A2(G114), .ZN(n520) );
  XOR2_X1 U562 ( .A(KEYINPUT66), .B(G2104), .Z(n516) );
  NAND2_X1 U563 ( .A1(G102), .A2(n863), .ZN(n518) );
  AND2_X1 U564 ( .A1(G2105), .A2(n516), .ZN(n870) );
  NAND2_X1 U565 ( .A1(G126), .A2(n870), .ZN(n517) );
  NAND2_X1 U566 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n862), .A2(G137), .ZN(n525) );
  NAND2_X1 U569 ( .A1(G101), .A2(n863), .ZN(n523) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  NAND2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U572 ( .A1(G113), .A2(n867), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G125), .A2(n870), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U575 ( .A1(n529), .A2(n528), .ZN(G160) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n530) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n530), .Z(n778) );
  NAND2_X1 U578 ( .A1(G85), .A2(n778), .ZN(n532) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n572) );
  INV_X1 U580 ( .A(G651), .ZN(n534) );
  NOR2_X1 U581 ( .A1(n572), .A2(n534), .ZN(n782) );
  NAND2_X1 U582 ( .A1(G72), .A2(n782), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U584 ( .A(KEYINPUT67), .B(n533), .ZN(n539) );
  NOR2_X1 U585 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n535), .Z(n779) );
  NAND2_X1 U587 ( .A1(G60), .A2(n779), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G47), .A2(n783), .ZN(n536) );
  AND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n539), .A2(n538), .ZN(G290) );
  NAND2_X1 U591 ( .A1(n778), .A2(G90), .ZN(n540) );
  XOR2_X1 U592 ( .A(KEYINPUT69), .B(n540), .Z(n542) );
  NAND2_X1 U593 ( .A1(n782), .A2(G77), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U595 ( .A(KEYINPUT9), .B(n543), .ZN(n548) );
  NAND2_X1 U596 ( .A1(G64), .A2(n779), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G52), .A2(n783), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U599 ( .A(KEYINPUT68), .B(n546), .Z(n547) );
  NAND2_X1 U600 ( .A1(n548), .A2(n547), .ZN(G301) );
  INV_X1 U601 ( .A(G301), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G63), .A2(n779), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G51), .A2(n783), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U605 ( .A(KEYINPUT6), .B(n551), .ZN(n559) );
  XOR2_X1 U606 ( .A(KEYINPUT4), .B(KEYINPUT77), .Z(n553) );
  NAND2_X1 U607 ( .A1(G89), .A2(n778), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U609 ( .A(KEYINPUT76), .B(n554), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n782), .A2(G76), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U612 ( .A(n557), .B(KEYINPUT5), .Z(n558) );
  NOR2_X1 U613 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(n560), .Z(n561) );
  XNOR2_X1 U615 ( .A(KEYINPUT78), .B(n561), .ZN(G168) );
  XOR2_X1 U616 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U617 ( .A1(G75), .A2(n782), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G50), .A2(n783), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U620 ( .A1(G88), .A2(n778), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G62), .A2(n779), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U624 ( .A(n568), .B(KEYINPUT83), .ZN(G303) );
  INV_X1 U625 ( .A(G303), .ZN(G166) );
  NAND2_X1 U626 ( .A1(G49), .A2(n783), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U629 ( .A1(n779), .A2(n571), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n572), .A2(G87), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(G288) );
  NAND2_X1 U632 ( .A1(G86), .A2(n778), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G61), .A2(n779), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n782), .A2(G73), .ZN(n577) );
  XOR2_X1 U636 ( .A(KEYINPUT2), .B(n577), .Z(n578) );
  NOR2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n783), .A2(G48), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U640 ( .A1(G160), .A2(G40), .ZN(n600) );
  NOR2_X1 U641 ( .A1(n601), .A2(n600), .ZN(n739) );
  NAND2_X1 U642 ( .A1(G107), .A2(n867), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G119), .A2(n870), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n862), .A2(G131), .ZN(n584) );
  XOR2_X1 U646 ( .A(KEYINPUT94), .B(n584), .Z(n585) );
  NOR2_X1 U647 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n863), .A2(G95), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n588), .A2(n587), .ZN(n875) );
  NAND2_X1 U650 ( .A1(G1991), .A2(n875), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT95), .B(n589), .Z(n598) );
  NAND2_X1 U652 ( .A1(G141), .A2(n862), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G117), .A2(n867), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U655 ( .A1(n863), .A2(G105), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT38), .B(n592), .Z(n593) );
  NOR2_X1 U657 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U658 ( .A1(n870), .A2(G129), .ZN(n595) );
  NAND2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n860) );
  NAND2_X1 U660 ( .A1(G1996), .A2(n860), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n911) );
  NAND2_X1 U662 ( .A1(n739), .A2(n911), .ZN(n727) );
  XNOR2_X1 U663 ( .A(G1986), .B(G290), .ZN(n957) );
  NAND2_X1 U664 ( .A1(n739), .A2(n957), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n727), .A2(n599), .ZN(n712) );
  INV_X1 U666 ( .A(n600), .ZN(n602) );
  NAND2_X2 U667 ( .A1(n602), .A2(n601), .ZN(n666) );
  XNOR2_X1 U668 ( .A(G2078), .B(KEYINPUT25), .ZN(n928) );
  NAND2_X1 U669 ( .A1(n643), .A2(n928), .ZN(n604) );
  INV_X1 U670 ( .A(G1961), .ZN(n979) );
  NAND2_X1 U671 ( .A1(n979), .A2(n666), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n656) );
  NAND2_X1 U673 ( .A1(n656), .A2(G171), .ZN(n655) );
  NAND2_X1 U674 ( .A1(G65), .A2(n779), .ZN(n606) );
  NAND2_X1 U675 ( .A1(G53), .A2(n783), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U677 ( .A1(G91), .A2(n778), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G78), .A2(n782), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n901) );
  NAND2_X1 U681 ( .A1(G2072), .A2(n643), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT27), .ZN(n614) );
  INV_X1 U683 ( .A(G1956), .ZN(n612) );
  NOR2_X1 U684 ( .A1(n643), .A2(n612), .ZN(n613) );
  NOR2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n617) );
  NOR2_X1 U686 ( .A1(n901), .A2(n617), .ZN(n616) );
  INV_X1 U687 ( .A(KEYINPUT28), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n653) );
  NAND2_X1 U689 ( .A1(n901), .A2(n617), .ZN(n651) );
  NAND2_X1 U690 ( .A1(G54), .A2(n783), .ZN(n624) );
  NAND2_X1 U691 ( .A1(G79), .A2(n782), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G66), .A2(n779), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n778), .A2(G92), .ZN(n620) );
  XOR2_X1 U695 ( .A(KEYINPUT74), .B(n620), .Z(n621) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(KEYINPUT15), .ZN(n963) );
  NAND2_X1 U699 ( .A1(G56), .A2(n779), .ZN(n626) );
  XOR2_X1 U700 ( .A(KEYINPUT14), .B(n626), .Z(n634) );
  XOR2_X1 U701 ( .A(KEYINPUT12), .B(KEYINPUT72), .Z(n628) );
  NAND2_X1 U702 ( .A1(G81), .A2(n778), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n628), .B(n627), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n782), .A2(G68), .ZN(n629) );
  XNOR2_X1 U705 ( .A(KEYINPUT73), .B(n629), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n632), .B(KEYINPUT13), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n783), .A2(G43), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n961) );
  INV_X1 U711 ( .A(G1996), .ZN(n929) );
  NOR2_X1 U712 ( .A1(n666), .A2(n929), .ZN(n638) );
  XOR2_X1 U713 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n637) );
  XNOR2_X1 U714 ( .A(n638), .B(n637), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n666), .A2(G1341), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n961), .A2(n641), .ZN(n642) );
  OR2_X1 U718 ( .A1(n963), .A2(n642), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n963), .A2(n642), .ZN(n647) );
  NAND2_X1 U720 ( .A1(G2067), .A2(n643), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G1348), .A2(n666), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n512), .ZN(n677) );
  NOR2_X1 U728 ( .A1(G171), .A2(n656), .ZN(n662) );
  NAND2_X1 U729 ( .A1(G8), .A2(n666), .ZN(n706) );
  NOR2_X1 U730 ( .A1(G1966), .A2(n706), .ZN(n679) );
  NOR2_X1 U731 ( .A1(G2084), .A2(n666), .ZN(n675) );
  NOR2_X1 U732 ( .A1(n679), .A2(n675), .ZN(n657) );
  XOR2_X1 U733 ( .A(KEYINPUT97), .B(n657), .Z(n658) );
  NAND2_X1 U734 ( .A1(G8), .A2(n658), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(KEYINPUT30), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n660), .A2(G168), .ZN(n661) );
  NOR2_X1 U737 ( .A1(n662), .A2(n661), .ZN(n664) );
  XOR2_X1 U738 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n663) );
  XNOR2_X1 U739 ( .A(n664), .B(n663), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n665), .A2(G286), .ZN(n672) );
  NOR2_X1 U742 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U743 ( .A(KEYINPUT99), .B(n667), .ZN(n670) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n706), .ZN(n668) );
  NOR2_X1 U745 ( .A1(G166), .A2(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U748 ( .A1(n673), .A2(G8), .ZN(n674) );
  NAND2_X1 U749 ( .A1(G8), .A2(n675), .ZN(n681) );
  AND2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n700) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n953) );
  AND2_X1 U754 ( .A1(n700), .A2(n953), .ZN(n682) );
  NAND2_X1 U755 ( .A1(n699), .A2(n682), .ZN(n689) );
  INV_X1 U756 ( .A(n953), .ZN(n687) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n683) );
  XOR2_X1 U759 ( .A(KEYINPUT100), .B(n683), .Z(n954) );
  INV_X1 U760 ( .A(n954), .ZN(n684) );
  NOR2_X1 U761 ( .A1(n685), .A2(n684), .ZN(n686) );
  OR2_X1 U762 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U763 ( .A1(n689), .A2(n688), .ZN(n692) );
  NOR2_X1 U764 ( .A1(n954), .A2(n706), .ZN(n690) );
  AND2_X1 U765 ( .A1(KEYINPUT33), .A2(n690), .ZN(n691) );
  XNOR2_X1 U766 ( .A(G1981), .B(G305), .ZN(n970) );
  OR2_X1 U767 ( .A1(n691), .A2(n970), .ZN(n693) );
  INV_X1 U768 ( .A(n693), .ZN(n694) );
  AND2_X1 U769 ( .A1(n694), .A2(KEYINPUT33), .ZN(n695) );
  NOR2_X1 U770 ( .A1(n696), .A2(n695), .ZN(n710) );
  NAND2_X1 U771 ( .A1(G8), .A2(G166), .ZN(n697) );
  NOR2_X1 U772 ( .A1(G2090), .A2(n697), .ZN(n698) );
  XNOR2_X1 U773 ( .A(n698), .B(KEYINPUT101), .ZN(n702) );
  NAND2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U776 ( .A1(n703), .A2(n706), .ZN(n708) );
  NOR2_X1 U777 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U778 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  NOR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U781 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n725) );
  NAND2_X1 U783 ( .A1(G140), .A2(n862), .ZN(n714) );
  NAND2_X1 U784 ( .A1(G104), .A2(n863), .ZN(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U786 ( .A(KEYINPUT34), .B(n715), .ZN(n720) );
  NAND2_X1 U787 ( .A1(G116), .A2(n867), .ZN(n717) );
  NAND2_X1 U788 ( .A1(G128), .A2(n870), .ZN(n716) );
  NAND2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U790 ( .A(n718), .B(KEYINPUT35), .Z(n719) );
  NOR2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U792 ( .A(KEYINPUT36), .B(n721), .Z(n722) );
  XOR2_X1 U793 ( .A(KEYINPUT92), .B(n722), .Z(n884) );
  XOR2_X1 U794 ( .A(G2067), .B(KEYINPUT37), .Z(n723) );
  XNOR2_X1 U795 ( .A(KEYINPUT91), .B(n723), .ZN(n736) );
  NOR2_X1 U796 ( .A1(n884), .A2(n736), .ZN(n919) );
  NAND2_X1 U797 ( .A1(n919), .A2(n739), .ZN(n724) );
  XOR2_X1 U798 ( .A(KEYINPUT93), .B(n724), .Z(n734) );
  NAND2_X1 U799 ( .A1(n725), .A2(n734), .ZN(n726) );
  XNOR2_X1 U800 ( .A(n726), .B(KEYINPUT102), .ZN(n742) );
  NOR2_X1 U801 ( .A1(G1996), .A2(n860), .ZN(n903) );
  INV_X1 U802 ( .A(n727), .ZN(n730) );
  NOR2_X1 U803 ( .A1(G1991), .A2(n875), .ZN(n916) );
  NOR2_X1 U804 ( .A1(G1986), .A2(G290), .ZN(n728) );
  NOR2_X1 U805 ( .A1(n916), .A2(n728), .ZN(n729) );
  NOR2_X1 U806 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U807 ( .A(KEYINPUT103), .B(n731), .Z(n732) );
  NOR2_X1 U808 ( .A1(n903), .A2(n732), .ZN(n733) );
  XNOR2_X1 U809 ( .A(KEYINPUT39), .B(n733), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n884), .A2(n736), .ZN(n910) );
  NAND2_X1 U812 ( .A1(n737), .A2(n910), .ZN(n738) );
  XNOR2_X1 U813 ( .A(KEYINPUT104), .B(n738), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U815 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U816 ( .A(n743), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U817 ( .A(G2443), .B(G2446), .Z(n745) );
  XNOR2_X1 U818 ( .A(G2427), .B(G2451), .ZN(n744) );
  XNOR2_X1 U819 ( .A(n745), .B(n744), .ZN(n751) );
  XOR2_X1 U820 ( .A(G2430), .B(G2454), .Z(n747) );
  XNOR2_X1 U821 ( .A(G1341), .B(G1348), .ZN(n746) );
  XNOR2_X1 U822 ( .A(n747), .B(n746), .ZN(n749) );
  XOR2_X1 U823 ( .A(G2435), .B(G2438), .Z(n748) );
  XNOR2_X1 U824 ( .A(n749), .B(n748), .ZN(n750) );
  XOR2_X1 U825 ( .A(n751), .B(n750), .Z(n752) );
  AND2_X1 U826 ( .A1(G14), .A2(n752), .ZN(G401) );
  AND2_X1 U827 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U828 ( .A1(G135), .A2(n862), .ZN(n754) );
  NAND2_X1 U829 ( .A1(G111), .A2(n867), .ZN(n753) );
  NAND2_X1 U830 ( .A1(n754), .A2(n753), .ZN(n757) );
  NAND2_X1 U831 ( .A1(n870), .A2(G123), .ZN(n755) );
  XOR2_X1 U832 ( .A(KEYINPUT18), .B(n755), .Z(n756) );
  NOR2_X1 U833 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U834 ( .A1(n863), .A2(G99), .ZN(n758) );
  NAND2_X1 U835 ( .A1(n759), .A2(n758), .ZN(n917) );
  XNOR2_X1 U836 ( .A(G2096), .B(n917), .ZN(n760) );
  OR2_X1 U837 ( .A1(G2100), .A2(n760), .ZN(G156) );
  INV_X1 U838 ( .A(G132), .ZN(G219) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U841 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U842 ( .A(G223), .B(KEYINPUT71), .ZN(n819) );
  NAND2_X1 U843 ( .A1(n819), .A2(G567), .ZN(n762) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U845 ( .A(G860), .ZN(n769) );
  OR2_X1 U846 ( .A1(n961), .A2(n769), .ZN(G153) );
  NAND2_X1 U847 ( .A1(G868), .A2(G171), .ZN(n764) );
  INV_X1 U848 ( .A(G868), .ZN(n799) );
  NAND2_X1 U849 ( .A1(n963), .A2(n799), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n765), .B(KEYINPUT75), .ZN(G284) );
  NAND2_X1 U852 ( .A1(n901), .A2(n799), .ZN(n766) );
  XNOR2_X1 U853 ( .A(n766), .B(KEYINPUT79), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G286), .A2(n799), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n769), .A2(G559), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n770), .A2(n963), .ZN(n771) );
  XNOR2_X1 U858 ( .A(n771), .B(KEYINPUT16), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT80), .B(n772), .ZN(G148) );
  NOR2_X1 U860 ( .A1(G868), .A2(n961), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G868), .A2(n963), .ZN(n773) );
  NOR2_X1 U862 ( .A1(G559), .A2(n773), .ZN(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(G282) );
  NAND2_X1 U864 ( .A1(G559), .A2(n963), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT81), .B(n776), .Z(n777) );
  XNOR2_X1 U866 ( .A(n961), .B(n777), .ZN(n796) );
  NOR2_X1 U867 ( .A1(G860), .A2(n796), .ZN(n789) );
  NAND2_X1 U868 ( .A1(G93), .A2(n778), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G67), .A2(n779), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G80), .A2(n782), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G55), .A2(n783), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n800) );
  XOR2_X1 U875 ( .A(n800), .B(KEYINPUT82), .Z(n788) );
  XNOR2_X1 U876 ( .A(n789), .B(n788), .ZN(G145) );
  XOR2_X1 U877 ( .A(n800), .B(G288), .Z(n795) );
  XNOR2_X1 U878 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n791) );
  XNOR2_X1 U879 ( .A(G290), .B(n901), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U881 ( .A(G166), .B(n792), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(G305), .ZN(n794) );
  XNOR2_X1 U883 ( .A(n795), .B(n794), .ZN(n887) );
  XNOR2_X1 U884 ( .A(n887), .B(n796), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n797), .A2(G868), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT85), .B(n798), .Z(n802) );
  NAND2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n802), .A2(n801), .ZN(G295) );
  NAND2_X1 U889 ( .A1(G2084), .A2(G2078), .ZN(n804) );
  XOR2_X1 U890 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n803) );
  XNOR2_X1 U891 ( .A(n804), .B(n803), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n805), .A2(G2090), .ZN(n806) );
  XOR2_X1 U893 ( .A(KEYINPUT21), .B(n806), .Z(n807) );
  XNOR2_X1 U894 ( .A(KEYINPUT87), .B(n807), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U896 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U897 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NAND2_X1 U898 ( .A1(G69), .A2(G120), .ZN(n809) );
  NOR2_X1 U899 ( .A1(G237), .A2(n809), .ZN(n810) );
  NAND2_X1 U900 ( .A1(G108), .A2(n810), .ZN(n899) );
  NAND2_X1 U901 ( .A1(n899), .A2(G567), .ZN(n816) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n811) );
  XNOR2_X1 U903 ( .A(KEYINPUT22), .B(n811), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n812), .A2(G96), .ZN(n813) );
  NOR2_X1 U905 ( .A1(G218), .A2(n813), .ZN(n814) );
  XOR2_X1 U906 ( .A(KEYINPUT88), .B(n814), .Z(n900) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n900), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n825) );
  NAND2_X1 U909 ( .A1(G661), .A2(G483), .ZN(n817) );
  XOR2_X1 U910 ( .A(KEYINPUT89), .B(n817), .Z(n818) );
  NOR2_X1 U911 ( .A1(n825), .A2(n818), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U913 ( .A1(n819), .A2(G2106), .ZN(n820) );
  XOR2_X1 U914 ( .A(KEYINPUT105), .B(n820), .Z(G217) );
  NAND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT106), .B(n821), .Z(n822) );
  NAND2_X1 U917 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(G188) );
  XNOR2_X1 U920 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  INV_X1 U921 ( .A(n825), .ZN(G319) );
  XOR2_X1 U922 ( .A(KEYINPUT110), .B(G1981), .Z(n827) );
  XNOR2_X1 U923 ( .A(G1966), .B(G1961), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U925 ( .A(n828), .B(KEYINPUT41), .Z(n830) );
  XNOR2_X1 U926 ( .A(G1996), .B(G1991), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U928 ( .A(G1976), .B(G1971), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1986), .B(G1956), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U931 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U932 ( .A(KEYINPUT109), .B(G2474), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(G229) );
  XOR2_X1 U934 ( .A(G2096), .B(KEYINPUT43), .Z(n838) );
  XNOR2_X1 U935 ( .A(G2072), .B(G2678), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U937 ( .A(n839), .B(KEYINPUT108), .Z(n841) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2090), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2100), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2078), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(G227) );
  NAND2_X1 U944 ( .A1(G136), .A2(n862), .ZN(n847) );
  NAND2_X1 U945 ( .A1(G112), .A2(n867), .ZN(n846) );
  NAND2_X1 U946 ( .A1(n847), .A2(n846), .ZN(n852) );
  NAND2_X1 U947 ( .A1(G124), .A2(n870), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n863), .A2(G100), .ZN(n849) );
  NAND2_X1 U950 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U951 ( .A1(n852), .A2(n851), .ZN(G162) );
  NAND2_X1 U952 ( .A1(G139), .A2(n862), .ZN(n854) );
  NAND2_X1 U953 ( .A1(G103), .A2(n863), .ZN(n853) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G115), .A2(n867), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G127), .A2(n870), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U958 ( .A(KEYINPUT47), .B(n857), .Z(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n906) );
  XNOR2_X1 U960 ( .A(G160), .B(n906), .ZN(n883) );
  XNOR2_X1 U961 ( .A(G162), .B(n860), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(n917), .ZN(n879) );
  XNOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n877) );
  NAND2_X1 U964 ( .A1(G142), .A2(n862), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G106), .A2(n863), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT45), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G118), .A2(n867), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G130), .A2(n870), .ZN(n871) );
  XNOR2_X1 U971 ( .A(KEYINPUT111), .B(n871), .ZN(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U976 ( .A(G164), .B(KEYINPUT48), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n883), .B(n882), .ZN(n885) );
  XNOR2_X1 U979 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U980 ( .A1(G37), .A2(n886), .ZN(G395) );
  XNOR2_X1 U981 ( .A(n887), .B(n961), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n888), .B(G286), .ZN(n890) );
  XOR2_X1 U983 ( .A(n963), .B(G171), .Z(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U985 ( .A1(G37), .A2(n891), .ZN(G397) );
  NOR2_X1 U986 ( .A1(G229), .A2(G227), .ZN(n893) );
  XNOR2_X1 U987 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n896) );
  NOR2_X1 U989 ( .A1(G395), .A2(G397), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(KEYINPUT114), .ZN(n895) );
  NAND2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G401), .A2(n897), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G319), .A2(n898), .ZN(G225) );
  XNOR2_X1 U994 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U996 ( .A(G120), .ZN(G236) );
  INV_X1 U997 ( .A(G69), .ZN(G235) );
  NOR2_X1 U998 ( .A1(n900), .A2(n899), .ZN(G325) );
  INV_X1 U999 ( .A(G325), .ZN(G261) );
  INV_X1 U1000 ( .A(G108), .ZN(G238) );
  INV_X1 U1001 ( .A(n901), .ZN(G299) );
  XOR2_X1 U1002 ( .A(G2090), .B(G162), .Z(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT51), .B(n904), .Z(n925) );
  XNOR2_X1 U1005 ( .A(G164), .B(G2078), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n905), .B(KEYINPUT117), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n906), .B(G2072), .Z(n907) );
  NOR2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT50), .B(n909), .ZN(n914) );
  INV_X1 U1010 ( .A(n910), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n923) );
  XOR2_X1 U1013 ( .A(G160), .B(G2084), .Z(n915) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1017 ( .A(KEYINPUT116), .B(n921), .Z(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(KEYINPUT52), .B(n926), .ZN(n927) );
  NAND2_X1 U1021 ( .A1(n927), .A2(G29), .ZN(n1010) );
  XNOR2_X1 U1022 ( .A(n928), .B(G27), .ZN(n931) );
  XNOR2_X1 U1023 ( .A(n929), .B(G32), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1025 ( .A(KEYINPUT119), .B(n932), .ZN(n938) );
  XOR2_X1 U1026 ( .A(G2072), .B(G33), .Z(n933) );
  NAND2_X1 U1027 ( .A1(n933), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(KEYINPUT118), .B(G2067), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G26), .B(n934), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(G25), .B(G1991), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1034 ( .A(KEYINPUT53), .B(n941), .Z(n944) );
  XOR2_X1 U1035 ( .A(KEYINPUT54), .B(G34), .Z(n942) );
  XNOR2_X1 U1036 ( .A(G2084), .B(n942), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G35), .B(G2090), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(KEYINPUT120), .ZN(n948) );
  NOR2_X1 U1041 ( .A1(G29), .A2(n948), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT55), .B(n949), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(G11), .ZN(n1008) );
  XNOR2_X1 U1044 ( .A(G16), .B(KEYINPUT56), .ZN(n978) );
  XNOR2_X1 U1045 ( .A(G171), .B(G1961), .ZN(n976) );
  XNOR2_X1 U1046 ( .A(G299), .B(G1956), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G303), .B(G1971), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n959) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT122), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT123), .ZN(n968) );
  XNOR2_X1 U1054 ( .A(G1341), .B(KEYINPUT124), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(n961), .ZN(n966) );
  INV_X1 U1056 ( .A(n963), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G1348), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n974) );
  XOR2_X1 U1060 ( .A(G1966), .B(G168), .Z(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n971), .Z(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT121), .B(n972), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n1006) );
  INV_X1 U1067 ( .A(G16), .ZN(n1004) );
  XNOR2_X1 U1068 ( .A(G5), .B(n979), .ZN(n999) );
  XOR2_X1 U1069 ( .A(KEYINPUT127), .B(KEYINPUT58), .Z(n986) );
  XNOR2_X1 U1070 ( .A(G1986), .B(G24), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(G23), .B(G1976), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1073 ( .A(G1971), .B(KEYINPUT126), .Z(n982) );
  XNOR2_X1 U1074 ( .A(G22), .B(n982), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n986), .B(n985), .ZN(n997) );
  XNOR2_X1 U1077 ( .A(G1956), .B(G20), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G1341), .B(G19), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(G1981), .B(G6), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n989), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(G4), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(KEYINPUT60), .B(n995), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G21), .B(G1966), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT61), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(KEYINPUT62), .B(n1011), .Z(G311) );
  INV_X1 U1097 ( .A(G311), .ZN(G150) );
endmodule

