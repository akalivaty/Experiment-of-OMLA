//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n213), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n208), .A2(new_n210), .A3(new_n212), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT67), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(G169gat), .A3(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n217), .A2(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(G169gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n221), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n215), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT25), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n225), .A2(new_n231), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n225), .A2(new_n231), .A3(new_n233), .ZN(new_n235));
  NOR2_X1   g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n209), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n235), .A2(KEYINPUT66), .B1(new_n237), .B2(new_n211), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n228), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n219), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI22_X1  g044(.A1(new_n243), .A2(new_n245), .B1(new_n204), .B2(new_n206), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT28), .ZN(new_n247));
  NOR2_X1   g046(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n205), .A2(new_n207), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n249), .B2(KEYINPUT27), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(G190gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT27), .B(G183gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(KEYINPUT28), .A3(new_n206), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n246), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n202), .B1(new_n240), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G127gat), .ZN(new_n257));
  INV_X1    g056(.A(G127gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G120gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT27), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n248), .ZN(new_n275));
  AOI21_X1  g074(.A(G190gat), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n253), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n241), .B(KEYINPUT26), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(new_n244), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(new_n228), .A3(KEYINPUT70), .A4(new_n239), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n255), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n283), .B(KEYINPUT64), .Z(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n228), .A3(new_n239), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n262), .A2(new_n270), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n202), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n282), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT33), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G15gat), .B(G43gat), .Z(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n288), .B(KEYINPUT32), .C1(new_n290), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n284), .A2(KEYINPUT34), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(new_n282), .B2(new_n287), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n271), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n235), .A2(KEYINPUT66), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n237), .A2(new_n211), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n302), .A2(new_n234), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n304), .A2(new_n230), .B1(new_n227), .B2(KEYINPUT25), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT70), .B1(new_n305), .B2(new_n280), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n287), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n283), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n300), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n298), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT72), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT31), .B(G50gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n322));
  XNOR2_X1  g121(.A(G155gat), .B(G162gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G141gat), .B(G148gat), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G148gat), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G141gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n321), .B(new_n331), .C1(new_n334), .C2(KEYINPUT76), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G211gat), .B(G218gat), .ZN(new_n339));
  INV_X1    g138(.A(G218gat), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT73), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G211gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n338), .B(new_n339), .C1(new_n345), .C2(KEYINPUT22), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT22), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT73), .B(G211gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(new_n340), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n339), .B1(new_n350), .B2(new_n338), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n337), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n336), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G228gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n336), .B2(new_n353), .ZN(new_n359));
  INV_X1    g158(.A(new_n339), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n344), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT22), .B1(new_n361), .B2(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n338), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n346), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n357), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(new_n354), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n336), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n364), .B2(new_n346), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(KEYINPUT3), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n347), .A2(new_n351), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n326), .B2(new_n335), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n358), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(new_n357), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G22gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n357), .ZN(new_n378));
  INV_X1    g177(.A(new_n358), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n365), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n336), .B1(new_n380), .B2(new_n353), .ZN(new_n381));
  INV_X1    g180(.A(new_n374), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n376), .A2(new_n377), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n377), .B1(new_n376), .B2(new_n383), .ZN(new_n385));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n386), .B(KEYINPUT79), .Z(new_n387));
  NOR3_X1   g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n354), .A2(new_n366), .A3(KEYINPUT80), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n336), .A2(new_n353), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n379), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n378), .B1(new_n392), .B2(new_n372), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n371), .B1(new_n393), .B2(new_n370), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n383), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G22gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n377), .A3(new_n383), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n319), .B1(new_n388), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n295), .A2(new_n297), .A3(new_n311), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n387), .B1(new_n384), .B2(new_n385), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n389), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n318), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G1gat), .B(G29gat), .Z(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT0), .ZN(new_n406));
  XNOR2_X1  g205(.A(G57gat), .B(G85gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n286), .A2(new_n336), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n271), .A2(new_n335), .A3(new_n326), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT5), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n410), .B2(new_n411), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT5), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT78), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n271), .B1(new_n336), .B2(new_n353), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(new_n373), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n414), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n286), .B2(new_n336), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n271), .B1(new_n335), .B2(new_n326), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(KEYINPUT4), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n417), .A2(new_n420), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n286), .A2(new_n336), .A3(new_n424), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n426), .B2(KEYINPUT4), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n431), .A2(new_n423), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n409), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n421), .A2(new_n373), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n427), .A2(new_n434), .A3(new_n413), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n416), .B1(new_n415), .B2(KEYINPUT5), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n418), .A2(KEYINPUT78), .A3(new_n419), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n423), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n408), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT6), .B(new_n409), .C1(new_n428), .C2(new_n432), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(G8gat), .B(G36gat), .Z(new_n445));
  XOR2_X1   g244(.A(G64gat), .B(G92gat), .Z(new_n446));
  XOR2_X1   g245(.A(new_n445), .B(new_n446), .Z(new_n447));
  XOR2_X1   g246(.A(new_n447), .B(KEYINPUT75), .Z(new_n448));
  OAI21_X1  g247(.A(new_n379), .B1(new_n240), .B2(new_n254), .ZN(new_n449));
  NAND2_X1  g248(.A1(G226gat), .A2(G233gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n285), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n365), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n285), .B2(new_n337), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n450), .B1(new_n305), .B2(new_n280), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(new_n372), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n448), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n452), .B1(new_n285), .B2(new_n379), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n372), .B1(new_n459), .B2(new_n456), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT29), .B1(new_n305), .B2(new_n280), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n453), .B(new_n365), .C1(new_n461), .C2(new_n452), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n447), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT30), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT30), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n317), .A2(new_n404), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n458), .B2(new_n463), .ZN(new_n471));
  INV_X1    g270(.A(new_n467), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n313), .A2(new_n473), .A3(new_n470), .A4(new_n444), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n469), .A2(new_n470), .B1(new_n404), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n400), .A2(KEYINPUT36), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n314), .A2(new_n476), .A3(new_n316), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT36), .B1(new_n313), .B2(new_n400), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n401), .A2(new_n402), .A3(new_n318), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n318), .B1(new_n401), .B2(new_n402), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n468), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n442), .A2(new_n443), .A3(new_n463), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n486), .A3(new_n462), .ZN(new_n487));
  INV_X1    g286(.A(new_n447), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT37), .B1(new_n454), .B2(new_n457), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n448), .A2(new_n485), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n365), .B1(new_n459), .B2(new_n456), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n453), .B(new_n372), .C1(new_n461), .C2(new_n452), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT37), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT82), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT82), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(new_n495), .A3(new_n498), .A4(KEYINPUT37), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n484), .A2(new_n491), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n414), .C1(new_n430), .C2(new_n422), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n503), .A2(new_n408), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT39), .B1(new_n412), .B2(new_n414), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n414), .B1(new_n430), .B2(new_n422), .ZN(new_n508));
  OAI211_X1 g307(.A(KEYINPUT81), .B(KEYINPUT39), .C1(new_n412), .C2(new_n414), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(KEYINPUT40), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT40), .B1(new_n504), .B2(new_n510), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n408), .B1(new_n438), .B2(new_n439), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n511), .B(new_n514), .C1(new_n471), .C2(new_n472), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n399), .A2(new_n515), .A3(new_n403), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n480), .B(new_n483), .C1(new_n501), .C2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n475), .A2(KEYINPUT83), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT83), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n404), .A2(new_n474), .ZN(new_n520));
  AOI211_X1 g319(.A(KEYINPUT72), .B(new_n311), .C1(new_n295), .C2(new_n297), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n315), .B1(new_n298), .B2(new_n312), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n481), .A2(new_n482), .ZN(new_n524));
  INV_X1    g323(.A(new_n468), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n400), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n520), .B1(new_n526), .B2(KEYINPUT35), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n478), .B1(new_n523), .B2(new_n476), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n483), .B1(new_n516), .B2(new_n501), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n519), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n518), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT16), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(G1gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(G1gat), .B2(new_n534), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G8gat), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n536), .B(new_n539), .C1(G1gat), .C2(new_n534), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n544), .A2(new_n546), .A3(KEYINPUT15), .A4(new_n547), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n541), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n553), .A2(new_n554), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT86), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n538), .A2(new_n540), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n555), .A2(new_n560), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT85), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n533), .B(new_n556), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT87), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n563), .A2(new_n570), .A3(new_n557), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT87), .B1(new_n541), .B2(new_n555), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n556), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n533), .B(KEYINPUT13), .Z(new_n574));
  AOI21_X1  g373(.A(KEYINPUT88), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n573), .A2(KEYINPUT88), .A3(new_n574), .ZN(new_n576));
  OAI22_X1  g375(.A1(new_n575), .A2(new_n576), .B1(new_n567), .B2(new_n568), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n569), .B1(new_n577), .B2(KEYINPUT89), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n565), .B(KEYINPUT85), .Z(new_n579));
  AOI21_X1  g378(.A(new_n541), .B1(new_n558), .B2(new_n561), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n579), .A2(new_n580), .B1(new_n541), .B2(new_n555), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(KEYINPUT18), .A3(new_n533), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n573), .A2(new_n574), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n573), .A2(KEYINPUT88), .A3(new_n574), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G197gat), .ZN(new_n592));
  XOR2_X1   g391(.A(KEYINPUT11), .B(G169gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n587), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n567), .A2(new_n600), .A3(new_n568), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n600), .B1(new_n567), .B2(new_n568), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G64gat), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n605), .A2(G57gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(G57gat), .ZN(new_n607));
  AND2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  OAI22_X1  g407(.A1(new_n606), .A2(new_n607), .B1(KEYINPUT9), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G71gat), .B(G78gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT20), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT94), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n541), .B1(KEYINPUT21), .B2(new_n611), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT93), .Z(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n630), .B(new_n631), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n625), .A3(new_n627), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  XNOR2_X1  g437(.A(G99gat), .B(G106gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(G85gat), .A2(G92gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT7), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT95), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  INV_X1    g442(.A(G85gat), .ZN(new_n644));
  INV_X1    g443(.A(G92gat), .ZN(new_n645));
  AOI22_X1  g444(.A1(KEYINPUT8), .A2(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n642), .B1(new_n641), .B2(new_n646), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n639), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  INV_X1    g450(.A(new_n639), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n611), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n650), .A2(new_n612), .A3(new_n653), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n654), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n638), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n638), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n655), .B2(new_n657), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n660), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n660), .B2(new_n662), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT98), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n670), .B(new_n666), .C1(new_n660), .C2(new_n662), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n654), .A2(new_n555), .ZN(new_n674));
  NAND3_X1  g473(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n562), .A2(new_n653), .A3(new_n650), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n674), .B(new_n675), .C1(new_n676), .C2(new_n566), .ZN(new_n677));
  XOR2_X1   g476(.A(G190gat), .B(G218gat), .Z(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  XNOR2_X1  g479(.A(G134gat), .B(G162gat), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n679), .A2(new_n680), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n680), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n677), .A2(new_n678), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n691), .B2(new_n684), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n636), .A2(new_n673), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n532), .A2(new_n604), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n444), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g497(.A1(new_n465), .A2(new_n467), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT16), .B(G8gat), .Z(new_n700));
  NAND3_X1  g499(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT42), .ZN(new_n702));
  OAI21_X1  g501(.A(G8gat), .B1(new_n694), .B2(new_n473), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(G1325gat));
  OAI21_X1  g506(.A(G15gat), .B1(new_n694), .B2(new_n480), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n313), .A2(new_n400), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(G15gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n694), .B2(new_n710), .ZN(G1326gat));
  NOR2_X1   g510(.A1(new_n694), .A2(new_n524), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  AOI21_X1  g513(.A(new_n598), .B1(new_n578), .B2(new_n589), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n636), .A2(new_n672), .A3(new_n692), .ZN(new_n718));
  AOI211_X1 g517(.A(new_n717), .B(new_n718), .C1(new_n518), .C2(new_n531), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n719), .A2(new_n542), .A3(new_n696), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT45), .ZN(new_n721));
  INV_X1    g520(.A(new_n692), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n518), .B2(new_n531), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n475), .A2(new_n517), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT44), .B1(new_n727), .B2(new_n692), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n636), .B(KEYINPUT100), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n604), .A3(new_n672), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n444), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT45), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n735), .A3(new_n736), .ZN(G1328gat));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n543), .A3(new_n699), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT101), .B(KEYINPUT46), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G36gat), .B1(new_n734), .B2(new_n473), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n739), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(G1329gat));
  AND4_X1   g542(.A1(G43gat), .A2(new_n729), .A3(new_n528), .A4(new_n733), .ZN(new_n744));
  INV_X1    g543(.A(new_n709), .ZN(new_n745));
  AOI21_X1  g544(.A(G43gat), .B1(new_n719), .B2(new_n745), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT47), .B1(new_n744), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1330gat));
  OAI21_X1  g548(.A(G50gat), .B1(new_n734), .B2(new_n524), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n524), .A2(G50gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n719), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n750), .A2(KEYINPUT102), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n751), .A2(KEYINPUT102), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(KEYINPUT102), .ZN(new_n756));
  INV_X1    g555(.A(G50gat), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n726), .A2(new_n728), .A3(new_n732), .ZN(new_n758));
  INV_X1    g557(.A(new_n524), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n753), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n755), .B(new_n756), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n754), .A2(new_n762), .ZN(G1331gat));
  NOR3_X1   g562(.A1(new_n604), .A2(new_n636), .A3(new_n692), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n727), .A2(new_n673), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(new_n444), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n765), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n699), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT49), .B(G64gat), .Z(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(G71gat), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n480), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n765), .B2(new_n709), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n769), .A2(new_n759), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT104), .B(G78gat), .Z(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1335gat));
  INV_X1    g581(.A(new_n636), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT105), .B1(new_n604), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n717), .A2(new_n785), .A3(new_n636), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n672), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT106), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n729), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n444), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n784), .A2(new_n786), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n692), .B(new_n792), .C1(new_n527), .C2(new_n530), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT108), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n722), .B1(new_n475), .B2(new_n517), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT51), .A4(new_n792), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT107), .B1(new_n793), .B2(new_n794), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n673), .A2(new_n644), .A3(new_n696), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n791), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  AOI21_X1  g603(.A(KEYINPUT83), .B1(new_n475), .B2(new_n517), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n527), .A2(new_n530), .A3(new_n519), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n724), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n527), .A2(new_n530), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n723), .B1(new_n808), .B2(new_n722), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n807), .A2(new_n699), .A3(new_n809), .A4(new_n789), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(new_n810), .B2(G92gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n672), .A2(new_n473), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(G92gat), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n802), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n810), .A2(KEYINPUT109), .A3(G92gat), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT109), .B1(new_n810), .B2(G92gat), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n814), .B(KEYINPUT110), .Z(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n793), .A2(new_n820), .A3(new_n794), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n793), .B2(new_n794), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n819), .B1(new_n823), .B2(new_n801), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n817), .A2(new_n818), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n816), .B1(new_n825), .B2(new_n826), .ZN(G1337gat));
  OAI21_X1  g626(.A(G99gat), .B1(new_n790), .B2(new_n480), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n709), .A2(new_n672), .A3(G99gat), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT112), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n802), .B2(new_n830), .ZN(G1338gat));
  NOR3_X1   g630(.A1(new_n524), .A2(G106gat), .A3(new_n672), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT113), .Z(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n823), .B2(new_n801), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n729), .A2(new_n759), .A3(new_n789), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(G106gat), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(G106gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n833), .B1(new_n796), .B2(new_n801), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n836), .A2(new_n837), .B1(new_n839), .B2(new_n840), .ZN(G1339gat));
  NAND2_X1  g640(.A1(new_n764), .A2(new_n672), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n581), .A2(new_n533), .B1(new_n574), .B2(new_n573), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n594), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n594), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n603), .A2(new_n848), .A3(new_n692), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n658), .A2(new_n659), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n661), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n658), .A2(new_n659), .A3(new_n638), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n665), .B1(new_n660), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(KEYINPUT55), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n667), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(KEYINPUT114), .A3(new_n667), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n853), .A2(new_n855), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n673), .A2(new_n603), .A3(new_n848), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n717), .B2(new_n864), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(new_n722), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n842), .B1(new_n868), .B2(new_n730), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n759), .A2(new_n709), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n699), .A2(new_n444), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n265), .A3(new_n717), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n696), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n317), .A3(new_n404), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n604), .A3(new_n473), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(new_n877), .B2(new_n265), .ZN(G1340gat));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n473), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n673), .A2(new_n263), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n869), .A2(new_n673), .A3(new_n872), .A4(new_n870), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT116), .B1(new_n881), .B2(G120gat), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n879), .A2(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n884), .B(new_n885), .ZN(G1341gat));
  OAI21_X1  g685(.A(G127gat), .B1(new_n873), .B2(new_n731), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n783), .A2(new_n258), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n879), .B2(new_n888), .ZN(G1342gat));
  OAI21_X1  g688(.A(G134gat), .B1(new_n873), .B2(new_n722), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n722), .A2(new_n699), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n256), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT56), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n892), .B2(KEYINPUT56), .ZN(new_n895));
  OAI221_X1 g694(.A(new_n890), .B1(KEYINPUT56), .B2(new_n892), .C1(new_n894), .C2(new_n895), .ZN(G1343gat));
  INV_X1    g695(.A(new_n857), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n897), .B(new_n863), .C1(new_n715), .C2(new_n716), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n692), .B1(new_n898), .B2(new_n866), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n636), .B1(new_n899), .B2(new_n865), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n842), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n759), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT57), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n869), .A2(new_n904), .A3(new_n759), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n480), .A2(new_n872), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G141gat), .B1(new_n907), .B2(new_n717), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n528), .A2(new_n524), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n869), .A2(new_n696), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n699), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n717), .A2(G141gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT58), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n915));
  INV_X1    g714(.A(new_n905), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n524), .B1(new_n900), .B2(new_n842), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n906), .B1(new_n917), .B2(new_n904), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n903), .A2(KEYINPUT119), .A3(new_n905), .A4(new_n906), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n604), .A3(new_n920), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n921), .A2(G141gat), .B1(new_n911), .B2(new_n912), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n914), .B1(new_n922), .B2(new_n923), .ZN(G1344gat));
  NAND3_X1  g723(.A1(new_n911), .A2(new_n329), .A3(new_n673), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n673), .A3(new_n920), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n329), .A2(KEYINPUT59), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n902), .A2(new_n930), .A3(new_n904), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n869), .A2(KEYINPUT57), .A3(new_n759), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT120), .B1(new_n917), .B2(KEYINPUT57), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n673), .A3(new_n906), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n929), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n925), .B1(new_n928), .B2(new_n936), .ZN(G1345gat));
  INV_X1    g736(.A(G155gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n911), .A2(new_n938), .A3(new_n783), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n919), .A2(new_n730), .A3(new_n920), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n938), .ZN(G1346gat));
  AND3_X1   g740(.A1(new_n919), .A2(new_n692), .A3(new_n920), .ZN(new_n942));
  INV_X1    g741(.A(G162gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n891), .A2(new_n943), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n942), .A2(new_n943), .B1(new_n910), .B2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n696), .A2(new_n473), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT121), .ZN(new_n947));
  AND4_X1   g746(.A1(G169gat), .A2(new_n871), .A3(new_n604), .A4(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n869), .A2(new_n444), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n317), .A2(new_n404), .A3(new_n473), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n604), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n220), .B2(new_n952), .ZN(G1348gat));
  AOI21_X1  g752(.A(G176gat), .B1(new_n951), .B2(new_n673), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n672), .B1(new_n231), .B2(new_n233), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n871), .A2(new_n947), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(G1349gat));
  NAND4_X1  g759(.A1(new_n869), .A2(new_n730), .A3(new_n870), .A4(new_n947), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n961), .A2(KEYINPUT123), .B1(new_n205), .B2(new_n207), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(KEYINPUT123), .B2(new_n961), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n951), .A2(new_n252), .A3(new_n783), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n965), .B(new_n966), .ZN(G1350gat));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n206), .A3(new_n692), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n869), .A2(new_n692), .A3(new_n870), .A4(new_n947), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G190gat), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(G1351gat));
  NAND2_X1  g775(.A1(new_n947), .A2(new_n480), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT127), .Z(new_n978));
  NAND2_X1  g777(.A1(new_n934), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(G197gat), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n979), .A2(new_n980), .A3(new_n717), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n949), .A2(new_n699), .A3(new_n909), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT126), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(new_n604), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n981), .B1(new_n984), .B2(new_n980), .ZN(G1352gat));
  NOR2_X1   g784(.A1(new_n813), .A2(G204gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n949), .A2(new_n909), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT62), .Z(new_n988));
  OAI21_X1  g787(.A(G204gat), .B1(new_n979), .B2(new_n672), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1353gat));
  NAND3_X1  g789(.A1(new_n983), .A2(new_n349), .A3(new_n783), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n934), .A2(new_n783), .A3(new_n978), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n992), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  NAND3_X1  g794(.A1(new_n983), .A2(new_n340), .A3(new_n692), .ZN(new_n996));
  OAI21_X1  g795(.A(G218gat), .B1(new_n979), .B2(new_n722), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1355gat));
endmodule


