

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751;

  XNOR2_X1 U369 ( .A(n602), .B(n601), .ZN(n656) );
  XNOR2_X1 U370 ( .A(KEYINPUT96), .B(n599), .ZN(n641) );
  AND2_X1 U371 ( .A1(n395), .A2(n356), .ZN(n441) );
  XNOR2_X1 U372 ( .A(n506), .B(n386), .ZN(n385) );
  XNOR2_X1 U373 ( .A(G143), .B(G104), .ZN(n536) );
  XNOR2_X1 U374 ( .A(n412), .B(n410), .ZN(n506) );
  XNOR2_X1 U375 ( .A(KEYINPUT76), .B(G104), .ZN(n413) );
  NAND2_X1 U376 ( .A1(n370), .A2(n372), .ZN(n366) );
  AND2_X4 U377 ( .A1(n707), .A2(n706), .ZN(n458) );
  XNOR2_X2 U378 ( .A(n347), .B(n627), .ZN(n726) );
  NAND2_X1 U379 ( .A1(n464), .A2(n459), .ZN(n347) );
  XNOR2_X1 U380 ( .A(n606), .B(n607), .ZN(n695) );
  INV_X1 U381 ( .A(n548), .ZN(n614) );
  OR2_X2 U382 ( .A1(n708), .A2(G902), .ZN(n465) );
  NOR2_X2 U383 ( .A1(n416), .A2(n415), .ZN(n579) );
  NOR2_X2 U384 ( .A1(n588), .A2(n349), .ZN(n404) );
  XNOR2_X2 U385 ( .A(n511), .B(n456), .ZN(n530) );
  XNOR2_X2 U386 ( .A(n721), .B(n516), .ZN(n703) );
  XNOR2_X2 U387 ( .A(n385), .B(n504), .ZN(n721) );
  NOR2_X2 U388 ( .A1(n517), .A2(n703), .ZN(n522) );
  AND2_X1 U389 ( .A1(n401), .A2(n678), .ZN(n638) );
  AND2_X1 U390 ( .A1(n367), .A2(n594), .ZN(n659) );
  AND2_X1 U391 ( .A1(n613), .A2(n374), .ZN(n646) );
  XNOR2_X1 U392 ( .A(n375), .B(n360), .ZN(n620) );
  INV_X1 U393 ( .A(n596), .ZN(n608) );
  XNOR2_X1 U394 ( .A(n376), .B(KEYINPUT41), .ZN(n694) );
  XNOR2_X1 U395 ( .A(n404), .B(n358), .ZN(n596) );
  XNOR2_X1 U396 ( .A(n563), .B(KEYINPUT1), .ZN(n676) );
  XNOR2_X1 U397 ( .A(n500), .B(n501), .ZN(n635) );
  XNOR2_X1 U398 ( .A(n530), .B(G137), .ZN(n472) );
  XNOR2_X1 U399 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U400 ( .A(n505), .B(n409), .ZN(n386) );
  INV_X1 U401 ( .A(G122), .ZN(n505) );
  XNOR2_X1 U402 ( .A(G953), .B(KEYINPUT64), .ZN(n477) );
  INV_X2 U403 ( .A(G143), .ZN(n457) );
  NAND2_X2 U404 ( .A1(n633), .A2(n632), .ZN(n707) );
  INV_X1 U405 ( .A(KEYINPUT38), .ZN(n380) );
  NOR2_X1 U406 ( .A1(G953), .A2(G237), .ZN(n533) );
  OR2_X1 U407 ( .A1(n635), .A2(n443), .ZN(n442) );
  NAND2_X1 U408 ( .A1(n502), .A2(n444), .ZN(n443) );
  INV_X1 U409 ( .A(G902), .ZN(n444) );
  XNOR2_X1 U410 ( .A(n626), .B(KEYINPUT65), .ZN(n627) );
  XNOR2_X1 U411 ( .A(n454), .B(G140), .ZN(n453) );
  INV_X1 U412 ( .A(KEYINPUT10), .ZN(n454) );
  NAND2_X1 U413 ( .A1(n426), .A2(n351), .ZN(n428) );
  XNOR2_X1 U414 ( .A(n366), .B(KEYINPUT105), .ZN(n464) );
  XNOR2_X1 U415 ( .A(n497), .B(n498), .ZN(n504) );
  XNOR2_X1 U416 ( .A(n496), .B(KEYINPUT3), .ZN(n497) );
  XNOR2_X1 U417 ( .A(G116), .B(G119), .ZN(n496) );
  XNOR2_X1 U418 ( .A(n455), .B(G146), .ZN(n510) );
  INV_X1 U419 ( .A(G125), .ZN(n455) );
  XNOR2_X1 U420 ( .A(n411), .B(G101), .ZN(n410) );
  XNOR2_X1 U421 ( .A(n413), .B(n474), .ZN(n412) );
  INV_X1 U422 ( .A(G107), .ZN(n411) );
  INV_X1 U423 ( .A(KEYINPUT6), .ZN(n394) );
  XOR2_X1 U424 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n480) );
  XNOR2_X1 U425 ( .A(G128), .B(G119), .ZN(n481) );
  XOR2_X1 U426 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n483) );
  INV_X1 U427 ( .A(G134), .ZN(n456) );
  XNOR2_X1 U428 ( .A(n452), .B(n542), .ZN(n543) );
  AND2_X1 U429 ( .A1(n393), .A2(n391), .ZN(n664) );
  AND2_X1 U430 ( .A1(n750), .A2(n392), .ZN(n391) );
  INV_X1 U431 ( .A(n661), .ZN(n392) );
  NAND2_X1 U432 ( .A1(n431), .A2(n357), .ZN(n430) );
  OR2_X1 U433 ( .A1(n433), .A2(n550), .ZN(n431) );
  NAND2_X1 U434 ( .A1(n583), .A2(n669), .ZN(n558) );
  NAND2_X1 U435 ( .A1(n608), .A2(n381), .ZN(n375) );
  AND2_X1 U436 ( .A1(n593), .A2(n348), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n600), .B(KEYINPUT97), .ZN(n685) );
  NAND2_X1 U438 ( .A1(n369), .A2(n598), .ZN(n503) );
  XNOR2_X1 U439 ( .A(n561), .B(n389), .ZN(n562) );
  XNOR2_X1 U440 ( .A(n390), .B(KEYINPUT28), .ZN(n389) );
  INV_X1 U441 ( .A(n616), .ZN(n403) );
  NOR2_X1 U442 ( .A1(n620), .A2(n594), .ZN(n613) );
  INV_X1 U443 ( .A(KEYINPUT103), .ZN(n371) );
  XNOR2_X1 U444 ( .A(G113), .B(KEYINPUT93), .ZN(n495) );
  INV_X1 U445 ( .A(G110), .ZN(n474) );
  INV_X1 U446 ( .A(n746), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n569), .B(n418), .ZN(n417) );
  INV_X1 U448 ( .A(KEYINPUT84), .ZN(n418) );
  NAND2_X1 U449 ( .A1(n669), .A2(KEYINPUT30), .ZN(n440) );
  OR2_X1 U450 ( .A1(G902), .A2(G237), .ZN(n518) );
  NAND2_X1 U451 ( .A1(n748), .A2(KEYINPUT44), .ZN(n373) );
  INV_X1 U452 ( .A(KEYINPUT16), .ZN(n409) );
  XOR2_X1 U453 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n535) );
  XNOR2_X1 U454 ( .A(G122), .B(G113), .ZN(n541) );
  XOR2_X1 U455 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n537) );
  XNOR2_X1 U456 ( .A(G902), .B(KEYINPUT15), .ZN(n630) );
  XOR2_X1 U457 ( .A(KEYINPUT17), .B(KEYINPUT78), .Z(n508) );
  NAND2_X1 U458 ( .A1(G237), .A2(G234), .ZN(n468) );
  NOR2_X1 U459 ( .A1(n441), .A2(n440), .ZN(n436) );
  NAND2_X1 U460 ( .A1(n439), .A2(n438), .ZN(n437) );
  OR2_X1 U461 ( .A1(n669), .A2(KEYINPUT30), .ZN(n438) );
  OR2_X1 U462 ( .A1(n442), .A2(n440), .ZN(n439) );
  NOR2_X1 U463 ( .A1(n550), .A2(n549), .ZN(n560) );
  INV_X1 U464 ( .A(KEYINPUT109), .ZN(n390) );
  XOR2_X1 U465 ( .A(G101), .B(KEYINPUT5), .Z(n494) );
  INV_X1 U466 ( .A(G953), .ZN(n725) );
  XNOR2_X1 U467 ( .A(G122), .B(G116), .ZN(n523) );
  XNOR2_X1 U468 ( .A(n500), .B(n466), .ZN(n708) );
  XNOR2_X1 U469 ( .A(n475), .B(G140), .ZN(n476) );
  INV_X1 U470 ( .A(n666), .ZN(n451) );
  XNOR2_X1 U471 ( .A(n580), .B(n553), .ZN(n554) );
  INV_X1 U472 ( .A(KEYINPUT111), .ZN(n553) );
  XNOR2_X1 U473 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U474 ( .A(n484), .B(n483), .ZN(n485) );
  AND2_X1 U475 ( .A1(n388), .A2(n350), .ZN(n665) );
  NOR2_X1 U476 ( .A1(n425), .A2(n427), .ZN(n578) );
  NAND2_X1 U477 ( .A1(n428), .A2(n432), .ZN(n425) );
  NAND2_X1 U478 ( .A1(n430), .A2(n651), .ZN(n427) );
  INV_X1 U479 ( .A(KEYINPUT80), .ZN(n383) );
  NAND2_X1 U480 ( .A1(n608), .A2(n685), .ZN(n602) );
  NOR2_X1 U481 ( .A1(n588), .A2(n564), .ZN(n652) );
  NOR2_X1 U482 ( .A1(n683), .A2(n548), .ZN(n374) );
  NOR2_X1 U483 ( .A1(n596), .A2(n683), .ZN(n597) );
  XNOR2_X1 U484 ( .A(n402), .B(n595), .ZN(n401) );
  INV_X1 U485 ( .A(KEYINPUT88), .ZN(n595) );
  NAND2_X1 U486 ( .A1(n613), .A2(n403), .ZN(n402) );
  XNOR2_X1 U487 ( .A(n420), .B(KEYINPUT119), .ZN(G63) );
  NAND2_X1 U488 ( .A1(n422), .A2(n421), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n422) );
  INV_X1 U490 ( .A(KEYINPUT60), .ZN(n405) );
  NAND2_X1 U491 ( .A1(n407), .A2(n421), .ZN(n406) );
  XNOR2_X1 U492 ( .A(n408), .B(n363), .ZN(n407) );
  INV_X1 U493 ( .A(KEYINPUT56), .ZN(n447) );
  NAND2_X1 U494 ( .A1(n449), .A2(n421), .ZN(n448) );
  XNOR2_X1 U495 ( .A(n450), .B(n362), .ZN(n449) );
  XOR2_X1 U496 ( .A(KEYINPUT21), .B(n492), .Z(n348) );
  NOR2_X1 U497 ( .A1(n592), .A2(n591), .ZN(n349) );
  OR2_X1 U498 ( .A1(n664), .A2(n663), .ZN(n350) );
  AND2_X1 U499 ( .A1(n668), .A2(n429), .ZN(n351) );
  AND2_X1 U500 ( .A1(n706), .A2(G478), .ZN(n352) );
  OR2_X1 U501 ( .A1(n503), .A2(n550), .ZN(n353) );
  AND2_X1 U502 ( .A1(n428), .A2(n430), .ZN(n354) );
  AND2_X1 U503 ( .A1(n442), .A2(n445), .ZN(n355) );
  BUF_X1 U504 ( .A(n676), .Z(n382) );
  NAND2_X1 U505 ( .A1(n446), .A2(G902), .ZN(n356) );
  XOR2_X1 U506 ( .A(KEYINPUT74), .B(KEYINPUT39), .Z(n357) );
  XOR2_X1 U507 ( .A(KEYINPUT0), .B(KEYINPUT68), .Z(n358) );
  XOR2_X1 U508 ( .A(KEYINPUT72), .B(G469), .Z(n359) );
  XOR2_X1 U509 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n360) );
  XOR2_X1 U510 ( .A(n556), .B(n555), .Z(n361) );
  INV_X1 U511 ( .A(KEYINPUT30), .ZN(n445) );
  XOR2_X1 U512 ( .A(n705), .B(n704), .Z(n362) );
  XNOR2_X1 U513 ( .A(n714), .B(KEYINPUT59), .ZN(n363) );
  XNOR2_X1 U514 ( .A(n510), .B(n453), .ZN(n735) );
  INV_X1 U515 ( .A(n735), .ZN(n452) );
  XOR2_X1 U516 ( .A(n637), .B(n636), .Z(n364) );
  XOR2_X1 U517 ( .A(KEYINPUT63), .B(KEYINPUT113), .Z(n365) );
  INV_X1 U518 ( .A(n720), .ZN(n421) );
  XNOR2_X1 U519 ( .A(n603), .B(KEYINPUT98), .ZN(n400) );
  NAND2_X1 U520 ( .A1(n400), .A2(n565), .ZN(n399) );
  XNOR2_X1 U521 ( .A(n557), .B(n361), .ZN(n367) );
  AND2_X1 U522 ( .A1(n461), .A2(n460), .ZN(n459) );
  NOR2_X1 U523 ( .A1(n751), .A2(n646), .ZN(n624) );
  XNOR2_X1 U524 ( .A(n621), .B(KEYINPUT32), .ZN(n751) );
  NOR2_X1 U525 ( .A1(n618), .A2(n617), .ZN(n384) );
  NOR2_X1 U526 ( .A1(n624), .A2(n622), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n435), .A2(n434), .ZN(n369) );
  XNOR2_X1 U528 ( .A(n377), .B(KEYINPUT46), .ZN(n415) );
  INV_X1 U529 ( .A(n749), .ZN(n378) );
  NAND2_X1 U530 ( .A1(n656), .A2(n641), .ZN(n603) );
  XNOR2_X1 U531 ( .A(n399), .B(n371), .ZN(n370) );
  INV_X1 U532 ( .A(n638), .ZN(n372) );
  AND2_X1 U533 ( .A1(n625), .A2(n373), .ZN(n460) );
  NAND2_X1 U534 ( .A1(n695), .A2(n608), .ZN(n609) );
  NAND2_X1 U535 ( .A1(n451), .A2(n593), .ZN(n376) );
  NAND2_X1 U536 ( .A1(n379), .A2(n378), .ZN(n377) );
  NAND2_X1 U537 ( .A1(n668), .A2(n669), .ZN(n666) );
  XNOR2_X1 U538 ( .A(n583), .B(n380), .ZN(n668) );
  XNOR2_X2 U539 ( .A(n414), .B(G146), .ZN(n500) );
  NOR2_X1 U540 ( .A1(n554), .A2(n558), .ZN(n557) );
  XNOR2_X1 U541 ( .A(n384), .B(n383), .ZN(n619) );
  NOR2_X1 U542 ( .A1(n701), .A2(G953), .ZN(n702) );
  XNOR2_X1 U543 ( .A(n662), .B(KEYINPUT85), .ZN(n388) );
  XNOR2_X1 U544 ( .A(n387), .B(n490), .ZN(n548) );
  NOR2_X1 U545 ( .A1(n716), .A2(G902), .ZN(n387) );
  NOR2_X1 U546 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X2 U547 ( .A(n558), .B(n559), .ZN(n588) );
  XNOR2_X2 U548 ( .A(n683), .B(n394), .ZN(n616) );
  NAND2_X4 U549 ( .A1(n441), .A2(n442), .ZN(n683) );
  NAND2_X1 U550 ( .A1(n635), .A2(n446), .ZN(n395) );
  NAND2_X1 U551 ( .A1(n664), .A2(KEYINPUT2), .ZN(n587) );
  XNOR2_X1 U552 ( .A(n579), .B(KEYINPUT48), .ZN(n393) );
  XNOR2_X1 U553 ( .A(n396), .B(n365), .ZN(G57) );
  NAND2_X1 U554 ( .A1(n397), .A2(n421), .ZN(n396) );
  XNOR2_X1 U555 ( .A(n398), .B(n364), .ZN(n397) );
  NAND2_X1 U556 ( .A1(n634), .A2(n707), .ZN(n398) );
  XNOR2_X1 U557 ( .A(n406), .B(n405), .ZN(G60) );
  NAND2_X1 U558 ( .A1(n458), .A2(G475), .ZN(n408) );
  XNOR2_X1 U559 ( .A(n414), .B(n452), .ZN(n740) );
  XNOR2_X2 U560 ( .A(n472), .B(n473), .ZN(n414) );
  NAND2_X1 U561 ( .A1(n419), .A2(n417), .ZN(n416) );
  NOR2_X1 U562 ( .A1(n659), .A2(n571), .ZN(n419) );
  INV_X1 U563 ( .A(n715), .ZN(n423) );
  NAND2_X1 U564 ( .A1(n352), .A2(n707), .ZN(n424) );
  NAND2_X1 U565 ( .A1(n503), .A2(n357), .ZN(n432) );
  INV_X1 U566 ( .A(n503), .ZN(n426) );
  NAND2_X1 U567 ( .A1(n354), .A2(n432), .ZN(n577) );
  NOR2_X1 U568 ( .A1(n550), .A2(n357), .ZN(n429) );
  INV_X1 U569 ( .A(n668), .ZN(n433) );
  NAND2_X1 U570 ( .A1(n441), .A2(n355), .ZN(n434) );
  NOR2_X1 U571 ( .A1(n437), .A2(n436), .ZN(n435) );
  INV_X1 U572 ( .A(n502), .ZN(n446) );
  XNOR2_X1 U573 ( .A(n448), .B(n447), .ZN(G51) );
  NAND2_X1 U574 ( .A1(n458), .A2(G210), .ZN(n450) );
  INV_X1 U575 ( .A(n593), .ZN(n671) );
  NAND2_X1 U576 ( .A1(n574), .A2(n694), .ZN(n576) );
  XNOR2_X2 U577 ( .A(n457), .B(G128), .ZN(n511) );
  NAND2_X1 U578 ( .A1(n458), .A2(G469), .ZN(n711) );
  NAND2_X1 U579 ( .A1(n458), .A2(G217), .ZN(n717) );
  XNOR2_X1 U580 ( .A(n463), .B(n462), .ZN(n461) );
  INV_X1 U581 ( .A(KEYINPUT66), .ZN(n462) );
  XNOR2_X2 U582 ( .A(n465), .B(n359), .ZN(n563) );
  XNOR2_X1 U583 ( .A(n506), .B(n476), .ZN(n466) );
  XOR2_X1 U584 ( .A(KEYINPUT77), .B(KEYINPUT25), .Z(n467) );
  INV_X1 U585 ( .A(KEYINPUT112), .ZN(n555) );
  XNOR2_X1 U586 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U587 ( .A(n489), .B(n467), .ZN(n490) );
  INV_X1 U588 ( .A(KEYINPUT82), .ZN(n519) );
  NOR2_X1 U589 ( .A1(G952), .A2(n742), .ZN(n720) );
  INV_X1 U590 ( .A(n477), .ZN(n742) );
  XNOR2_X1 U591 ( .A(n468), .B(KEYINPUT14), .ZN(n469) );
  NAND2_X1 U592 ( .A1(G952), .A2(n469), .ZN(n693) );
  NOR2_X1 U593 ( .A1(G953), .A2(n693), .ZN(n592) );
  AND2_X1 U594 ( .A1(G902), .A2(n469), .ZN(n589) );
  NAND2_X1 U595 ( .A1(n477), .A2(n589), .ZN(n470) );
  NOR2_X1 U596 ( .A1(G900), .A2(n470), .ZN(n471) );
  NOR2_X1 U597 ( .A1(n592), .A2(n471), .ZN(n550) );
  XOR2_X1 U598 ( .A(KEYINPUT71), .B(G131), .Z(n540) );
  XOR2_X1 U599 ( .A(KEYINPUT4), .B(KEYINPUT69), .Z(n509) );
  XOR2_X1 U600 ( .A(n540), .B(n509), .Z(n473) );
  NAND2_X1 U601 ( .A1(G227), .A2(n742), .ZN(n475) );
  INV_X1 U602 ( .A(G234), .ZN(n478) );
  OR2_X1 U603 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U604 ( .A(n480), .B(n479), .ZN(n525) );
  NAND2_X1 U605 ( .A1(G221), .A2(n525), .ZN(n486) );
  XOR2_X1 U606 ( .A(G137), .B(G110), .Z(n482) );
  XNOR2_X1 U607 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U608 ( .A(n487), .B(n735), .ZN(n716) );
  NAND2_X1 U609 ( .A1(G234), .A2(n630), .ZN(n488) );
  XNOR2_X1 U610 ( .A(KEYINPUT20), .B(n488), .ZN(n491) );
  NAND2_X1 U611 ( .A1(n491), .A2(G217), .ZN(n489) );
  NAND2_X1 U612 ( .A1(n491), .A2(G221), .ZN(n492) );
  NAND2_X1 U613 ( .A1(n548), .A2(n348), .ZN(n675) );
  NOR2_X1 U614 ( .A1(n563), .A2(n675), .ZN(n598) );
  XNOR2_X1 U615 ( .A(KEYINPUT95), .B(G472), .ZN(n502) );
  NAND2_X1 U616 ( .A1(n533), .A2(G210), .ZN(n493) );
  XNOR2_X1 U617 ( .A(n494), .B(n493), .ZN(n499) );
  XNOR2_X1 U618 ( .A(n495), .B(KEYINPUT73), .ZN(n498) );
  XNOR2_X1 U619 ( .A(n499), .B(n504), .ZN(n501) );
  NAND2_X1 U620 ( .A1(G214), .A2(n518), .ZN(n669) );
  INV_X1 U621 ( .A(n630), .ZN(n517) );
  NAND2_X1 U622 ( .A1(G224), .A2(n742), .ZN(n507) );
  XNOR2_X1 U623 ( .A(n508), .B(n507), .ZN(n515) );
  XOR2_X1 U624 ( .A(KEYINPUT18), .B(n509), .Z(n513) );
  XNOR2_X1 U625 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U626 ( .A(n513), .B(n512), .ZN(n514) );
  AND2_X1 U627 ( .A1(G210), .A2(n518), .ZN(n520) );
  XNOR2_X2 U628 ( .A(n522), .B(n521), .ZN(n583) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(G107), .Z(n524) );
  XNOR2_X1 U630 ( .A(n524), .B(n523), .ZN(n529) );
  XOR2_X1 U631 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n527) );
  NAND2_X1 U632 ( .A1(G217), .A2(n525), .ZN(n526) );
  XNOR2_X1 U633 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U634 ( .A(n529), .B(n528), .ZN(n531) );
  XNOR2_X1 U635 ( .A(n530), .B(n531), .ZN(n715) );
  NOR2_X1 U636 ( .A1(n715), .A2(G902), .ZN(n532) );
  XNOR2_X1 U637 ( .A(G478), .B(n532), .ZN(n566) );
  XNOR2_X1 U638 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n546) );
  NAND2_X1 U639 ( .A1(G214), .A2(n533), .ZN(n534) );
  XNOR2_X1 U640 ( .A(n535), .B(n534), .ZN(n539) );
  XNOR2_X1 U641 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U642 ( .A(n539), .B(n538), .Z(n544) );
  XNOR2_X1 U643 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U644 ( .A(n544), .B(n543), .ZN(n714) );
  NOR2_X1 U645 ( .A1(G902), .A2(n714), .ZN(n545) );
  XNOR2_X1 U646 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U647 ( .A(G475), .B(n547), .Z(n572) );
  NOR2_X1 U648 ( .A1(n566), .A2(n572), .ZN(n647) );
  INV_X1 U649 ( .A(n647), .ZN(n657) );
  NOR2_X1 U650 ( .A1(n577), .A2(n657), .ZN(n661) );
  NAND2_X1 U651 ( .A1(n614), .A2(n348), .ZN(n549) );
  NAND2_X1 U652 ( .A1(n616), .A2(n560), .ZN(n551) );
  XNOR2_X1 U653 ( .A(n551), .B(KEYINPUT107), .ZN(n552) );
  NAND2_X1 U654 ( .A1(n566), .A2(n572), .ZN(n654) );
  INV_X1 U655 ( .A(n654), .ZN(n651) );
  NAND2_X1 U656 ( .A1(n552), .A2(n651), .ZN(n580) );
  XOR2_X1 U657 ( .A(KEYINPUT36), .B(KEYINPUT89), .Z(n556) );
  XNOR2_X1 U658 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n559) );
  NAND2_X1 U659 ( .A1(n560), .A2(n683), .ZN(n561) );
  NOR2_X1 U660 ( .A1(n563), .A2(n562), .ZN(n574) );
  INV_X1 U661 ( .A(n574), .ZN(n564) );
  NOR2_X1 U662 ( .A1(n651), .A2(n647), .ZN(n667) );
  INV_X1 U663 ( .A(n667), .ZN(n565) );
  NAND2_X1 U664 ( .A1(n652), .A2(n565), .ZN(n570) );
  NAND2_X1 U665 ( .A1(n570), .A2(KEYINPUT47), .ZN(n568) );
  INV_X1 U666 ( .A(n566), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n573), .A2(n572), .ZN(n604) );
  NOR2_X1 U668 ( .A1(n604), .A2(n353), .ZN(n567) );
  NAND2_X1 U669 ( .A1(n567), .A2(n583), .ZN(n650) );
  NAND2_X1 U670 ( .A1(n568), .A2(n650), .ZN(n569) );
  NOR2_X1 U671 ( .A1(KEYINPUT47), .A2(n570), .ZN(n571) );
  NOR2_X1 U672 ( .A1(n573), .A2(n572), .ZN(n593) );
  XOR2_X1 U673 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n575) );
  XNOR2_X1 U674 ( .A(n576), .B(n575), .ZN(n746) );
  XNOR2_X1 U675 ( .A(n578), .B(KEYINPUT40), .ZN(n749) );
  INV_X1 U676 ( .A(n382), .ZN(n594) );
  NOR2_X1 U677 ( .A1(n594), .A2(n580), .ZN(n581) );
  NAND2_X1 U678 ( .A1(n581), .A2(n669), .ZN(n582) );
  XNOR2_X1 U679 ( .A(KEYINPUT43), .B(n582), .ZN(n585) );
  INV_X1 U680 ( .A(n583), .ZN(n584) );
  NAND2_X1 U681 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U682 ( .A(KEYINPUT108), .B(n586), .ZN(n750) );
  XNOR2_X1 U683 ( .A(n587), .B(KEYINPUT87), .ZN(n628) );
  XOR2_X1 U684 ( .A(KEYINPUT104), .B(n614), .Z(n678) );
  NOR2_X1 U685 ( .A1(G898), .A2(n725), .ZN(n722) );
  NAND2_X1 U686 ( .A1(n722), .A2(n589), .ZN(n590) );
  XOR2_X1 U687 ( .A(KEYINPUT94), .B(n590), .Z(n591) );
  NAND2_X1 U688 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U689 ( .A1(n676), .A2(n675), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n605), .A2(n683), .ZN(n600) );
  INV_X1 U691 ( .A(KEYINPUT31), .ZN(n601) );
  XNOR2_X1 U692 ( .A(n604), .B(KEYINPUT79), .ZN(n611) );
  XOR2_X1 U693 ( .A(KEYINPUT91), .B(KEYINPUT33), .Z(n607) );
  NAND2_X1 U694 ( .A1(n605), .A2(n616), .ZN(n606) );
  XOR2_X1 U695 ( .A(KEYINPUT34), .B(n609), .Z(n610) );
  NAND2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U697 ( .A(n612), .B(KEYINPUT35), .ZN(n748) );
  NOR2_X1 U698 ( .A1(n678), .A2(n676), .ZN(n615) );
  XOR2_X1 U699 ( .A(KEYINPUT106), .B(n615), .Z(n618) );
  XOR2_X1 U700 ( .A(n616), .B(KEYINPUT81), .Z(n617) );
  INV_X1 U701 ( .A(KEYINPUT44), .ZN(n622) );
  NOR2_X1 U702 ( .A1(KEYINPUT44), .A2(n748), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U704 ( .A(KEYINPUT45), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n628), .A2(n726), .ZN(n706) );
  AND2_X1 U706 ( .A1(G472), .A2(n706), .ZN(n634) );
  INV_X1 U707 ( .A(n664), .ZN(n741) );
  NOR2_X1 U708 ( .A1(n630), .A2(n741), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n629), .A2(n726), .ZN(n633) );
  XOR2_X1 U710 ( .A(n630), .B(KEYINPUT86), .Z(n631) );
  NAND2_X1 U711 ( .A1(n631), .A2(KEYINPUT2), .ZN(n632) );
  INV_X1 U712 ( .A(n635), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT62), .B(KEYINPUT92), .Z(n636) );
  XOR2_X1 U714 ( .A(n638), .B(G101), .Z(n639) );
  XNOR2_X1 U715 ( .A(KEYINPUT114), .B(n639), .ZN(G3) );
  NOR2_X1 U716 ( .A1(n641), .A2(n654), .ZN(n640) );
  XOR2_X1 U717 ( .A(G104), .B(n640), .Z(G6) );
  NOR2_X1 U718 ( .A1(n657), .A2(n641), .ZN(n645) );
  XOR2_X1 U719 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n643) );
  XNOR2_X1 U720 ( .A(G107), .B(KEYINPUT115), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U722 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U723 ( .A(n646), .B(G110), .Z(G12) );
  XOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .Z(n649) );
  NAND2_X1 U725 ( .A1(n652), .A2(n647), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n649), .B(n648), .ZN(G30) );
  XNOR2_X1 U727 ( .A(G143), .B(n650), .ZN(G45) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(G146), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n654), .A2(n656), .ZN(n655) );
  XOR2_X1 U731 ( .A(G113), .B(n655), .Z(G15) );
  NOR2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U733 ( .A(G116), .B(n658), .Z(G18) );
  XNOR2_X1 U734 ( .A(n659), .B(G125), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n660), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U736 ( .A(G134), .B(n661), .Z(G36) );
  XOR2_X1 U737 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n663) );
  NOR2_X1 U738 ( .A1(n726), .A2(n663), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n706), .A2(n665), .ZN(n700) );
  NOR2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n673) );
  NOR2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n674), .A2(n695), .ZN(n689) );
  NAND2_X1 U745 ( .A1(n382), .A2(n675), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT50), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n348), .A2(n678), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n679), .B(KEYINPUT49), .ZN(n680) );
  NAND2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U752 ( .A(KEYINPUT51), .B(n686), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n687), .A2(n694), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  XOR2_X1 U756 ( .A(KEYINPUT116), .B(n691), .Z(n692) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n698) );
  NAND2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U759 ( .A(KEYINPUT117), .B(n696), .ZN(n697) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U762 ( .A(n702), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U763 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n705) );
  XNOR2_X1 U764 ( .A(n703), .B(KEYINPUT90), .ZN(n704) );
  XNOR2_X1 U765 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n710) );
  XNOR2_X1 U766 ( .A(n708), .B(KEYINPUT57), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n710), .B(n709), .ZN(n712) );
  XOR2_X1 U768 ( .A(n712), .B(n711), .Z(n713) );
  NOR2_X1 U769 ( .A1(n720), .A2(n713), .ZN(G54) );
  XNOR2_X1 U770 ( .A(n716), .B(KEYINPUT120), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n720), .A2(n719), .ZN(G66) );
  XNOR2_X1 U773 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n724) );
  NOR2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n734) );
  NAND2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n727), .B(KEYINPUT122), .ZN(n732) );
  XOR2_X1 U778 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n729) );
  NAND2_X1 U779 ( .A1(G224), .A2(G953), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U781 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U783 ( .A(n734), .B(n733), .Z(G69) );
  XOR2_X1 U784 ( .A(G227), .B(n740), .Z(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(G900), .ZN(n737) );
  XOR2_X1 U786 ( .A(KEYINPUT125), .B(n737), .Z(n738) );
  NAND2_X1 U787 ( .A1(G953), .A2(n738), .ZN(n739) );
  XNOR2_X1 U788 ( .A(n739), .B(KEYINPUT126), .ZN(n745) );
  XOR2_X1 U789 ( .A(n741), .B(n740), .Z(n743) );
  NAND2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n745), .A2(n744), .ZN(G72) );
  XNOR2_X1 U792 ( .A(G137), .B(n746), .ZN(n747) );
  XNOR2_X1 U793 ( .A(n747), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U794 ( .A(n748), .B(G122), .Z(G24) );
  XOR2_X1 U795 ( .A(G131), .B(n749), .Z(G33) );
  XNOR2_X1 U796 ( .A(G140), .B(n750), .ZN(G42) );
  XOR2_X1 U797 ( .A(n751), .B(G119), .Z(G21) );
endmodule

