//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  OR2_X1    g001(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(G141gat), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n212), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n208), .A2(new_n213), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT29), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G211gat), .A2(G218gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT71), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G197gat), .A2(G204gat), .ZN(new_n232));
  AND2_X1   g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(new_n229), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n227), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n235), .A2(new_n229), .ZN(new_n238));
  XNOR2_X1  g037(.A(G197gat), .B(G204gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n238), .A2(new_n226), .A3(new_n239), .A4(new_n231), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(G228gat), .B(G233gat), .C1(new_n225), .C2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G141gat), .B(G148gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n212), .B(new_n220), .C1(new_n243), .C2(KEYINPUT2), .ZN(new_n244));
  INV_X1    g043(.A(new_n207), .ZN(new_n245));
  AND2_X1   g044(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(new_n248), .B2(G141gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n213), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT29), .B1(new_n237), .B2(new_n240), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n242), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT81), .B(new_n251), .C1(new_n252), .C2(KEYINPUT3), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT82), .B1(new_n225), .B2(new_n241), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n244), .B(new_n224), .C1(new_n249), .C2(new_n250), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n241), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n257), .A2(new_n258), .A3(new_n259), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G228gat), .A2(G233gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n255), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT84), .ZN(new_n269));
  OAI21_X1  g068(.A(G22gat), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI211_X1 g069(.A(KEYINPUT84), .B(new_n255), .C1(new_n267), .C2(new_n266), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n202), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n267), .ZN(new_n273));
  INV_X1    g072(.A(new_n255), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT84), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n268), .A2(new_n269), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(KEYINPUT85), .A3(G22gat), .A4(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT83), .B(G22gat), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G78gat), .B(G106gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G50gat), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n272), .A2(new_n278), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n284), .B(KEYINPUT80), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n268), .A2(new_n279), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n280), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n286), .A2(KEYINPUT86), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT86), .B1(new_n286), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT0), .ZN(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G85gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n205), .A2(new_n207), .B1(new_n212), .B2(new_n211), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n221), .B1(new_n210), .B2(new_n216), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G113gat), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G127gat), .ZN(new_n309));
  INV_X1    g108(.A(G127gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G134gat), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n306), .A2(new_n307), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n311), .ZN(new_n313));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(KEYINPUT1), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n260), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n301), .A2(new_n260), .A3(KEYINPUT75), .A4(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n251), .B2(new_n316), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n312), .A2(new_n315), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n223), .A3(KEYINPUT4), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n322), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT5), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n223), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n251), .A2(new_n316), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n322), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n327), .B1(new_n319), .B2(new_n320), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(KEYINPUT5), .A3(new_n322), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n298), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT76), .B1(new_n340), .B2(KEYINPUT6), .ZN(new_n341));
  AND4_X1   g140(.A1(KEYINPUT5), .A2(new_n321), .A3(new_n322), .A4(new_n328), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n335), .B1(new_n338), .B2(new_n322), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n297), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n337), .A2(new_n298), .A3(new_n339), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT77), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n337), .A2(new_n350), .A3(new_n298), .A4(new_n339), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n341), .A2(new_n347), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n298), .A4(new_n339), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  NOR4_X1   g160(.A1(KEYINPUT67), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT67), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n361), .B2(new_n360), .ZN(new_n364));
  OAI221_X1 g163(.A(new_n359), .B1(new_n360), .B2(new_n361), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT27), .B(G183gat), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n368), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n370), .A3(new_n367), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n365), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G169gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT23), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  OAI221_X1 g175(.A(KEYINPUT25), .B1(G176gat), .B2(new_n374), .C1(new_n376), .C2(new_n361), .ZN(new_n377));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT24), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT24), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(G183gat), .A3(G190gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT66), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(KEYINPUT66), .A3(new_n383), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n377), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n361), .B1(KEYINPUT23), .B2(new_n359), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT65), .B(G176gat), .Z(new_n390));
  INV_X1    g189(.A(new_n374), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n383), .A2(KEYINPUT64), .ZN(new_n393));
  NOR2_X1   g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n382), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT25), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n372), .B1(new_n388), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT73), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n372), .B(new_n401), .C1(new_n388), .C2(new_n398), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n399), .B2(new_n261), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n403), .A2(new_n405), .B1(new_n406), .B2(KEYINPUT72), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT72), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n382), .A2(new_n393), .A3(new_n396), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT65), .B(G176gat), .ZN(new_n411));
  OAI22_X1  g210(.A1(new_n411), .A2(new_n374), .B1(new_n376), .B2(new_n361), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT25), .B1(new_n374), .B2(G176gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n389), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT66), .B1(new_n382), .B2(new_n383), .ZN(new_n416));
  AOI211_X1 g215(.A(new_n385), .B(new_n394), .C1(new_n379), .C2(new_n381), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT29), .B1(new_n419), .B2(new_n372), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n408), .B1(new_n420), .B2(new_n405), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n241), .B1(new_n407), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n405), .A2(KEYINPUT29), .ZN(new_n423));
  INV_X1    g222(.A(new_n402), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n401), .B1(new_n419), .B2(new_n372), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n419), .A2(new_n372), .A3(new_n405), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n263), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n358), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n405), .B1(new_n424), .B2(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n399), .A2(new_n261), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT72), .A3(new_n404), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n421), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n263), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n427), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n241), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n357), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n429), .A2(KEYINPUT30), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n428), .B1(new_n263), .B2(new_n433), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n357), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n293), .B1(new_n354), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n354), .A2(new_n293), .A3(new_n442), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n292), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n434), .B2(new_n436), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n448), .B2(new_n357), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT90), .B(new_n358), .C1(new_n439), .C2(new_n447), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n436), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT38), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n447), .B1(new_n435), .B2(new_n263), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n241), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n357), .A2(KEYINPUT38), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n452), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n460));
  AND4_X1   g259(.A1(new_n353), .A2(new_n459), .A3(new_n460), .A4(new_n437), .ZN(new_n461));
  INV_X1    g260(.A(new_n338), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n334), .ZN(new_n464));
  INV_X1    g263(.A(new_n333), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n465), .B2(new_n322), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n338), .B2(new_n322), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n467), .A3(new_n297), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n348), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n438), .A2(new_n472), .A3(new_n441), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n464), .A2(new_n467), .A3(new_n475), .A4(new_n297), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT88), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n474), .A2(new_n479), .A3(new_n469), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n454), .A2(new_n461), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n286), .A2(new_n289), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n286), .A2(KEYINPUT86), .A3(new_n289), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n489));
  XOR2_X1   g288(.A(G15gat), .B(G43gat), .Z(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n399), .A2(new_n316), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n419), .A2(new_n325), .A3(new_n372), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n492), .B1(new_n496), .B2(KEYINPUT33), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT32), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n494), .A2(new_n495), .ZN(new_n502));
  INV_X1    g301(.A(new_n493), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n501), .B(KEYINPUT34), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n497), .A2(new_n499), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n500), .A2(new_n504), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n504), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n497), .A2(new_n499), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n497), .A2(new_n499), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n513), .A3(KEYINPUT69), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT69), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n489), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n509), .A2(new_n513), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT70), .B1(new_n518), .B2(new_n489), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n520));
  AOI211_X1 g319(.A(new_n520), .B(KEYINPUT36), .C1(new_n509), .C2(new_n513), .ZN(new_n521));
  OR3_X1    g320(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n445), .A2(new_n488), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n444), .A2(new_n443), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n485), .A2(new_n486), .B1(new_n516), .B2(new_n514), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n518), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n460), .A2(new_n353), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n524), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n441), .B2(new_n438), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n528), .B(new_n531), .C1(new_n290), .C2(new_n291), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n523), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(G1gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n537), .B(new_n538), .C1(G1gat), .C2(new_n535), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G8gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n545));
  AOI21_X1  g344(.A(G36gat), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G36gat), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n542), .A2(new_n547), .A3(G29gat), .ZN(new_n548));
  OR3_X1    g347(.A1(new_n546), .A2(KEYINPUT15), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT15), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT17), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n552), .B2(new_n553), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n541), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n554), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n540), .B(new_n554), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n559), .B(KEYINPUT13), .Z(new_n564));
  AOI22_X1  g363(.A1(new_n561), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n558), .A2(KEYINPUT18), .A3(new_n559), .A4(new_n560), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G197gat), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT11), .B(G169gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT93), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n575), .B(new_n565), .C1(new_n568), .C2(new_n569), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n570), .A2(KEYINPUT93), .A3(new_n576), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT95), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(KEYINPUT9), .ZN(new_n589));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590));
  OAI22_X1  g389(.A1(new_n589), .A2(new_n590), .B1(KEYINPUT94), .B2(new_n588), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n587), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n598), .A2(new_n587), .A3(new_n599), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n584), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  INV_X1    g403(.A(new_n584), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n605), .A3(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G183gat), .B(G211gat), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n541), .B1(new_n594), .B2(new_n593), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n615), .A3(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT98), .ZN(new_n623));
  XOR2_X1   g422(.A(G134gat), .B(G162gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT101), .B(G92gat), .Z(new_n627));
  INV_X1    g426(.A(G85gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n629), .A2(KEYINPUT100), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT8), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n629), .B2(KEYINPUT100), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n627), .A2(new_n628), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT7), .ZN(new_n634));
  INV_X1    g433(.A(G92gat), .ZN(new_n635));
  OAI211_X1 g434(.A(KEYINPUT99), .B(new_n634), .C1(new_n628), .C2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT99), .B1(new_n628), .B2(new_n635), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(G85gat), .A3(G92gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n639), .A3(KEYINPUT7), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G99gat), .B(G106gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n633), .A2(new_n640), .A3(new_n642), .A4(new_n636), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(KEYINPUT102), .A3(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n649), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n648), .B(new_n647), .C1(new_n555), .C2(new_n557), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n650), .A2(new_n654), .A3(new_n651), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n626), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(KEYINPUT103), .B(new_n626), .C1(new_n655), .C2(new_n656), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n652), .A2(KEYINPUT104), .A3(new_n654), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT104), .B1(new_n652), .B2(new_n654), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n656), .A2(new_n626), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n659), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G230gat), .ZN(new_n666));
  INV_X1    g465(.A(G233gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n647), .A2(new_n593), .A3(new_n648), .ZN(new_n669));
  INV_X1    g468(.A(new_n593), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n644), .A3(new_n646), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n649), .A2(KEYINPUT10), .A3(new_n670), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n669), .A2(new_n671), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n668), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(G120gat), .B(G148gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT105), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n676), .A2(new_n678), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR4_X1   g486(.A1(new_n583), .A2(new_n620), .A3(new_n665), .A4(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n534), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n354), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  INV_X1    g491(.A(new_n442), .ZN(new_n693));
  OR2_X1    g492(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n689), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT106), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  INV_X1    g497(.A(new_n689), .ZN(new_n699));
  OAI21_X1  g498(.A(G8gat), .B1(new_n699), .B2(new_n442), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(G1325gat));
  OR3_X1    g501(.A1(new_n699), .A2(G15gat), .A3(new_n518), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n522), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT107), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n699), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n703), .A2(new_n709), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n689), .A2(new_n292), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NOR3_X1   g512(.A1(new_n583), .A2(new_n619), .A3(new_n687), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n534), .A2(new_n665), .A3(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n354), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n445), .A2(new_n488), .A3(new_n522), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n354), .A2(new_n442), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT78), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n514), .A2(new_n516), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n354), .A2(new_n293), .A3(new_n442), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n487), .A2(new_n722), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n533), .B1(new_n725), .B2(KEYINPUT35), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n719), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n523), .B(KEYINPUT109), .C1(new_n527), .C2(new_n533), .ZN(new_n728));
  INV_X1    g527(.A(new_n665), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT44), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n725), .A2(KEYINPUT35), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n722), .A2(new_n724), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n706), .B1(new_n733), .B2(new_n292), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n732), .A2(new_n532), .B1(new_n734), .B2(new_n488), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT44), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(KEYINPUT110), .A3(new_n714), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT110), .B1(new_n737), .B2(new_n714), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n739), .A2(new_n354), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n718), .B1(new_n741), .B2(new_n543), .ZN(G1328gat));
  NAND2_X1  g541(.A1(new_n693), .A2(new_n547), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n715), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT111), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(KEYINPUT112), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n739), .A2(new_n442), .A3(new_n740), .ZN(new_n749));
  OAI221_X1 g548(.A(new_n747), .B1(new_n745), .B2(new_n748), .C1(new_n749), .C2(new_n547), .ZN(G1329gat));
  NAND2_X1  g549(.A1(new_n737), .A2(new_n714), .ZN(new_n751));
  OAI21_X1  g550(.A(G43gat), .B1(new_n751), .B2(new_n522), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n715), .A2(G43gat), .A3(new_n518), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n708), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(new_n758), .A3(new_n738), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n753), .B1(new_n759), .B2(G43gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n760), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n715), .A2(KEYINPUT114), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n715), .A2(KEYINPUT114), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n487), .A2(G50gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G50gat), .B1(new_n751), .B2(new_n487), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n768), .B(new_n769), .C1(new_n767), .C2(new_n766), .ZN(new_n770));
  INV_X1    g569(.A(new_n766), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n757), .A2(new_n292), .A3(new_n738), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G50gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(G1331gat));
  INV_X1    g574(.A(new_n687), .ZN(new_n776));
  NOR4_X1   g575(.A1(new_n620), .A2(new_n582), .A3(new_n665), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n727), .A2(new_n728), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n354), .B(KEYINPUT116), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(G57gat), .Z(G1332gat));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n778), .A2(new_n782), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n693), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT49), .B(G64gat), .Z(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(G1333gat));
  INV_X1    g587(.A(G71gat), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n708), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n783), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n727), .A2(new_n728), .A3(new_n528), .A4(new_n777), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n789), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n783), .A2(new_n792), .A3(new_n784), .A4(new_n790), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(G1334gat));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n292), .A3(new_n784), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT119), .B(G78gat), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(G1335gat));
  NOR2_X1   g602(.A1(new_n735), .A2(new_n729), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n582), .A2(new_n619), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(KEYINPUT51), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n628), .A3(new_n690), .A4(new_n687), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n737), .A2(new_n687), .A3(new_n805), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n690), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n628), .ZN(G1336gat));
  NOR3_X1   g613(.A1(new_n442), .A2(new_n776), .A3(G92gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  AND4_X1   g615(.A1(new_n693), .A2(new_n737), .A3(new_n687), .A4(new_n805), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n627), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n816), .B(new_n820), .C1(new_n817), .C2(new_n627), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1337gat));
  XOR2_X1   g621(.A(KEYINPUT120), .B(G99gat), .Z(new_n823));
  NAND4_X1  g622(.A1(new_n810), .A2(new_n528), .A3(new_n687), .A4(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n812), .A2(new_n758), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(new_n823), .ZN(G1338gat));
  NOR2_X1   g625(.A1(new_n776), .A2(G106gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n292), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(G106gat), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n292), .A2(new_n737), .A3(new_n687), .A4(new_n805), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n828), .B(new_n833), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1339gat));
  NOR4_X1   g634(.A1(new_n620), .A2(new_n582), .A3(new_n665), .A4(new_n687), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n673), .A2(new_n674), .A3(new_n668), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n676), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n685), .B1(new_n675), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n843), .A2(new_n686), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n563), .A2(new_n564), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n574), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n579), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n665), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n687), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n582), .B2(new_n845), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n853), .B2(new_n665), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n836), .B1(new_n854), .B2(new_n620), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n779), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n526), .A2(new_n442), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n582), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n855), .A2(new_n292), .A3(new_n518), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n862), .A2(new_n690), .A3(new_n442), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n583), .A2(new_n304), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(G1340gat));
  AOI21_X1  g664(.A(G120gat), .B1(new_n860), .B2(new_n687), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n776), .A2(new_n302), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n863), .B2(new_n867), .ZN(G1341gat));
  NAND3_X1  g667(.A1(new_n863), .A2(G127gat), .A3(new_n619), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n871));
  AOI21_X1  g670(.A(G127gat), .B1(new_n860), .B2(new_n619), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1342gat));
  NOR3_X1   g672(.A1(new_n859), .A2(G134gat), .A3(new_n729), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n308), .B1(new_n863), .B2(new_n665), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(KEYINPUT56), .B2(new_n875), .ZN(G1343gat));
  OAI21_X1  g678(.A(KEYINPUT57), .B1(new_n855), .B2(new_n487), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n706), .A2(new_n354), .A3(new_n693), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n844), .A2(new_n686), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n580), .A2(new_n882), .A3(new_n581), .A4(new_n843), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n665), .B1(new_n883), .B2(new_n851), .ZN(new_n884));
  INV_X1    g683(.A(new_n850), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n620), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n583), .A2(new_n619), .A3(new_n729), .A4(new_n776), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n292), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n880), .A2(new_n881), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(G141gat), .A3(new_n582), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n758), .A2(new_n487), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n856), .A2(new_n893), .A3(new_n442), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n206), .B1(new_n894), .B2(new_n583), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g696(.A(new_n894), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n248), .A3(new_n687), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n292), .A2(new_n901), .A3(new_n889), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n890), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n902), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n687), .A3(new_n881), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n900), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n248), .C1(new_n891), .C2(new_n687), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(G1345gat));
  NOR3_X1   g708(.A1(new_n894), .A2(KEYINPUT123), .A3(new_n620), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(G155gat), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT123), .B1(new_n894), .B2(new_n620), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n620), .A2(new_n218), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n911), .A2(new_n912), .B1(new_n891), .B2(new_n913), .ZN(G1346gat));
  AOI21_X1  g713(.A(G162gat), .B1(new_n898), .B2(new_n665), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n729), .A2(new_n219), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n891), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n855), .A2(new_n690), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n693), .A3(new_n526), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n582), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n779), .A2(new_n693), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n862), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n373), .A3(new_n583), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT124), .Z(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n920), .B2(new_n687), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n923), .A2(new_n390), .A3(new_n776), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  NAND3_X1  g728(.A1(new_n920), .A2(new_n366), .A3(new_n619), .ZN(new_n930));
  OAI21_X1  g729(.A(G183gat), .B1(new_n923), .B2(new_n620), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n923), .B2(new_n729), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT61), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n367), .A3(new_n665), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1351gat));
  AOI21_X1  g736(.A(new_n889), .B1(new_n888), .B2(new_n292), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT57), .B(new_n487), .C1(new_n886), .C2(new_n887), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n902), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n903), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT125), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n940), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n708), .A2(new_n922), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n943), .A2(new_n582), .A3(new_n945), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT126), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n905), .B2(new_n944), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n950), .A2(new_n951), .A3(new_n582), .A4(new_n943), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n952), .A3(G197gat), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n918), .A2(new_n693), .A3(new_n893), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n955), .A2(G197gat), .A3(new_n583), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n953), .A2(new_n956), .ZN(G1352gat));
  NOR3_X1   g756(.A1(new_n955), .A2(G204gat), .A3(new_n776), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n950), .A2(new_n687), .A3(new_n943), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G204gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1353gat));
  OR3_X1    g761(.A1(new_n955), .A2(G211gat), .A3(new_n620), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n620), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n940), .A2(new_n941), .A3(new_n964), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n963), .B(KEYINPUT127), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1354gat));
  AND4_X1   g771(.A1(G218gat), .A2(new_n950), .A3(new_n665), .A4(new_n943), .ZN(new_n973));
  AOI21_X1  g772(.A(G218gat), .B1(new_n954), .B2(new_n665), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(G1355gat));
endmodule


