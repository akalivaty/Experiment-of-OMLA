

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585;

  INV_X1 U319 ( .A(n491), .ZN(n557) );
  INV_X1 U320 ( .A(n476), .ZN(n484) );
  XNOR2_X1 U321 ( .A(n450), .B(KEYINPUT38), .ZN(n510) );
  NOR2_X1 U322 ( .A1(n485), .A2(n496), .ZN(n450) );
  XNOR2_X1 U323 ( .A(n411), .B(n410), .ZN(n485) );
  OR2_X1 U324 ( .A1(n409), .A2(n495), .ZN(n411) );
  NOR2_X1 U325 ( .A1(n471), .A2(n528), .ZN(n472) );
  XOR2_X2 U326 ( .A(KEYINPUT94), .B(n403), .Z(n528) );
  XNOR2_X1 U327 ( .A(n380), .B(KEYINPUT95), .ZN(n381) );
  NOR2_X1 U328 ( .A1(n535), .A2(n392), .ZN(n393) );
  NOR2_X1 U329 ( .A1(n401), .A2(n400), .ZN(n402) );
  AND2_X1 U330 ( .A1(n528), .A2(n391), .ZN(n549) );
  XNOR2_X1 U331 ( .A(n469), .B(KEYINPUT48), .ZN(n548) );
  XNOR2_X1 U332 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U333 ( .A(KEYINPUT89), .B(n430), .Z(n287) );
  XNOR2_X1 U334 ( .A(n455), .B(KEYINPUT113), .ZN(n456) );
  XNOR2_X1 U335 ( .A(n457), .B(n456), .ZN(n459) );
  XNOR2_X1 U336 ( .A(n353), .B(G50GAT), .ZN(n354) );
  XNOR2_X1 U337 ( .A(n405), .B(KEYINPUT100), .ZN(n406) );
  XNOR2_X1 U338 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U339 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U340 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U341 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U342 ( .A(n437), .B(n384), .ZN(n385) );
  XOR2_X1 U343 ( .A(n361), .B(n387), .Z(n471) );
  XNOR2_X1 U344 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U345 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U346 ( .A(n451), .B(G43GAT), .ZN(n452) );
  XNOR2_X1 U347 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G78GAT), .B(G211GAT), .Z(n289) );
  XNOR2_X1 U350 ( .A(G127GAT), .B(G183GAT), .ZN(n288) );
  XNOR2_X1 U351 ( .A(n289), .B(n288), .ZN(n290) );
  XOR2_X1 U352 ( .A(G71GAT), .B(KEYINPUT13), .Z(n439) );
  XOR2_X1 U353 ( .A(n290), .B(n439), .Z(n292) );
  XNOR2_X1 U354 ( .A(G155GAT), .B(G57GAT), .ZN(n291) );
  XNOR2_X1 U355 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U356 ( .A(KEYINPUT67), .B(G22GAT), .Z(n294) );
  XNOR2_X1 U357 ( .A(G1GAT), .B(G15GAT), .ZN(n293) );
  XNOR2_X1 U358 ( .A(n294), .B(n293), .ZN(n412) );
  XOR2_X1 U359 ( .A(n412), .B(KEYINPUT12), .Z(n296) );
  NAND2_X1 U360 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U361 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U362 ( .A(n298), .B(n297), .Z(n306) );
  XOR2_X1 U363 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n300) );
  XNOR2_X1 U364 ( .A(G64GAT), .B(G8GAT), .ZN(n299) );
  XNOR2_X1 U365 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U366 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n302) );
  XNOR2_X1 U367 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n301) );
  XNOR2_X1 U368 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U369 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U370 ( .A(n306), .B(n305), .Z(n564) );
  XOR2_X1 U371 ( .A(KEYINPUT9), .B(G106GAT), .Z(n308) );
  NAND2_X1 U372 ( .A1(G232GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U373 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U374 ( .A(n309), .B(KEYINPUT10), .ZN(n317) );
  XOR2_X1 U375 ( .A(KEYINPUT70), .B(G99GAT), .Z(n311) );
  XNOR2_X1 U376 ( .A(KEYINPUT71), .B(G92GAT), .ZN(n310) );
  XNOR2_X1 U377 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U378 ( .A(G85GAT), .B(n312), .ZN(n447) );
  XOR2_X1 U379 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n314) );
  XNOR2_X1 U380 ( .A(G162GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U381 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U382 ( .A(n447), .B(n315), .ZN(n316) );
  XNOR2_X1 U383 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U384 ( .A(G190GAT), .B(G36GAT), .Z(n388) );
  XNOR2_X1 U385 ( .A(n318), .B(n388), .ZN(n322) );
  XOR2_X1 U386 ( .A(G29GAT), .B(G134GAT), .Z(n365) );
  XOR2_X1 U387 ( .A(G43GAT), .B(G50GAT), .Z(n320) );
  XNOR2_X1 U388 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n319) );
  XNOR2_X1 U389 ( .A(n320), .B(n319), .ZN(n418) );
  XNOR2_X1 U390 ( .A(n365), .B(n418), .ZN(n321) );
  XNOR2_X1 U391 ( .A(n322), .B(n321), .ZN(n491) );
  XNOR2_X1 U392 ( .A(KEYINPUT36), .B(n557), .ZN(n581) );
  NAND2_X1 U393 ( .A1(n564), .A2(n581), .ZN(n409) );
  XOR2_X1 U394 ( .A(KEYINPUT83), .B(G169GAT), .Z(n324) );
  XNOR2_X1 U395 ( .A(G120GAT), .B(KEYINPUT82), .ZN(n323) );
  XNOR2_X1 U396 ( .A(n324), .B(n323), .ZN(n333) );
  XOR2_X1 U397 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n326) );
  XNOR2_X1 U398 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n325) );
  XNOR2_X1 U399 ( .A(n326), .B(n325), .ZN(n382) );
  XOR2_X1 U400 ( .A(KEYINPUT20), .B(n382), .Z(n331) );
  XOR2_X1 U401 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n328) );
  XNOR2_X1 U402 ( .A(G127GAT), .B(G113GAT), .ZN(n327) );
  XNOR2_X1 U403 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U404 ( .A(KEYINPUT80), .B(n329), .Z(n376) );
  XNOR2_X1 U405 ( .A(n376), .B(G15GAT), .ZN(n330) );
  XNOR2_X1 U406 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U407 ( .A(n333), .B(n332), .ZN(n341) );
  NAND2_X1 U408 ( .A1(G227GAT), .A2(G233GAT), .ZN(n339) );
  XOR2_X1 U409 ( .A(G176GAT), .B(G71GAT), .Z(n335) );
  XNOR2_X1 U410 ( .A(G43GAT), .B(G190GAT), .ZN(n334) );
  XNOR2_X1 U411 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U412 ( .A(G134GAT), .B(G99GAT), .Z(n336) );
  XNOR2_X1 U413 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U414 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U415 ( .A(n341), .B(n340), .Z(n522) );
  INV_X1 U416 ( .A(n522), .ZN(n535) );
  XOR2_X1 U417 ( .A(KEYINPUT2), .B(G162GAT), .Z(n343) );
  XNOR2_X1 U418 ( .A(G155GAT), .B(G141GAT), .ZN(n342) );
  XNOR2_X1 U419 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U420 ( .A(KEYINPUT3), .B(n344), .Z(n377) );
  XNOR2_X1 U421 ( .A(G106GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U422 ( .A(n345), .B(G204GAT), .ZN(n430) );
  NAND2_X1 U423 ( .A1(G228GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U424 ( .A(n287), .B(n346), .ZN(n355) );
  XOR2_X1 U425 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n348) );
  XNOR2_X1 U426 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n347) );
  XNOR2_X1 U427 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U428 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n350) );
  XNOR2_X1 U429 ( .A(G148GAT), .B(G22GAT), .ZN(n349) );
  XNOR2_X1 U430 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U431 ( .A(n352), .B(n351), .Z(n353) );
  XNOR2_X1 U432 ( .A(n377), .B(n356), .ZN(n361) );
  XNOR2_X1 U433 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n357) );
  XNOR2_X1 U434 ( .A(n357), .B(KEYINPUT88), .ZN(n358) );
  XOR2_X1 U435 ( .A(n358), .B(KEYINPUT21), .Z(n360) );
  XNOR2_X1 U436 ( .A(G218GAT), .B(G211GAT), .ZN(n359) );
  XOR2_X1 U437 ( .A(n360), .B(n359), .Z(n387) );
  XOR2_X1 U438 ( .A(KEYINPUT28), .B(n471), .Z(n525) );
  XNOR2_X1 U439 ( .A(G120GAT), .B(G148GAT), .ZN(n362) );
  XNOR2_X1 U440 ( .A(n362), .B(G57GAT), .ZN(n440) );
  XOR2_X1 U441 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n364) );
  XNOR2_X1 U442 ( .A(G85GAT), .B(G1GAT), .ZN(n363) );
  XNOR2_X1 U443 ( .A(n364), .B(n363), .ZN(n366) );
  XNOR2_X1 U444 ( .A(n366), .B(n365), .ZN(n368) );
  AND2_X1 U445 ( .A1(G225GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U446 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U447 ( .A(n440), .B(n369), .Z(n371) );
  XNOR2_X1 U448 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n370) );
  XNOR2_X1 U449 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U450 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n373) );
  XNOR2_X1 U451 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n372) );
  XNOR2_X1 U452 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U453 ( .A(n375), .B(n374), .Z(n379) );
  XNOR2_X1 U454 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U455 ( .A(n379), .B(n378), .ZN(n403) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n380) );
  XOR2_X1 U457 ( .A(G8GAT), .B(G169GAT), .Z(n413) );
  XNOR2_X1 U458 ( .A(n383), .B(n413), .ZN(n386) );
  XOR2_X1 U459 ( .A(G64GAT), .B(G176GAT), .Z(n437) );
  XOR2_X1 U460 ( .A(G92GAT), .B(G204GAT), .Z(n384) );
  XOR2_X1 U461 ( .A(n388), .B(n387), .Z(n389) );
  XOR2_X1 U462 ( .A(n390), .B(n389), .Z(n520) );
  XNOR2_X1 U463 ( .A(n520), .B(KEYINPUT27), .ZN(n399) );
  INV_X1 U464 ( .A(n399), .ZN(n391) );
  NAND2_X1 U465 ( .A1(n525), .A2(n549), .ZN(n537) );
  XNOR2_X1 U466 ( .A(KEYINPUT96), .B(n537), .ZN(n392) );
  XNOR2_X1 U467 ( .A(n393), .B(KEYINPUT97), .ZN(n407) );
  OR2_X1 U468 ( .A1(n520), .A2(n522), .ZN(n394) );
  XNOR2_X1 U469 ( .A(n394), .B(KEYINPUT98), .ZN(n396) );
  INV_X1 U470 ( .A(n471), .ZN(n395) );
  NAND2_X1 U471 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U472 ( .A(KEYINPUT25), .B(n397), .ZN(n401) );
  NAND2_X1 U473 ( .A1(n471), .A2(n522), .ZN(n398) );
  XNOR2_X1 U474 ( .A(n398), .B(KEYINPUT26), .ZN(n568) );
  NOR2_X1 U475 ( .A1(n399), .A2(n568), .ZN(n400) );
  XNOR2_X1 U476 ( .A(KEYINPUT99), .B(n402), .ZN(n404) );
  NAND2_X1 U477 ( .A1(n404), .A2(n403), .ZN(n405) );
  NAND2_X1 U478 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n408), .B(KEYINPUT101), .ZN(n495) );
  XOR2_X1 U480 ( .A(KEYINPUT104), .B(KEYINPUT37), .Z(n410) );
  XOR2_X1 U481 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n417) );
  INV_X1 U484 ( .A(KEYINPUT66), .ZN(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n418), .B(KEYINPUT68), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n428) );
  XOR2_X1 U488 ( .A(G197GAT), .B(G36GAT), .Z(n422) );
  XNOR2_X1 U489 ( .A(G29GAT), .B(G113GAT), .ZN(n421) );
  XNOR2_X1 U490 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U491 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n424) );
  XNOR2_X1 U492 ( .A(G141GAT), .B(KEYINPUT29), .ZN(n423) );
  XNOR2_X1 U493 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U494 ( .A(n426), .B(n425), .Z(n427) );
  XOR2_X1 U495 ( .A(n428), .B(n427), .Z(n571) );
  INV_X1 U496 ( .A(n571), .ZN(n561) );
  INV_X1 U497 ( .A(KEYINPUT33), .ZN(n429) );
  XNOR2_X1 U498 ( .A(n430), .B(n429), .ZN(n434) );
  INV_X1 U499 ( .A(n434), .ZN(n432) );
  NAND2_X1 U500 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  INV_X1 U501 ( .A(n433), .ZN(n431) );
  NAND2_X1 U502 ( .A1(n432), .A2(n431), .ZN(n436) );
  NAND2_X1 U503 ( .A1(n434), .A2(n433), .ZN(n435) );
  NAND2_X1 U504 ( .A1(n436), .A2(n435), .ZN(n438) );
  XNOR2_X1 U505 ( .A(n438), .B(n437), .ZN(n446) );
  XOR2_X1 U506 ( .A(n440), .B(n439), .Z(n444) );
  XOR2_X1 U507 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n442) );
  XNOR2_X1 U508 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n441) );
  XNOR2_X1 U509 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n454) );
  NOR2_X1 U511 ( .A1(n561), .A2(n454), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n449), .B(KEYINPUT73), .ZN(n496) );
  NAND2_X1 U513 ( .A1(n510), .A2(n535), .ZN(n453) );
  XOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n451) );
  XNOR2_X1 U515 ( .A(KEYINPUT41), .B(n454), .ZN(n476) );
  INV_X1 U516 ( .A(n520), .ZN(n530) );
  NAND2_X1 U517 ( .A1(n571), .A2(n484), .ZN(n457) );
  XOR2_X1 U518 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n455) );
  INV_X1 U519 ( .A(n564), .ZN(n579) );
  NOR2_X1 U520 ( .A1(n557), .A2(n579), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n460), .B(KEYINPUT115), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n461), .B(KEYINPUT47), .ZN(n468) );
  XOR2_X1 U524 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n463) );
  NAND2_X1 U525 ( .A1(n579), .A2(n581), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n464) );
  NAND2_X1 U527 ( .A1(n464), .A2(n561), .ZN(n465) );
  NOR2_X1 U528 ( .A1(n454), .A2(n465), .ZN(n466) );
  XOR2_X1 U529 ( .A(KEYINPUT116), .B(n466), .Z(n467) );
  NAND2_X1 U530 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n530), .A2(n548), .ZN(n470) );
  XOR2_X1 U532 ( .A(KEYINPUT54), .B(n470), .Z(n567) );
  AND2_X1 U533 ( .A1(n567), .A2(n472), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT55), .ZN(n474) );
  NOR2_X1 U535 ( .A1(n522), .A2(n474), .ZN(n475) );
  XNOR2_X1 U536 ( .A(KEYINPUT121), .B(n475), .ZN(n563) );
  NOR2_X1 U537 ( .A1(n476), .A2(n563), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n477), .B(G176GAT), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  NOR2_X1 U541 ( .A1(n491), .A2(n563), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n481) );
  XNOR2_X1 U543 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n480) );
  NAND2_X1 U544 ( .A1(n561), .A2(n484), .ZN(n514) );
  NOR2_X1 U545 ( .A1(n514), .A2(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT110), .ZN(n533) );
  INV_X1 U547 ( .A(n525), .ZN(n509) );
  NAND2_X1 U548 ( .A1(n533), .A2(n509), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n488) );
  INV_X1 U550 ( .A(G106GAT), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1339GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n498) );
  XOR2_X1 U553 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n493) );
  NAND2_X1 U554 ( .A1(n579), .A2(n491), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  OR2_X1 U556 ( .A1(n495), .A2(n494), .ZN(n513) );
  NOR2_X1 U557 ( .A1(n496), .A2(n513), .ZN(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n528), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U560 ( .A(G1GAT), .B(n499), .Z(G1324GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n530), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n502) );
  NAND2_X1 U564 ( .A1(n504), .A2(n535), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U566 ( .A(G15GAT), .B(n503), .Z(G1326GAT) );
  NAND2_X1 U567 ( .A1(n509), .A2(n504), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT39), .Z(n507) );
  NAND2_X1 U570 ( .A1(n528), .A2(n510), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NAND2_X1 U572 ( .A1(n510), .A2(n530), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U574 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT106), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(n512), .ZN(G1331GAT) );
  NOR2_X1 U577 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(n515), .Z(n524) );
  INV_X1 U579 ( .A(n528), .ZN(n566) );
  NOR2_X1 U580 ( .A1(n524), .A2(n566), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n519) );
  XOR2_X1 U583 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1332GAT) );
  NOR2_X1 U585 ( .A1(n524), .A2(n520), .ZN(n521) );
  XOR2_X1 U586 ( .A(G64GAT), .B(n521), .Z(G1333GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n524), .ZN(n523) );
  XOR2_X1 U588 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n533), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n529), .ZN(G1336GAT) );
  XOR2_X1 U594 ( .A(G92GAT), .B(KEYINPUT111), .Z(n532) );
  NAND2_X1 U595 ( .A1(n530), .A2(n533), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n535), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U600 ( .A1(n548), .A2(n535), .ZN(n536) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n544), .A2(n571), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U605 ( .A1(n544), .A2(n484), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n544), .A2(n579), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U611 ( .A1(n544), .A2(n557), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U615 ( .A1(n568), .A2(n550), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n558), .A2(n571), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n553) );
  NAND2_X1 U619 ( .A1(n558), .A2(n484), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .Z(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n579), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT120), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n563), .ZN(n562) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n562), .Z(G1348GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  XOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .Z(n573) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT124), .ZN(n582) );
  NAND2_X1 U636 ( .A1(n571), .A2(n582), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n582), .A2(n454), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

