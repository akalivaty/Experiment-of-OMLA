//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT85), .ZN(new_n204));
  OR3_X1    g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT88), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT87), .B(G29gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G36gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n213), .B1(new_n212), .B2(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n205), .B(KEYINPUT86), .ZN(new_n216));
  INV_X1    g015(.A(new_n204), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n209), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT15), .A3(new_n210), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G1gat), .B2(new_n222), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(G8gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT89), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n215), .A2(new_n219), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n221), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n226), .A2(new_n232), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n228), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n202), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n236), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT91), .B1(new_n235), .B2(new_n228), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n228), .B2(new_n235), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n238), .B(KEYINPUT13), .Z(new_n244));
  INV_X1    g043(.A(new_n235), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(KEYINPUT91), .A3(new_n220), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n240), .A2(new_n241), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT84), .ZN(new_n250));
  XOR2_X1   g049(.A(G113gat), .B(G141gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G169gat), .B(G197gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT12), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n240), .A2(new_n247), .A3(new_n255), .A4(new_n241), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(KEYINPUT92), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT92), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n248), .A2(new_n260), .A3(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT93), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(KEYINPUT93), .A3(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT27), .B(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT28), .ZN(new_n271));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n272), .A2(KEYINPUT26), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  INV_X1    g080(.A(G183gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n269), .A2(G183gat), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(G183gat), .A3(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n280), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G183gat), .B(G190gat), .ZN(new_n289));
  OAI211_X1 g088(.A(KEYINPUT65), .B(new_n286), .C1(new_n289), .C2(new_n281), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n272), .A2(KEYINPUT23), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n275), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n288), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n286), .B1(new_n289), .B2(new_n281), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n291), .A2(new_n293), .A3(KEYINPUT25), .A4(new_n275), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT66), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n304));
  AOI211_X1 g103(.A(new_n304), .B(new_n301), .C1(new_n296), .C2(new_n297), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n279), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  NAND2_X1  g109(.A1(G113gat), .A2(G120gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G134gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G127gat), .ZN(new_n314));
  INV_X1    g113(.A(G127gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G134gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n311), .ZN(new_n319));
  NOR2_X1   g118(.A1(G113gat), .A2(G120gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT68), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT68), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n309), .A2(new_n322), .A3(new_n311), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n323), .A3(new_n310), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G127gat), .B(G134gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n318), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G227gat), .ZN(new_n331));
  INV_X1    g130(.A(G233gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n324), .A2(new_n328), .ZN(new_n334));
  INV_X1    g133(.A(new_n318), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(new_n279), .C1(new_n303), .C2(new_n305), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n330), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n339));
  XNOR2_X1  g138(.A(G15gat), .B(G43gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n338), .B(KEYINPUT32), .C1(new_n339), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n342), .B1(new_n338), .B2(KEYINPUT32), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(new_n339), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n344), .A2(KEYINPUT70), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT70), .B1(new_n344), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n337), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT34), .ZN(new_n350));
  INV_X1    g149(.A(new_n333), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT71), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n333), .B1(new_n330), .B2(new_n337), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n355), .A2(new_n350), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT71), .A3(new_n350), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n358), .B(new_n343), .C1(new_n347), .C2(new_n346), .ZN(new_n361));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365));
  INV_X1    g164(.A(G211gat), .ZN(new_n366));
  INV_X1    g165(.A(G218gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G211gat), .B(G218gat), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n363), .B1(new_n372), .B2(KEYINPUT29), .ZN(new_n373));
  NAND2_X1  g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374));
  INV_X1    g173(.A(G155gat), .ZN(new_n375));
  INV_X1    g174(.A(G162gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G141gat), .B(G148gat), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n374), .B(new_n377), .C1(new_n378), .C2(KEYINPUT2), .ZN(new_n379));
  INV_X1    g178(.A(G141gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G148gat), .ZN(new_n381));
  INV_X1    g180(.A(G148gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G141gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n377), .A2(new_n374), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(KEYINPUT2), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n362), .B1(new_n373), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n379), .A2(new_n363), .A3(new_n387), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n371), .B1(new_n392), .B2(KEYINPUT75), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(KEYINPUT75), .B2(new_n392), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n379), .A2(new_n387), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n370), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n391), .B(new_n397), .C1(new_n371), .C2(KEYINPUT74), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n398), .B2(new_n363), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n371), .B1(new_n391), .B2(new_n390), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n362), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(KEYINPUT76), .A2(G22gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(KEYINPUT76), .A2(G22gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G78gat), .B(G106gat), .Z(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n406), .B(new_n409), .C1(new_n403), .C2(new_n404), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n402), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n402), .B2(new_n412), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n360), .A2(new_n361), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT35), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n336), .A2(new_n419), .A3(new_n390), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n329), .B2(new_n396), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n329), .A2(new_n396), .A3(new_n421), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT72), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n336), .A2(new_n388), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n329), .A2(new_n396), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n425), .A2(new_n428), .B1(new_n431), .B2(KEYINPUT5), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n433), .B(new_n427), .C1(new_n423), .C2(new_n424), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n418), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n436));
  INV_X1    g235(.A(new_n424), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n420), .B2(new_n422), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n438), .B2(new_n427), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n425), .A2(KEYINPUT5), .A3(new_n428), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT79), .A3(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G1gat), .B(G29gat), .Z(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT73), .B(KEYINPUT0), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n435), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n440), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT6), .B1(new_n449), .B2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n447), .A4(new_n440), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G8gat), .B(G36gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n301), .B1(new_n296), .B2(new_n297), .ZN(new_n458));
  INV_X1    g257(.A(G226gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n332), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n458), .A2(new_n278), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n460), .A2(KEYINPUT29), .ZN(new_n463));
  AOI211_X1 g262(.A(new_n371), .B(new_n462), .C1(new_n306), .C2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n279), .B(new_n460), .C1(new_n303), .C2(new_n305), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n458), .B2(new_n278), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n372), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n457), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n462), .ZN(new_n469));
  INV_X1    g268(.A(new_n297), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n294), .B1(new_n299), .B2(new_n280), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(new_n290), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n304), .B1(new_n472), .B2(new_n301), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n278), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n463), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n469), .B(new_n372), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n465), .A2(new_n466), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n477), .B(new_n456), .C1(new_n478), .C2(new_n372), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n467), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n477), .A4(new_n456), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n453), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT80), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n453), .A2(new_n484), .A3(KEYINPUT80), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n417), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n416), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n417), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n453), .A2(new_n484), .A3(KEYINPUT80), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT80), .B1(new_n453), .B2(new_n484), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n360), .A2(new_n361), .A3(new_n415), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT82), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n439), .A2(new_n447), .A3(new_n440), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n450), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n452), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT35), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n491), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n348), .A2(new_n359), .ZN(new_n504));
  INV_X1    g303(.A(new_n361), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n415), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT39), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n429), .A2(new_n430), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n428), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n428), .B2(new_n425), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n438), .A2(new_n427), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n513), .B(new_n446), .C1(KEYINPUT39), .C2(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(KEYINPUT78), .A2(KEYINPUT40), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n517), .A2(new_n448), .ZN(new_n518));
  INV_X1    g317(.A(new_n484), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n509), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n468), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n456), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n481), .B2(new_n477), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT38), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n451), .A2(new_n452), .A3(new_n479), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n469), .B(new_n371), .C1(new_n475), .C2(new_n476), .ZN(new_n528));
  OAI211_X1 g327(.A(KEYINPUT37), .B(new_n528), .C1(new_n478), .C2(new_n371), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT38), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n526), .B(new_n527), .C1(new_n524), .C2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n520), .A2(new_n532), .B1(new_n501), .B2(new_n509), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n507), .B1(new_n360), .B2(new_n361), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n267), .B1(new_n503), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G71gat), .B(G78gat), .Z(new_n541));
  OR2_X1    g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT21), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n245), .B1(new_n545), .B2(new_n544), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT20), .ZN(new_n554));
  XOR2_X1   g353(.A(G127gat), .B(G155gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G183gat), .B(G211gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT96), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n552), .A2(new_n559), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  OAI21_X1  g363(.A(G92gat), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G92gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n565), .A2(new_n567), .B1(new_n563), .B2(new_n564), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n571), .B2(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  NAND3_X1  g375(.A1(new_n221), .A2(new_n230), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n574), .B(new_n575), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n228), .A2(new_n578), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT99), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n581), .B(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT97), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n584), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT100), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT102), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n543), .A3(new_n542), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT10), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n544), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n595), .A3(new_n594), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n593), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n594), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(new_n592), .ZN(new_n601));
  XOR2_X1   g400(.A(G120gat), .B(G148gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT101), .ZN(new_n603));
  XOR2_X1   g402(.A(G176gat), .B(G204gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n596), .A2(new_n598), .ZN(new_n607));
  INV_X1    g406(.A(new_n592), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n600), .A2(new_n592), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n605), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n562), .A2(new_n590), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n537), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n500), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G1gat), .ZN(G1324gat));
  INV_X1    g416(.A(new_n614), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G8gat), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n618), .A2(new_n484), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G8gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n614), .B2(new_n519), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT42), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(KEYINPUT42), .B2(new_n621), .ZN(G1325gat));
  NAND3_X1  g424(.A1(new_n508), .A2(KEYINPUT104), .A3(new_n535), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT36), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(new_n534), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(G15gat), .B1(new_n618), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n506), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n633), .A2(G15gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n618), .B2(new_n634), .ZN(G1326gat));
  NAND2_X1  g434(.A1(new_n614), .A2(new_n509), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT43), .B(G22gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  INV_X1    g437(.A(new_n612), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n562), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n590), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n537), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n643), .A2(new_n500), .A3(new_n208), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT45), .Z(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n503), .A2(new_n536), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(new_n590), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT105), .ZN(new_n650));
  AOI211_X1 g449(.A(new_n641), .B(new_n650), .C1(new_n503), .C2(new_n536), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n640), .A2(new_n262), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n208), .B1(new_n654), .B2(new_n500), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n645), .A2(new_n655), .ZN(G1328gat));
  OAI21_X1  g455(.A(G36gat), .B1(new_n654), .B2(new_n484), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n643), .A2(G36gat), .A3(new_n484), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT46), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(G1329gat));
  NOR2_X1   g459(.A1(new_n628), .A2(new_n534), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n652), .A2(new_n662), .A3(new_n653), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G43gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n633), .A2(G43gat), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n537), .A2(new_n642), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(KEYINPUT47), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n630), .B(new_n653), .C1(new_n648), .C2(new_n651), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n668), .A2(new_n667), .B1(new_n671), .B2(G43gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(KEYINPUT47), .B2(new_n672), .ZN(G1330gat));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674));
  INV_X1    g473(.A(G50gat), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n415), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n653), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n643), .B2(new_n415), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n674), .B(KEYINPUT48), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n674), .A2(KEYINPUT48), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(KEYINPUT48), .ZN(new_n681));
  AND4_X1   g480(.A1(new_n680), .A2(new_n677), .A3(new_n681), .A4(new_n678), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n679), .A2(new_n682), .ZN(G1331gat));
  INV_X1    g482(.A(new_n262), .ZN(new_n684));
  NOR4_X1   g483(.A1(new_n684), .A2(new_n562), .A3(new_n590), .A4(new_n639), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n647), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n615), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g488(.A(new_n484), .B(KEYINPUT108), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  AND2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n692), .B2(new_n693), .ZN(G1333gat));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697));
  INV_X1    g496(.A(G71gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n631), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n699), .B2(new_n687), .ZN(new_n700));
  NOR4_X1   g499(.A1(new_n686), .A2(new_n631), .A3(KEYINPUT109), .A4(new_n698), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT110), .B1(new_n686), .B2(new_n633), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n698), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n686), .A2(KEYINPUT110), .A3(new_n633), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n700), .A2(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT50), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n707));
  OAI221_X1 g506(.A(new_n707), .B1(new_n703), .B2(new_n704), .C1(new_n700), .C2(new_n701), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1334gat));
  NOR2_X1   g508(.A1(new_n686), .A2(new_n415), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT111), .B(G78gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1335gat));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n647), .A2(KEYINPUT113), .A3(new_n590), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n262), .A2(new_n562), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n641), .B1(new_n503), .B2(new_n536), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(KEYINPUT113), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n713), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n718), .A2(KEYINPUT113), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n715), .B1(new_n718), .B2(KEYINPUT113), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT51), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n615), .A2(new_n612), .A3(new_n564), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT114), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n715), .A2(new_n639), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT112), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n615), .B(new_n729), .C1(new_n648), .C2(new_n651), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G85gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(KEYINPUT115), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT115), .ZN(new_n733));
  INV_X1    g532(.A(new_n726), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n720), .B2(new_n723), .ZN(new_n735));
  INV_X1    g534(.A(new_n731), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(G1336gat));
  NOR3_X1   g537(.A1(new_n691), .A2(G92gat), .A3(new_n639), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n690), .B(new_n729), .C1(new_n648), .C2(new_n651), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n566), .A2(KEYINPUT52), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(KEYINPUT52), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n519), .B(new_n729), .C1(new_n648), .C2(new_n651), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(G92gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n739), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n720), .B2(new_n723), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(new_n743), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n750), .B2(new_n751), .ZN(G1337gat));
  XOR2_X1   g551(.A(KEYINPUT117), .B(G99gat), .Z(new_n753));
  NOR2_X1   g552(.A1(new_n639), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n724), .A2(new_n506), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n652), .A2(new_n630), .A3(new_n729), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1338gat));
  NOR3_X1   g557(.A1(new_n639), .A2(G106gat), .A3(new_n415), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n724), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n509), .B(new_n729), .C1(new_n648), .C2(new_n651), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n759), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n720), .B2(new_n723), .ZN(new_n766));
  INV_X1    g565(.A(new_n763), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT53), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(G1339gat));
  NOR2_X1   g568(.A1(new_n262), .A2(G113gat), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n593), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n609), .B(KEYINPUT54), .C1(new_n607), .C2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n605), .B1(new_n599), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n611), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT118), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(KEYINPUT118), .A3(new_n777), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n259), .A2(new_n780), .A3(new_n781), .A4(new_n261), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n237), .A2(new_n239), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(KEYINPUT119), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(KEYINPUT119), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n244), .B1(new_n243), .B2(new_n246), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n258), .B(new_n612), .C1(new_n787), .C2(new_n254), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n590), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n590), .A2(new_n781), .A3(new_n780), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n258), .B1(new_n787), .B2(new_n254), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n562), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n613), .A2(new_n262), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n496), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n690), .A2(new_n500), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT120), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n771), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n307), .B1(new_n798), .B2(new_n266), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT121), .B1(new_n802), .B2(new_n805), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1340gat));
  AOI211_X1 g608(.A(G120gat), .B(new_n639), .C1(new_n799), .C2(new_n801), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n308), .B1(new_n798), .B2(new_n612), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n810), .A2(new_n811), .ZN(G1341gat));
  INV_X1    g611(.A(new_n562), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n813), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n814), .A2(KEYINPUT122), .A3(new_n315), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT122), .B1(new_n814), .B2(new_n315), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n315), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(G1342gat));
  NAND2_X1  g617(.A1(new_n590), .A2(new_n484), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT123), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n795), .A2(new_n313), .A3(new_n615), .A4(new_n821), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT56), .Z(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n797), .B2(new_n641), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT124), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(KEYINPUT124), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  NAND2_X1  g626(.A1(new_n661), .A2(new_n796), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n793), .A2(new_n794), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n509), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n831), .B2(KEYINPUT57), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n776), .A2(KEYINPUT125), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT55), .B1(new_n776), .B2(KEYINPUT125), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(new_n778), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n264), .B2(new_n265), .ZN(new_n837));
  INV_X1    g636(.A(new_n788), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n641), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n792), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n813), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n794), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n509), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n832), .B1(new_n843), .B2(KEYINPUT57), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n380), .B1(new_n844), .B2(new_n266), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n415), .B1(new_n793), .B2(new_n794), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n631), .A3(new_n615), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n690), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n267), .A2(G141gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n828), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n835), .A2(new_n778), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n259), .A2(KEYINPUT93), .A3(new_n261), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT93), .B1(new_n259), .B2(new_n261), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n590), .B1(new_n858), .B2(new_n788), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n562), .B1(new_n859), .B2(new_n792), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n415), .B1(new_n860), .B2(new_n794), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n684), .B(new_n854), .C1(new_n861), .C2(new_n853), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n862), .A2(G141gat), .B1(new_n848), .B2(new_n849), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n845), .A2(new_n852), .B1(new_n863), .B2(new_n851), .ZN(G1344gat));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n382), .A3(new_n612), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G148gat), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n844), .B2(new_n612), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n613), .A2(new_n264), .A3(new_n265), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT126), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n853), .B(new_n509), .C1(new_n841), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n831), .A2(KEYINPUT57), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n872), .A2(new_n612), .A3(new_n829), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n866), .B1(new_n874), .B2(G148gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n865), .B1(new_n868), .B2(new_n875), .ZN(G1345gat));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n375), .A3(new_n813), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n844), .A2(new_n813), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n879), .B2(new_n375), .ZN(G1346gat));
  NAND2_X1  g679(.A1(new_n844), .A2(new_n590), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G162gat), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n821), .A2(new_n376), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n847), .B2(new_n883), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n615), .A2(new_n484), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT127), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n795), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(G169gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(new_n267), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n615), .B1(new_n793), .B2(new_n794), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n416), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n691), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n684), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n893), .B2(new_n888), .ZN(G1348gat));
  OAI21_X1  g693(.A(G176gat), .B1(new_n887), .B2(new_n639), .ZN(new_n895));
  OR3_X1    g694(.A1(new_n691), .A2(G176gat), .A3(new_n639), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n891), .B2(new_n896), .ZN(G1349gat));
  NAND3_X1  g696(.A1(new_n892), .A2(new_n268), .A3(new_n813), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n887), .B2(new_n562), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n892), .A2(new_n269), .A3(new_n590), .ZN(new_n902));
  OAI21_X1  g701(.A(G190gat), .B1(new_n887), .B2(new_n641), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(KEYINPUT61), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(KEYINPUT61), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(G1351gat));
  AND2_X1   g705(.A1(new_n872), .A2(new_n873), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n631), .A2(new_n886), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n907), .A2(G197gat), .A3(new_n266), .A4(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(G197gat), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n890), .A2(new_n631), .A3(new_n509), .A4(new_n690), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n262), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n909), .A2(new_n912), .ZN(G1352gat));
  NAND4_X1  g712(.A1(new_n872), .A2(new_n612), .A3(new_n873), .A4(new_n908), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G204gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n639), .A2(G204gat), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT62), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n911), .A2(KEYINPUT62), .A3(new_n917), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n918), .A3(new_n919), .ZN(G1353gat));
  NAND4_X1  g719(.A1(new_n872), .A2(new_n813), .A3(new_n873), .A4(new_n908), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n813), .A2(new_n366), .ZN(new_n924));
  OAI22_X1  g723(.A1(new_n922), .A2(new_n923), .B1(new_n911), .B2(new_n924), .ZN(G1354gat));
  AND3_X1   g724(.A1(new_n907), .A2(new_n590), .A3(new_n908), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n590), .A2(new_n367), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n926), .A2(new_n367), .B1(new_n911), .B2(new_n927), .ZN(G1355gat));
endmodule


