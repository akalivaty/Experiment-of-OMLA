//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n208), .B(new_n209), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n207), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n207), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n212), .B(new_n223), .C1(new_n214), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(new_n225), .A2(KEYINPUT0), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(KEYINPUT0), .B2(new_n225), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n221), .A2(new_n233), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n224), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G226), .B(G232), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n239), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n258), .B(G45), .C1(new_n256), .C2(KEYINPUT5), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT84), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT5), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT84), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(G270), .B(new_n255), .C1(new_n261), .C2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n255), .A2(G274), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n259), .A2(new_n260), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n263), .A2(KEYINPUT84), .A3(new_n265), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n268), .A2(new_n269), .A3(new_n257), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G257), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G264), .A2(G1698), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n255), .ZN(new_n278));
  OR2_X1    g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n277), .B(new_n278), .C1(G303), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n267), .A2(new_n271), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G1), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n285), .A2(G20), .B1(new_n258), .B2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(new_n226), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n287), .B2(new_n226), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n286), .B(G116), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n284), .A2(new_n227), .A3(G1), .ZN(new_n293));
  INV_X1    g0093(.A(G116), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n287), .A2(new_n226), .B1(G20), .B2(new_n294), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G283), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n227), .C1(G33), .C2(new_n213), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n296), .A2(KEYINPUT20), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT20), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n292), .B(new_n295), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n283), .A2(new_n301), .A3(G169), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT21), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n283), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(new_n301), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n267), .A2(G190), .A3(new_n271), .A4(new_n282), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n283), .A2(new_n301), .A3(KEYINPUT21), .A4(G169), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n267), .A2(G179), .A3(new_n271), .A4(new_n282), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n301), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n304), .A2(new_n308), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT88), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n302), .A2(new_n303), .B1(new_n311), .B2(new_n301), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n316), .A2(KEYINPUT88), .A3(new_n309), .A4(new_n308), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G107), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n293), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g0120(.A(new_n320), .B(KEYINPUT25), .Z(new_n321));
  NAND2_X1  g0121(.A1(new_n287), .A2(new_n226), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT70), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n289), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n286), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n321), .B1(new_n325), .B2(new_n319), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT23), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n227), .B2(G107), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n319), .A2(KEYINPUT23), .A3(G20), .ZN(new_n329));
  INV_X1    g0129(.A(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n294), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n328), .A2(new_n329), .B1(new_n331), .B2(new_n227), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n227), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n333), .A2(KEYINPUT22), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(KEYINPUT22), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT24), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT24), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n332), .C1(new_n334), .C2(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n290), .A2(new_n291), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n326), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(G250), .B(new_n272), .C1(new_n275), .C2(new_n276), .ZN(new_n343));
  OAI211_X1 g0143(.A(G257), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n344));
  INV_X1    g0144(.A(G294), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n343), .B(new_n344), .C1(new_n330), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n278), .ZN(new_n347));
  OAI211_X1 g0147(.A(G264), .B(new_n255), .C1(new_n261), .C2(new_n266), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n271), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G179), .B2(new_n349), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(G200), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n347), .A2(G190), .A3(new_n271), .A4(new_n348), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n324), .B1(new_n337), .B2(new_n339), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n356), .A2(new_n357), .A3(new_n326), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n318), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT79), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT78), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n281), .A2(new_n364), .A3(G226), .A4(G1698), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n275), .A2(new_n276), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G226), .A2(G1698), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT78), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(G1698), .B1(new_n279), .B2(new_n280), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n255), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n268), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G232), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n255), .A2(new_n373), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n363), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  INV_X1    g0180(.A(G274), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n278), .A2(new_n381), .A3(new_n373), .ZN(new_n382));
  INV_X1    g0182(.A(new_n377), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(G232), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(G223), .B(new_n272), .C1(new_n275), .C2(new_n276), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n330), .B2(new_n211), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n365), .B2(new_n368), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n380), .B(new_n384), .C1(new_n387), .C2(new_n255), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n379), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n279), .A2(new_n227), .A3(new_n280), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n280), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n203), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n202), .A2(new_n203), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G20), .A2(G33), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G159), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n390), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n366), .B2(new_n227), .ZN(new_n403));
  INV_X1    g0203(.A(new_n394), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n401), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n407), .A3(new_n341), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT8), .B(G58), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n293), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n324), .B1(G1), .B2(new_n227), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n409), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n362), .B1(new_n389), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n405), .A2(new_n406), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n324), .B1(new_n419), .B2(new_n390), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n415), .B1(new_n420), .B2(new_n407), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n379), .A2(new_n388), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(KEYINPUT79), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n361), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(G169), .B1(new_n372), .B2(new_n378), .ZN(new_n425));
  INV_X1    g0225(.A(G179), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n384), .B1(new_n387), .B2(new_n255), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n417), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT18), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n417), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n421), .A2(new_n422), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n361), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n424), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT80), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n272), .A2(G222), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G223), .A2(G1698), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n281), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n278), .C1(G77), .C2(new_n281), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n383), .A2(G226), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n375), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G179), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n350), .B2(new_n444), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n204), .A2(G20), .ZN(new_n447));
  INV_X1    g0247(.A(G150), .ZN(new_n448));
  INV_X1    g0248(.A(new_n399), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n227), .A2(G33), .ZN(new_n450));
  OAI221_X1 g0250(.A(new_n447), .B1(new_n448), .B2(new_n449), .C1(new_n450), .C2(new_n409), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n341), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n414), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n453), .A2(KEYINPUT71), .B1(G50), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT71), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n452), .A2(new_n456), .B1(new_n201), .B2(new_n293), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n446), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(KEYINPUT9), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT9), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n462), .A3(new_n457), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT76), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n444), .A2(new_n380), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n444), .A2(G200), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n466), .B1(new_n461), .B2(new_n463), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT10), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n461), .A2(new_n463), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT74), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT74), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n464), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n469), .B(KEYINPUT75), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT10), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n467), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n460), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT12), .ZN(new_n485));
  OAI21_X1  g0285(.A(G68), .B1(new_n454), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n203), .A2(G20), .ZN(new_n487));
  INV_X1    g0287(.A(G77), .ZN(new_n488));
  OAI221_X1 g0288(.A(new_n487), .B1(new_n450), .B2(new_n488), .C1(new_n449), .C2(new_n201), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n341), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n490), .A2(KEYINPUT11), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(KEYINPUT11), .ZN(new_n492));
  INV_X1    g0292(.A(new_n487), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n485), .A2(new_n284), .A3(G1), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n411), .A2(new_n485), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n486), .A2(new_n491), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n376), .A2(G1698), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n281), .B(new_n497), .C1(G226), .C2(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G97), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n255), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT13), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n382), .B1(G238), .B2(new_n383), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G238), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n375), .B1(new_n505), .B2(new_n377), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT13), .B1(new_n506), .B2(new_n500), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G169), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n509), .A2(KEYINPUT14), .B1(new_n426), .B2(new_n508), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n509), .A2(KEYINPUT14), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n496), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n508), .A2(new_n380), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(new_n496), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(G200), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(KEYINPUT77), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(KEYINPUT77), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G238), .A2(G1698), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n281), .B(new_n519), .C1(new_n376), .C2(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n278), .C1(G107), .C2(new_n281), .ZN(new_n521));
  INV_X1    g0321(.A(G244), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n375), .C1(new_n522), .C2(new_n377), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n380), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n449), .A2(KEYINPUT73), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n449), .A2(KEYINPUT73), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n527), .A2(new_n409), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g0329(.A(KEYINPUT15), .B(G87), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n530), .A2(new_n450), .B1(new_n227), .B2(new_n488), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n341), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n293), .A2(new_n488), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n533), .C1(new_n488), .C2(new_n414), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(G200), .B2(new_n523), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n525), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n523), .A2(G179), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n350), .B2(new_n523), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n534), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n512), .A2(new_n518), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n438), .A2(KEYINPUT81), .A3(new_n484), .A4(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n471), .A2(new_n465), .B1(G200), .B2(new_n444), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT76), .B1(new_n474), .B2(new_n466), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n480), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n481), .B1(new_n475), .B2(new_n477), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n540), .B(new_n459), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n389), .A2(new_n417), .A3(new_n362), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT79), .B1(new_n421), .B2(new_n422), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT17), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n432), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n431), .B1(new_n428), .B2(new_n417), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n553), .A3(new_n435), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n554), .B(KEYINPUT80), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n542), .B1(new_n547), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n541), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n293), .A2(new_n213), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n325), .B2(new_n213), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n319), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT6), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n564), .A2(new_n227), .B1(new_n488), .B2(new_n449), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n319), .B1(new_n393), .B2(new_n394), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n341), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n403), .B2(new_n404), .ZN(new_n570));
  AND2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G97), .A2(G107), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n563), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n319), .A2(KEYINPUT6), .A3(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(G20), .B1(G77), .B2(new_n399), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(KEYINPUT82), .A3(new_n341), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n560), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n272), .B1(new_n279), .B2(new_n280), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT83), .ZN(new_n582));
  OAI211_X1 g0382(.A(G244), .B(new_n272), .C1(new_n275), .C2(new_n276), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n370), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(G244), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n581), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n278), .ZN(new_n589));
  OAI211_X1 g0389(.A(G257), .B(new_n255), .C1(new_n261), .C2(new_n266), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n271), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G200), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n579), .B(new_n594), .C1(new_n380), .C2(new_n593), .ZN(new_n595));
  XOR2_X1   g0395(.A(KEYINPUT15), .B(G87), .Z(new_n596));
  INV_X1    g0396(.A(KEYINPUT86), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n530), .A2(KEYINPUT86), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n324), .A2(new_n598), .A3(new_n286), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n211), .A2(new_n213), .A3(new_n319), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n499), .A2(new_n227), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT19), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n227), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n450), .B2(new_n213), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n341), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n530), .A2(new_n293), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n600), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n212), .B1(new_n262), .B2(G1), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n258), .A2(new_n381), .A3(G45), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n255), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(G238), .A2(G1698), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n522), .B2(G1698), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n331), .B1(new_n615), .B2(new_n281), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n426), .B(new_n613), .C1(new_n616), .C2(new_n255), .ZN(new_n617));
  INV_X1    g0417(.A(new_n613), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n281), .ZN(new_n619));
  INV_X1    g0419(.A(new_n331), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n621), .B2(new_n278), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n610), .B(new_n617), .C1(G169), .C2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n613), .B1(new_n616), .B2(new_n255), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G200), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n607), .A2(new_n341), .B1(new_n293), .B2(new_n530), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n324), .A2(G87), .A3(new_n286), .ZN(new_n627));
  OAI211_X1 g0427(.A(G190), .B(new_n613), .C1(new_n616), .C2(new_n255), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n589), .A2(new_n592), .A3(G179), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n350), .B1(new_n589), .B2(new_n592), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n579), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI211_X1 g0434(.A(KEYINPUT85), .B(new_n560), .C1(new_n569), .C2(new_n578), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n595), .B(new_n630), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n560), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT82), .B1(new_n577), .B2(new_n341), .ZN(new_n640));
  AOI211_X1 g0440(.A(new_n568), .B(new_n324), .C1(new_n570), .C2(new_n576), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT85), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n579), .A2(new_n631), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n591), .B1(new_n278), .B2(new_n588), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G179), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n350), .B2(new_n645), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(KEYINPUT87), .A3(new_n595), .A4(new_n630), .ZN(new_n649));
  AOI211_X1 g0449(.A(new_n360), .B(new_n558), .C1(new_n638), .C2(new_n649), .ZN(G372));
  INV_X1    g0450(.A(new_n518), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n512), .B1(new_n651), .B2(new_n539), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n435), .A3(new_n550), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n553), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n473), .A2(new_n483), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n460), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n255), .A2(new_n611), .A3(new_n612), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n613), .A2(KEYINPUT89), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n658), .B(new_n659), .C1(new_n616), .C2(new_n255), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G200), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n350), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n610), .A3(new_n617), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n354), .A2(new_n355), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n342), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n667), .B(new_n595), .C1(new_n634), .C2(new_n635), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n648), .A2(KEYINPUT90), .A3(new_n595), .A4(new_n667), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n316), .B(new_n309), .C1(new_n342), .C2(new_n352), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n665), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n647), .A2(new_n674), .A3(new_n675), .A4(new_n642), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n664), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n643), .A2(new_n644), .A3(new_n647), .A4(new_n630), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(KEYINPUT26), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n656), .B1(new_n558), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT91), .ZN(G369));
  NAND2_X1  g0483(.A1(new_n285), .A2(new_n227), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n306), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n315), .B2(new_n317), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n316), .A2(new_n309), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  INV_X1    g0493(.A(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n359), .B1(new_n342), .B2(new_n689), .ZN(new_n696));
  INV_X1    g0496(.A(new_n353), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n689), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n692), .A2(new_n689), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT92), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n689), .B(KEYINPUT93), .Z(new_n702));
  AOI22_X1  g0502(.A1(new_n698), .A2(new_n701), .B1(new_n353), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  NOR2_X1   g0504(.A1(new_n223), .A2(G41), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n258), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n601), .A2(G116), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n230), .B2(new_n705), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  NAND2_X1  g0509(.A1(new_n680), .A2(new_n702), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n689), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n678), .A2(new_n675), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT94), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n678), .A2(KEYINPUT94), .A3(new_n675), .ZN(new_n717));
  AND4_X1   g0517(.A1(KEYINPUT26), .A2(new_n647), .A3(new_n642), .A4(new_n674), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n648), .A2(new_n595), .A3(new_n667), .A4(new_n672), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n664), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n713), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n712), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n318), .A2(new_n359), .A3(new_n702), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n638), .B2(new_n649), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n283), .A2(new_n426), .A3(new_n660), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n593), .A3(new_n349), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n622), .A2(new_n348), .A3(new_n347), .ZN(new_n731));
  NOR4_X1   g0531(.A1(new_n593), .A2(new_n731), .A3(KEYINPUT30), .A4(new_n310), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n731), .A2(new_n310), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n645), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n730), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n702), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n736), .A2(new_n713), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(KEYINPUT31), .ZN(new_n740));
  OAI21_X1  g0540(.A(G330), .B1(new_n728), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n726), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n709), .B1(new_n743), .B2(G1), .ZN(G364));
  NAND2_X1  g0544(.A1(new_n227), .A2(G13), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G45), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n706), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n693), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n226), .B1(G20), .B2(new_n350), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n223), .A2(new_n281), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n262), .B2(new_n230), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n252), .B2(new_n262), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n223), .A2(new_n366), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G355), .B1(new_n294), .B2(new_n223), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n227), .A2(new_n426), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n380), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(G190), .A3(new_n363), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(G322), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n426), .A2(G20), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n773), .A2(new_n380), .A3(new_n363), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n772), .A2(G311), .B1(new_n774), .B2(G303), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n281), .B(new_n776), .C1(G326), .C2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n773), .A2(G190), .A3(new_n363), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G283), .A2(new_n780), .B1(new_n781), .B2(G329), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  NAND2_X1  g0583(.A1(new_n363), .A2(G190), .ZN(new_n784));
  OAI21_X1  g0584(.A(G20), .B1(new_n784), .B2(G179), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT96), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n779), .B(new_n783), .C1(new_n345), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n213), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n767), .A2(new_n202), .ZN(new_n792));
  INV_X1    g0592(.A(new_n780), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n319), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(G87), .C2(new_n774), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n764), .A2(new_n203), .B1(new_n777), .B2(new_n201), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n366), .B(new_n796), .C1(G77), .C2(new_n772), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n781), .A2(G159), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT32), .Z(new_n799));
  NAND3_X1  g0599(.A1(new_n795), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n790), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n762), .B1(new_n801), .B2(new_n753), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n748), .B1(new_n752), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n693), .B(new_n694), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(new_n748), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT98), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  INV_X1    g0607(.A(new_n748), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n538), .A2(new_n534), .A3(new_n689), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n534), .A2(new_n713), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n536), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n812), .B2(new_n539), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n710), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n680), .A2(new_n702), .A3(new_n813), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n808), .B1(new_n817), .B2(new_n741), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n741), .B2(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(new_n753), .ZN(new_n820));
  INV_X1    g0620(.A(new_n774), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n201), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n793), .A2(new_n203), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n778), .A2(G137), .B1(new_n772), .B2(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G143), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n825), .B2(new_n767), .C1(new_n448), .C2(new_n764), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT34), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n822), .B(new_n823), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n366), .B1(new_n781), .B2(G132), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT100), .Z(new_n830));
  OR2_X1    g0630(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  INV_X1    g0631(.A(new_n789), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G58), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n828), .A2(new_n830), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n781), .ZN(new_n835));
  INV_X1    g0635(.A(G311), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n366), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n764), .A2(new_n838), .B1(new_n771), .B2(new_n294), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT99), .Z(new_n840));
  OAI22_X1  g0640(.A1(new_n793), .A2(new_n211), .B1(new_n345), .B2(new_n767), .ZN(new_n841));
  INV_X1    g0641(.A(G303), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n821), .A2(new_n319), .B1(new_n842), .B2(new_n777), .ZN(new_n843));
  OR4_X1    g0643(.A1(new_n837), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n834), .B1(new_n791), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n820), .B1(new_n845), .B2(KEYINPUT101), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(KEYINPUT101), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n753), .A2(new_n749), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n748), .B1(new_n488), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n813), .C2(new_n750), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n819), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n746), .A2(new_n258), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT40), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n417), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n408), .A2(new_n416), .A3(KEYINPUT103), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n428), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n418), .A3(new_n423), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n856), .A2(new_n688), .A3(new_n857), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n418), .A2(new_n423), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n417), .A2(new_n688), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n429), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n554), .A2(new_n860), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n496), .A2(new_n713), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n512), .A2(new_n518), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n512), .B2(new_n518), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n813), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n638), .A2(new_n649), .ZN(new_n877));
  INV_X1    g0677(.A(new_n727), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT31), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT105), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n736), .A2(new_n713), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n736), .B2(new_n713), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n879), .A2(KEYINPUT106), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT106), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n883), .A2(new_n884), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n728), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n876), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT107), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n872), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g0692(.A(KEYINPUT107), .B(new_n876), .C1(new_n886), .C2(new_n889), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n854), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n862), .A2(new_n865), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n434), .A2(new_n429), .A3(new_n863), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n437), .A2(new_n863), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n871), .A2(KEYINPUT104), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT104), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n867), .A2(new_n868), .A3(new_n901), .A4(KEYINPUT38), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n854), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n890), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n558), .B1(new_n889), .B2(new_n886), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n694), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n898), .A2(new_n899), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n902), .ZN(new_n912));
  INV_X1    g0712(.A(new_n871), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT39), .B1(new_n913), .B2(new_n869), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n512), .A2(new_n713), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n874), .A2(new_n875), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n809), .B(KEYINPUT102), .Z(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n816), .B2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n921), .A2(new_n872), .B1(new_n433), .B2(new_n687), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n557), .A2(new_n712), .A3(new_n725), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n656), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n853), .B1(new_n908), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n908), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(G116), .A4(new_n228), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n396), .A2(new_n229), .A3(new_n488), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n203), .A2(G50), .ZN(new_n934));
  OAI211_X1 g0734(.A(G1), .B(new_n284), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n928), .A2(new_n932), .A3(new_n935), .ZN(G367));
  OAI211_X1 g0736(.A(new_n648), .B(new_n595), .C1(new_n579), .C2(new_n702), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n647), .A2(new_n642), .A3(new_n737), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n698), .A2(new_n939), .A3(new_n701), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT42), .Z(new_n941));
  AOI21_X1  g0741(.A(new_n697), .B1(new_n937), .B2(new_n938), .ZN(new_n942));
  INV_X1    g0742(.A(new_n648), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n702), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n626), .A2(new_n627), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n713), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n674), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n664), .B2(new_n946), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n941), .A2(new_n944), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n699), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n939), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n705), .B(KEYINPUT41), .Z(new_n955));
  OR2_X1    g0755(.A1(new_n695), .A2(new_n698), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n699), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n701), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n743), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n703), .A2(new_n939), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT45), .Z(new_n962));
  OR3_X1    g0762(.A1(new_n703), .A2(KEYINPUT108), .A3(new_n939), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT108), .B1(new_n703), .B2(new_n939), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(KEYINPUT44), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT44), .B1(new_n963), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n952), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n967), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(new_n962), .A3(new_n699), .A4(new_n965), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n960), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n955), .B1(new_n971), .B2(new_n743), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n747), .A2(G1), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n954), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n239), .A2(new_n756), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n755), .B1(new_n223), .B2(new_n596), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n748), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n751), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n366), .B1(new_n780), .B2(G77), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT110), .Z(new_n980));
  INV_X1    g0780(.A(G137), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n821), .A2(new_n202), .B1(new_n835), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(G159), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n448), .A2(new_n767), .B1(new_n764), .B2(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n777), .A2(new_n825), .B1(new_n771), .B2(new_n201), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n980), .B(new_n986), .C1(new_n203), .C2(new_n789), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n789), .A2(new_n319), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n764), .A2(new_n345), .B1(new_n771), .B2(new_n838), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n281), .B(new_n989), .C1(G303), .C2(new_n768), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n793), .A2(new_n213), .B1(new_n835), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(KEYINPUT109), .B(G311), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(new_n778), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n774), .A2(G116), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n990), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n987), .B1(new_n988), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT47), .Z(new_n999));
  OAI221_X1 g0799(.A(new_n977), .B1(new_n978), .B2(new_n948), .C1(new_n999), .C2(new_n820), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n974), .A2(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n705), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n960), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n743), .B2(new_n958), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n707), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n760), .A2(new_n1005), .B1(new_n319), .B2(new_n223), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n244), .A2(new_n262), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n410), .A2(new_n201), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n707), .B(new_n262), .C1(new_n203), .C2(new_n488), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n756), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1006), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n748), .B1(new_n1012), .B2(new_n754), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n698), .B2(new_n978), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n366), .B1(new_n780), .B2(G97), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n821), .B2(new_n488), .C1(new_n448), .C2(new_n835), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT111), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n598), .A2(new_n599), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n789), .A2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n778), .A2(G159), .B1(new_n772), .B2(G68), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n410), .A2(new_n765), .B1(new_n768), .B2(G50), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n767), .A2(new_n991), .B1(new_n771), .B2(new_n842), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT112), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(KEYINPUT112), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n993), .A2(new_n765), .B1(new_n778), .B2(G322), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT113), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1029), .A2(KEYINPUT48), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(KEYINPUT48), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n789), .A2(new_n838), .B1(new_n345), .B2(new_n821), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n793), .A2(new_n294), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n281), .B(new_n1035), .C1(G326), .C2(new_n781), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1022), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1014), .B1(new_n1039), .B2(new_n753), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n958), .B2(new_n973), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1004), .A2(new_n1041), .ZN(G393));
  NAND3_X1  g0842(.A1(new_n968), .A2(new_n970), .A3(new_n973), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n249), .A2(new_n757), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n754), .B1(new_n213), .B2(new_n222), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n808), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n767), .A2(new_n983), .B1(new_n777), .B2(new_n448), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT51), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n832), .A2(G77), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n366), .B1(new_n780), .B2(G87), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n821), .A2(new_n203), .B1(new_n201), .B2(new_n764), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n835), .A2(new_n825), .B1(new_n409), .B2(new_n771), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n765), .A2(G303), .B1(G322), .B2(new_n781), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n838), .B2(new_n821), .C1(new_n345), .C2(new_n771), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1056), .A2(new_n281), .A3(new_n794), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n294), .B2(new_n789), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n767), .A2(new_n836), .B1(new_n777), .B2(new_n991), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT52), .Z(new_n1060));
  OAI21_X1  g0860(.A(new_n1054), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1046), .B1(new_n1061), .B2(new_n753), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n939), .B2(new_n978), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1043), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n971), .A2(new_n705), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n968), .A2(new_n970), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n959), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1064), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  AOI21_X1  g0869(.A(new_n694), .B1(new_n886), .B2(new_n889), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n876), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(G330), .B(new_n813), .C1(new_n728), .C2(new_n740), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n919), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n816), .A2(new_n920), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n919), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1070), .B2(new_n813), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n812), .A2(new_n539), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n810), .B1(new_n724), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n919), .B2(new_n1073), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1079), .A2(new_n1082), .A3(KEYINPUT114), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT114), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT106), .B1(new_n879), .B2(new_n885), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n728), .A2(new_n888), .A3(new_n887), .ZN(new_n1086));
  OAI211_X1 g0886(.A(G330), .B(new_n813), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n919), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1073), .A2(new_n919), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n678), .A2(KEYINPUT94), .A3(new_n675), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT94), .B1(new_n678), .B2(new_n675), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n1091), .A3(new_n718), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n689), .B(new_n1080), .C1(new_n1092), .C2(new_n722), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n809), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1084), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1077), .B1(new_n1083), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n557), .A2(new_n1070), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n924), .A2(new_n656), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n914), .B(new_n912), .C1(new_n921), .C2(new_n917), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n909), .A2(new_n902), .A3(new_n911), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n916), .C1(new_n1081), .C2(new_n919), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1089), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1072), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1072), .A2(new_n1074), .B1(new_n816), .B2(new_n920), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT114), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1088), .A2(new_n1084), .A3(new_n1095), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(new_n1099), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1116), .A3(new_n705), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n912), .A2(new_n749), .A3(new_n914), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n748), .B1(new_n409), .B2(new_n848), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT115), .Z(new_n1120));
  NAND2_X1  g0920(.A1(new_n832), .A2(G159), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n774), .A2(G150), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT53), .Z(new_n1123));
  AOI22_X1  g0923(.A1(G132), .A2(new_n768), .B1(new_n765), .B2(G137), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n778), .A2(G128), .B1(new_n772), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n366), .B1(new_n781), .B2(G125), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n201), .B2(new_n793), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT116), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT117), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n768), .A2(G116), .B1(G294), .B2(new_n781), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n319), .B2(new_n764), .C1(new_n838), .C2(new_n777), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n823), .B(new_n1136), .C1(G97), .C2(new_n772), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n281), .B1(new_n774), .B2(G87), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT118), .Z(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1049), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1133), .A2(KEYINPUT117), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1120), .B1(new_n1142), .B2(new_n753), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1118), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n973), .B2(new_n1115), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1117), .A2(new_n1146), .ZN(G378));
  OAI22_X1  g0947(.A1(new_n767), .A2(new_n319), .B1(new_n777), .B2(new_n294), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n366), .A2(new_n256), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G77), .B2(new_n774), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n202), .B2(new_n793), .C1(new_n213), .C2(new_n764), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1148), .B(new_n1151), .C1(G283), .C2(new_n781), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n203), .B2(new_n789), .C1(new_n1018), .C2(new_n771), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT58), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1149), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT120), .Z(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n778), .A2(G125), .B1(new_n774), .B2(new_n1126), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n981), .B2(new_n771), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G128), .A2(new_n768), .B1(new_n765), .B2(G132), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n448), .C2(new_n789), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n780), .A2(G159), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n781), .C2(G124), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n753), .B1(new_n1159), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT121), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n748), .B1(new_n201), .B2(new_n848), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n484), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n484), .A2(new_n1175), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1177), .A2(new_n458), .A3(new_n688), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n458), .A2(new_n688), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1178), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n1176), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1172), .B(new_n1173), .C1(new_n1183), .C2(new_n750), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT122), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n694), .B1(new_n903), .B2(new_n890), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n894), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1183), .B1(new_n894), .B2(new_n1186), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n923), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1183), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n913), .A2(new_n869), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1071), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(KEYINPUT107), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n890), .A2(new_n891), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT40), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n904), .A2(G330), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1190), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n923), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n894), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1189), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1185), .B1(new_n1201), .B2(new_n973), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1099), .B1(new_n1115), .B2(new_n1097), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1200), .B2(new_n1189), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n705), .B1(new_n1204), .B2(KEYINPUT57), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1100), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1201), .A2(KEYINPUT57), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1202), .B1(new_n1205), .B2(new_n1208), .ZN(G375));
  INV_X1    g1009(.A(new_n955), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1099), .B(new_n1077), .C1(new_n1083), .C2(new_n1096), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1101), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n919), .A2(new_n749), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n821), .A2(new_n983), .B1(new_n981), .B2(new_n767), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n366), .B(new_n1214), .C1(G58), .C2(new_n780), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n832), .A2(G50), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n772), .A2(G150), .B1(new_n781), .B2(G128), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1126), .A2(new_n765), .B1(new_n778), .B2(G132), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n767), .A2(new_n838), .B1(new_n771), .B2(new_n319), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n281), .B(new_n1220), .C1(G77), .C2(new_n780), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G97), .A2(new_n774), .B1(new_n781), .B2(G303), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n765), .A2(G116), .B1(new_n778), .B2(G294), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n1019), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n820), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n748), .B(new_n1225), .C1(new_n203), .C2(new_n848), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1097), .A2(new_n973), .B1(new_n1213), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1212), .A2(new_n1227), .ZN(G381));
  NAND3_X1  g1028(.A1(new_n1068), .A2(new_n974), .A3(new_n1000), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1230), .A2(new_n851), .A3(new_n1227), .A4(new_n1212), .ZN(new_n1231));
  OR4_X1    g1031(.A1(G378), .A2(G375), .A3(new_n1229), .A4(new_n1231), .ZN(G407));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  INV_X1    g1033(.A(G343), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(G213), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G375), .C2(new_n1237), .ZN(G409));
  INV_X1    g1038(.A(new_n1229), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1068), .B1(new_n974), .B2(new_n1000), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n806), .B1(new_n1004), .B2(new_n1041), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1239), .A2(new_n1240), .B1(new_n1230), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1230), .A2(new_n1241), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1229), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1202), .C1(new_n1205), .C2(new_n1208), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1187), .A2(new_n1188), .A3(new_n923), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1198), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT123), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1189), .A2(new_n1252), .A3(new_n1200), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1251), .A2(new_n973), .A3(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1201), .A2(new_n1210), .A3(new_n1206), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1185), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1233), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1236), .B1(new_n1248), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1236), .A2(G2897), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1211), .A2(KEYINPUT124), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT60), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1211), .A2(KEYINPUT124), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n705), .B1(new_n1113), .B2(new_n1099), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1268), .A2(G384), .A3(new_n1227), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1268), .B2(new_n1227), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1227), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n851), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1268), .A2(G384), .A3(new_n1227), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1260), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1247), .B1(new_n1259), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT62), .B1(new_n1259), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1277), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1248), .A2(new_n1258), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1235), .A3(new_n1279), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1282), .A2(KEYINPUT62), .A3(new_n1235), .A4(new_n1279), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(KEYINPUT125), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1246), .B1(new_n1281), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1282), .A2(new_n1235), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1276), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1283), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1293), .A3(new_n1246), .A4(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT126), .B1(new_n1288), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1283), .A2(new_n1278), .A3(new_n1284), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1286), .A2(KEYINPUT125), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1291), .B(new_n1298), .C1(new_n1299), .C2(new_n1280), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1246), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1295), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1297), .A2(new_n1304), .ZN(G405));
  INV_X1    g1105(.A(new_n1279), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1246), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1246), .A2(new_n1306), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT127), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1233), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1311), .A2(new_n1248), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1301), .A2(new_n1279), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1307), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1310), .A2(new_n1312), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1312), .B1(new_n1310), .B2(new_n1315), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


