//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT80), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n208), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n209), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT65), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(G183gat), .A3(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G183gat), .B(G190gat), .Z(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT24), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G183gat), .B(G190gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n230), .B1(new_n237), .B2(new_n229), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n235), .B1(new_n214), .B2(KEYINPUT23), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT27), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT27), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G183gat), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n254), .A3(new_n215), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n214), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n251), .A2(new_n249), .A3(KEYINPUT66), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n253), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT29), .B1(new_n243), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT77), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n207), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G211gat), .A2(G218gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(G211gat), .A2(G218gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(G197gat), .A2(G204gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(G197gat), .A2(G204gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G197gat), .B(G204gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n273), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT75), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n280), .B(new_n269), .C1(new_n272), .C2(new_n273), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT65), .B1(new_n224), .B2(new_n227), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n238), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT25), .B1(new_n285), .B2(new_n228), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n262), .B1(new_n286), .B2(new_n241), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n265), .ZN(new_n288));
  INV_X1    g087(.A(new_n265), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n241), .B1(new_n234), .B2(new_n235), .ZN(new_n290));
  INV_X1    g089(.A(new_n262), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT79), .B(new_n289), .C1(new_n292), .C2(KEYINPUT29), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n266), .A2(new_n283), .A3(new_n288), .A4(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT78), .B1(new_n287), .B2(new_n265), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n288), .B1(new_n263), .B2(new_n265), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(KEYINPUT78), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n279), .A2(KEYINPUT76), .A3(new_n281), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n206), .B(new_n294), .C1(new_n297), .C2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n294), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n265), .B1(new_n287), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n289), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT78), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n295), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n205), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n289), .B1(new_n292), .B2(KEYINPUT29), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(new_n288), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n301), .B1(new_n316), .B2(new_n295), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n317), .A2(KEYINPUT30), .A3(new_n206), .A4(new_n294), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n305), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT35), .ZN(new_n320));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G57gat), .B(G85gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n330));
  OAI21_X1  g129(.A(G120gat), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI22_X1  g134(.A1(KEYINPUT70), .A2(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n331), .A2(new_n335), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G113gat), .ZN(new_n340));
  INV_X1    g139(.A(G120gat), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT1), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G113gat), .A2(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G134gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G127gat), .ZN(new_n346));
  INV_X1    g145(.A(G127gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G141gat), .B(G148gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(G155gat), .B2(G162gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G141gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G148gat), .ZN(new_n359));
  INV_X1    g158(.A(G148gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G141gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G155gat), .B(G162gat), .ZN(new_n363));
  INV_X1    g162(.A(G155gat), .ZN(new_n364));
  INV_X1    g163(.A(G162gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT2), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n339), .A2(new_n350), .A3(new_n357), .A4(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n339), .A2(new_n350), .B1(new_n357), .B2(new_n367), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n328), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT5), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n368), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n342), .A2(new_n343), .B1(new_n346), .B2(new_n348), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n349), .A2(new_n334), .A3(new_n336), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n331), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n357), .A2(new_n367), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT82), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n368), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n373), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n357), .A2(new_n367), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT3), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n357), .A2(new_n367), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n339), .A2(new_n350), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n389), .A2(new_n327), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n372), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n369), .A2(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n368), .A2(new_n378), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n327), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT5), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n326), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n390), .A2(new_n398), .A3(new_n392), .A4(new_n393), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n379), .A2(KEYINPUT82), .B1(new_n368), .B2(new_n381), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n400), .B2(new_n373), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n399), .B(new_n325), .C1(new_n401), .C2(new_n372), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n397), .A2(KEYINPUT87), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n401), .B2(new_n372), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n326), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT6), .B1(new_n405), .B2(new_n326), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT87), .B1(new_n408), .B2(new_n402), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n320), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n319), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n387), .A2(new_n307), .ZN(new_n412));
  INV_X1    g211(.A(new_n300), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT76), .B1(new_n279), .B2(new_n281), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n386), .B1(new_n282), .B2(KEYINPUT29), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n384), .ZN(new_n417));
  INV_X1    g216(.A(G228gat), .ZN(new_n418));
  INV_X1    g217(.A(G233gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n282), .A2(new_n412), .ZN(new_n422));
  INV_X1    g221(.A(new_n278), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT84), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n422), .B1(new_n427), .B2(new_n377), .ZN(new_n428));
  INV_X1    g227(.A(new_n420), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G22gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT31), .B(G50gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G22gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n432), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n429), .B1(new_n301), .B2(new_n412), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n441), .A2(new_n417), .B1(new_n429), .B2(new_n428), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n440), .B1(new_n442), .B2(new_n437), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(KEYINPUT86), .A3(G22gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n421), .A2(new_n430), .A3(KEYINPUT85), .A4(new_n437), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n439), .B1(new_n448), .B2(new_n435), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n376), .B1(new_n290), .B2(new_n291), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n388), .B(new_n262), .C1(new_n286), .C2(new_n241), .ZN(new_n451));
  INV_X1    g250(.A(G227gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(new_n419), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n454), .B(KEYINPUT32), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n454), .B2(new_n455), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n454), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT71), .B1(new_n454), .B2(KEYINPUT32), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT72), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n466), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n460), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n451), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n452), .B2(new_n419), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT34), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n449), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n454), .A2(KEYINPUT32), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n454), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n466), .B1(new_n478), .B2(new_n461), .ZN(new_n479));
  INV_X1    g278(.A(new_n467), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n459), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n471), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n411), .A2(new_n473), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n411), .A2(new_n473), .A3(new_n485), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT73), .B1(new_n468), .B2(new_n472), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n489), .A3(new_n471), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(new_n473), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n408), .A2(new_n402), .ZN(new_n494));
  INV_X1    g293(.A(new_n406), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n319), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n488), .A2(new_n490), .A3(new_n473), .A4(KEYINPUT89), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n487), .B1(new_n499), .B2(KEYINPUT35), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n407), .A2(new_n409), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n303), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n317), .A2(new_n504), .A3(new_n294), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n205), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n297), .A2(new_n302), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n288), .B1(new_n308), .B2(KEYINPUT79), .ZN(new_n508));
  INV_X1    g307(.A(new_n293), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n282), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n504), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n503), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT37), .B1(new_n306), .B2(new_n312), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(KEYINPUT38), .A3(new_n205), .A4(new_n505), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n449), .ZN(new_n516));
  INV_X1    g315(.A(new_n319), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n392), .A2(new_n389), .A3(new_n393), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n328), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n369), .A2(new_n370), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n519), .B(KEYINPUT39), .C1(new_n328), .C2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n521), .B(new_n325), .C1(KEYINPUT39), .C2(new_n519), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT40), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n397), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n516), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  OAI22_X1  g326(.A1(new_n515), .A2(new_n527), .B1(new_n516), .B2(new_n497), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n468), .A2(new_n472), .ZN(new_n530));
  AOI211_X1 g329(.A(new_n460), .B(new_n471), .C1(new_n465), .C2(new_n467), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n468), .A2(new_n472), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n482), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n529), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n490), .A2(new_n488), .A3(KEYINPUT36), .A4(new_n535), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n528), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n500), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT16), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(G1gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G1gat), .B2(new_n543), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n546), .B(G8gat), .Z(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  INV_X1    g347(.A(G36gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT14), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT14), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT91), .ZN(new_n554));
  XOR2_X1   g353(.A(G43gat), .B(G50gat), .Z(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G43gat), .B(G50gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  NAND2_X1  g358(.A1(G29gat), .A2(G36gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT92), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564));
  INV_X1    g363(.A(new_n560), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n553), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(new_n559), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n562), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(new_n567), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(new_n564), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n547), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT93), .B1(new_n547), .B2(new_n572), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n563), .A2(new_n568), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n546), .B(G8gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n542), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n574), .A2(new_n580), .A3(KEYINPUT18), .A4(new_n582), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n576), .A2(new_n578), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n575), .A2(new_n579), .A3(KEYINPUT94), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n582), .B(KEYINPUT13), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n584), .B(new_n585), .C1(new_n590), .C2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G197gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT11), .B(G169gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT12), .Z(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT90), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n586), .ZN(new_n601));
  INV_X1    g400(.A(new_n589), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT94), .B1(new_n575), .B2(new_n579), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n591), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(new_n584), .A3(new_n585), .A4(new_n598), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(new_n606), .A3(KEYINPUT95), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT95), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n608), .A3(new_n599), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n541), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n364), .ZN(new_n613));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT21), .ZN(new_n617));
  AND2_X1   g416(.A1(G71gat), .A2(G78gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  XOR2_X1   g418(.A(G57gat), .B(G64gat), .Z(new_n620));
  AOI211_X1 g419(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(KEYINPUT9), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n618), .B1(KEYINPUT9), .B2(new_n619), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT96), .B(G57gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(G64gat), .ZN(new_n624));
  INV_X1    g423(.A(G64gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G57gat), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n622), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n547), .B1(new_n617), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(new_n628), .B2(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(G127gat), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n634), .A2(G127gat), .A3(new_n635), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n630), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n637), .A2(new_n630), .A3(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n616), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(new_n639), .A3(new_n615), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G85gat), .A2(G92gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  XOR2_X1   g448(.A(G99gat), .B(G106gat), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g450(.A1(G99gat), .A2(G106gat), .ZN(new_n652));
  INV_X1    g451(.A(G85gat), .ZN(new_n653));
  INV_X1    g452(.A(G92gat), .ZN(new_n654));
  AOI22_X1  g453(.A1(KEYINPUT8), .A2(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI211_X1 g457(.A(KEYINPUT99), .B(new_n650), .C1(new_n649), .C2(new_n655), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n570), .B2(new_n573), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(G232gat), .A2(G233gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n662), .A2(new_n576), .B1(KEYINPUT41), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(G190gat), .B(G218gat), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n661), .A2(new_n669), .A3(new_n665), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n664), .A2(KEYINPUT41), .ZN(new_n671));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT100), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n668), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n668), .B2(new_n670), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n621), .A2(new_n627), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n662), .A2(KEYINPUT10), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682));
  INV_X1    g481(.A(new_n658), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n656), .A2(new_n657), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n628), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n680), .B1(new_n658), .B2(new_n659), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n681), .B(new_n682), .C1(new_n687), .C2(KEYINPUT10), .ZN(new_n688));
  NAND2_X1  g487(.A1(G230gat), .A2(G233gat), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n662), .A2(KEYINPUT101), .A3(KEYINPUT10), .A4(new_n680), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT102), .ZN(new_n692));
  INV_X1    g491(.A(new_n689), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(G176gat), .B(G204gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n688), .A2(new_n698), .A3(new_n689), .A4(new_n690), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n692), .A2(new_n694), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n697), .ZN(new_n701));
  INV_X1    g500(.A(new_n691), .ZN(new_n702));
  INV_X1    g501(.A(new_n694), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n646), .A2(new_n679), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n611), .A2(new_n496), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g507(.A1(new_n611), .A2(new_n319), .A3(new_n706), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT16), .B(G8gat), .Z(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR4_X1   g511(.A1(new_n709), .A2(KEYINPUT103), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n709), .B2(G8gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n709), .A2(new_n712), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n715), .B2(KEYINPUT42), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n713), .B1(new_n716), .B2(new_n718), .ZN(G1325gat));
  NAND2_X1  g518(.A1(new_n611), .A2(new_n706), .ZN(new_n720));
  INV_X1    g519(.A(G15gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n538), .A2(new_n539), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n720), .B2(new_n536), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(G1326gat));
  NOR2_X1   g526(.A1(new_n720), .A2(new_n516), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT43), .B(G22gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  NOR3_X1   g529(.A1(new_n705), .A2(new_n645), .A3(new_n678), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT105), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n611), .A2(new_n548), .A3(new_n496), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT45), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n679), .B1(new_n500), .B2(new_n540), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(KEYINPUT44), .B(new_n679), .C1(new_n500), .C2(new_n540), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n610), .A2(new_n645), .A3(new_n705), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n739), .A2(new_n496), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n734), .B1(new_n548), .B2(new_n741), .ZN(G1328gat));
  AND3_X1   g541(.A1(new_n593), .A2(new_n608), .A3(new_n599), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n608), .B1(new_n593), .B2(new_n599), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n606), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n745), .B(new_n732), .C1(new_n500), .C2(new_n540), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n746), .A2(G36gat), .A3(new_n517), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT46), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n739), .A2(new_n319), .A3(new_n740), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n549), .ZN(G1329gat));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT106), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n536), .A2(G43gat), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n722), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n737), .A2(new_n756), .A3(new_n738), .A4(new_n740), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n755), .B1(new_n757), .B2(G43gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n751), .A2(KEYINPUT106), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1330gat));
  OR3_X1    g559(.A1(new_n746), .A2(G50gat), .A3(new_n516), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(KEYINPUT48), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n737), .A2(new_n449), .A3(new_n738), .A4(new_n740), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G50gat), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(G50gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n761), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n771), .ZN(G1331gat));
  NAND3_X1  g571(.A1(new_n705), .A2(new_n645), .A3(new_n678), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n541), .A2(new_n745), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n496), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(new_n623), .Z(G1332gat));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n774), .B(new_n319), .C1(new_n777), .C2(new_n625), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n625), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1333gat));
  INV_X1    g579(.A(G71gat), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n541), .A2(new_n745), .A3(new_n773), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(new_n536), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n756), .A2(G71gat), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n774), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n774), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT50), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n783), .B(new_n791), .C1(new_n787), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1334gat));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n449), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g594(.A1(new_n745), .A2(new_n645), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n705), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT109), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n737), .A2(new_n496), .A3(new_n738), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G85gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n802));
  INV_X1    g601(.A(new_n528), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n722), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n487), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n679), .A4(new_n796), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n679), .B(new_n796), .C1(new_n500), .C2(new_n540), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n705), .A2(new_n653), .A3(new_n496), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT111), .Z(new_n814));
  OAI22_X1  g613(.A1(new_n801), .A2(new_n802), .B1(new_n812), .B2(new_n814), .ZN(G1336gat));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n737), .A2(new_n319), .A3(new_n738), .A4(new_n798), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G92gat), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n705), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n517), .A2(new_n822), .A3(G92gat), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n808), .A2(new_n809), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND4_X1   g625(.A1(new_n817), .A2(new_n819), .A3(new_n821), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n820), .B1(new_n811), .B2(new_n823), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n817), .B1(new_n828), .B2(new_n819), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(G1337gat));
  NAND3_X1  g629(.A1(new_n739), .A2(new_n756), .A3(new_n798), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G99gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n536), .A2(G99gat), .A3(new_n822), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n811), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1338gat));
  NAND4_X1  g634(.A1(new_n737), .A2(new_n449), .A3(new_n738), .A4(new_n798), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G106gat), .ZN(new_n837));
  OR3_X1    g636(.A1(new_n822), .A2(new_n516), .A3(G106gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n812), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT53), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n837), .B(new_n841), .C1(new_n812), .C2(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1339gat));
  OAI211_X1 g642(.A(new_n592), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n581), .A2(new_n583), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n597), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n593), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n598), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n688), .A2(new_n690), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n693), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n692), .A2(new_n850), .A3(KEYINPUT54), .A4(new_n699), .ZN(new_n851));
  XNOR2_X1  g650(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n697), .B1(new_n702), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(KEYINPUT55), .A3(new_n853), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n848), .A2(new_n856), .A3(new_n700), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n645), .B1(new_n858), .B2(new_n679), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n679), .B1(new_n848), .B2(new_n705), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n607), .A2(new_n856), .A3(new_n609), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n700), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n822), .A2(new_n645), .A3(new_n678), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n745), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n706), .A2(new_n610), .A3(KEYINPUT113), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n319), .A2(new_n495), .A3(new_n494), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n530), .A2(new_n531), .A3(new_n449), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n610), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n493), .A2(new_n498), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n610), .A2(new_n330), .A3(new_n329), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT115), .Z(new_n880));
  OAI21_X1  g679(.A(new_n876), .B1(new_n878), .B2(new_n880), .ZN(G1340gat));
  INV_X1    g680(.A(new_n878), .ZN(new_n882));
  AOI21_X1  g681(.A(G120gat), .B1(new_n882), .B2(new_n705), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n822), .A2(new_n341), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n874), .B2(new_n884), .ZN(G1341gat));
  OAI21_X1  g684(.A(G127gat), .B1(new_n875), .B2(new_n646), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n882), .A2(new_n347), .A3(new_n645), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1342gat));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n345), .A3(new_n679), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n889), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT116), .B1(new_n889), .B2(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n345), .B1(new_n874), .B2(new_n679), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(KEYINPUT56), .B2(new_n889), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1343gat));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n870), .A2(KEYINPUT57), .A3(new_n449), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n859), .A2(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n516), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n722), .A2(new_n871), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n722), .A2(new_n871), .A3(KEYINPUT117), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n901), .A2(new_n745), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(G141gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n899), .A2(new_n516), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n722), .A3(new_n871), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(G141gat), .A3(new_n610), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n896), .B(KEYINPUT58), .C1(new_n907), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(G141gat), .B2(new_n906), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT118), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT58), .B1(new_n910), .B2(KEYINPUT119), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(KEYINPUT119), .B2(new_n910), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n911), .B(new_n914), .C1(new_n907), .C2(new_n916), .ZN(G1344gat));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n859), .A2(new_n863), .B1(new_n610), .B2(new_n706), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n898), .B1(new_n919), .B2(new_n516), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n897), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n921), .A2(new_n705), .A3(new_n904), .A4(new_n905), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G148gat), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n901), .A2(new_n705), .A3(new_n904), .A4(new_n905), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n360), .A2(KEYINPUT59), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n923), .A2(KEYINPUT59), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n909), .A2(G148gat), .A3(new_n822), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n927), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n922), .B2(G148gat), .ZN(new_n932));
  OAI211_X1 g731(.A(KEYINPUT120), .B(new_n929), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n933), .ZN(G1345gat));
  INV_X1    g733(.A(new_n909), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n364), .A3(new_n645), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n904), .A2(new_n905), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n900), .B2(new_n897), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(new_n645), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n939), .B2(new_n364), .ZN(G1346gat));
  AOI21_X1  g739(.A(KEYINPUT121), .B1(new_n938), .B2(new_n679), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n365), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(KEYINPUT121), .A3(new_n679), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n935), .A2(new_n365), .A3(new_n679), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1347gat));
  NOR3_X1   g745(.A1(new_n899), .A2(new_n496), .A3(new_n517), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n873), .ZN(new_n948));
  OAI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n610), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n877), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n745), .A2(new_n222), .A3(new_n223), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(G1348gat));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n877), .A3(new_n705), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT122), .A3(new_n209), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT122), .B1(new_n953), .B2(new_n209), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n705), .A2(G176gat), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n954), .A2(new_n955), .B1(new_n948), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1349gat));
  NOR2_X1   g758(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n960));
  INV_X1    g759(.A(new_n950), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n961), .A2(new_n245), .A3(new_n247), .A4(new_n645), .ZN(new_n962));
  OAI21_X1  g761(.A(G183gat), .B1(new_n948), .B2(new_n646), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT125), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n964), .B(new_n966), .ZN(G1350gat));
  OAI21_X1  g766(.A(G190gat), .B1(new_n948), .B2(new_n678), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT61), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n961), .A2(new_n248), .A3(new_n679), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1351gat));
  NOR3_X1   g770(.A1(new_n756), .A2(new_n496), .A3(new_n517), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n908), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974), .B2(new_n745), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n921), .A2(new_n972), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n745), .A2(G197gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(G1352gat));
  OR3_X1    g777(.A1(new_n973), .A2(G204gat), .A3(new_n822), .ZN(new_n979));
  XNOR2_X1  g778(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n976), .A2(new_n705), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G204gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(G1353gat));
  NOR3_X1   g784(.A1(new_n973), .A2(G211gat), .A3(new_n646), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n921), .A2(new_n645), .A3(new_n972), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  INV_X1    g792(.A(G218gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n974), .A2(new_n994), .A3(new_n679), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n976), .A2(new_n679), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n996), .B2(new_n994), .ZN(G1355gat));
endmodule


