//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT16), .B1(new_n192), .B2(G125), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(KEYINPUT73), .A3(G125), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G125), .B(G140), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT73), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n193), .B1(new_n198), .B2(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT75), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT68), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT68), .A2(G128), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .A4(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT23), .B1(new_n205), .B2(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G110), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT24), .B(G110), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(G128), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n205), .A2(G119), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n204), .A2(new_n208), .A3(KEYINPUT74), .A4(new_n209), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n212), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n192), .A2(G125), .ZN(new_n221));
  INV_X1    g035(.A(G125), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G140), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g038(.A(KEYINPUT16), .B(new_n194), .C1(new_n224), .C2(KEYINPUT73), .ZN(new_n225));
  INV_X1    g039(.A(new_n193), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n200), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n196), .A2(new_n200), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n201), .A2(new_n220), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n226), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n225), .A2(new_n200), .A3(new_n226), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n209), .B1(new_n204), .B2(new_n208), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  OR3_X1    g052(.A1(new_n216), .A2(new_n217), .A3(new_n213), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n231), .A2(new_n240), .A3(KEYINPUT76), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT76), .B1(new_n231), .B2(new_n240), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n191), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n231), .A2(new_n240), .ZN(new_n244));
  INV_X1    g058(.A(new_n191), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G217), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT70), .B(G902), .Z(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G234), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G902), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n254));
  INV_X1    g068(.A(new_n249), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n247), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n243), .A2(new_n246), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n249), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n250), .B(KEYINPUT71), .Z(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT2), .B(G113), .Z(new_n262));
  XNOR2_X1  g076(.A(G116), .B(G119), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  OR2_X1    g080(.A1(KEYINPUT66), .A2(G134), .ZN(new_n267));
  INV_X1    g081(.A(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT11), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT66), .A2(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G131), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n268), .A2(KEYINPUT11), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(G134), .B2(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n267), .A2(new_n270), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G137), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n200), .B2(G143), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(KEYINPUT64), .A3(G146), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n287));
  AND2_X1   g101(.A1(KEYINPUT68), .A2(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(KEYINPUT68), .A2(G128), .ZN(new_n289));
  OAI22_X1  g103(.A1(new_n281), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n200), .A2(G143), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n280), .A2(G146), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n285), .A2(new_n286), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT69), .B1(new_n279), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n293), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n280), .A2(KEYINPUT64), .A3(G146), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT64), .B1(new_n280), .B2(G146), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n291), .B(new_n286), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n275), .A4(new_n278), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(KEYINPUT0), .A2(G128), .ZN(new_n304));
  AND2_X1   g118(.A1(KEYINPUT0), .A2(G128), .ZN(new_n305));
  AOI211_X1 g119(.A(new_n304), .B(new_n305), .C1(new_n291), .C2(new_n292), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n291), .B(new_n305), .C1(new_n297), .C2(new_n298), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT65), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n285), .A2(new_n309), .A3(new_n305), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n275), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(KEYINPUT67), .A3(G131), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n266), .B1(new_n303), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n300), .A2(new_n275), .A3(new_n278), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n266), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n265), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G237), .A2(G953), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G210), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT27), .Z(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G101), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n303), .A2(new_n264), .A3(new_n317), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT31), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n311), .A2(new_n315), .A3(new_n316), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n295), .A2(new_n302), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n332), .A2(new_n333), .A3(new_n265), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT30), .B1(new_n332), .B2(new_n333), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n320), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n336), .B2(new_n265), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT31), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n328), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n317), .A2(new_n319), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n265), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n265), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n342), .B(new_n343), .C1(new_n340), .C2(new_n329), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n327), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(G472), .A2(G902), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(KEYINPUT32), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n328), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n322), .A2(new_n327), .A3(new_n329), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n265), .B1(new_n332), .B2(new_n333), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n329), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n342), .B1(new_n353), .B2(new_n340), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n328), .A2(KEYINPUT29), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n249), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G472), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT32), .B1(new_n346), .B2(new_n347), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n261), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n261), .B(new_n362), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G214), .B1(G237), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n368));
  OR2_X1    g182(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G104), .ZN(new_n371));
  AND2_X1   g185(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G107), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(G107), .ZN(new_n377));
  NOR2_X1   g191(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n373), .A2(new_n374), .A3(new_n376), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n370), .A2(G104), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n378), .B2(new_n377), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n374), .B1(new_n383), .B2(new_n373), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n368), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n376), .B1(new_n369), .B2(new_n371), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n378), .B1(new_n377), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(KEYINPUT81), .A3(new_n380), .A4(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(G101), .B(new_n393), .C1(new_n386), .C2(new_n388), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT83), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n264), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G113), .ZN(new_n399));
  INV_X1    g213(.A(G116), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n400), .A2(KEYINPUT5), .A3(G119), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n399), .B(new_n401), .C1(KEYINPUT5), .C2(new_n263), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n263), .B2(new_n262), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n377), .B2(new_n382), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n380), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G122), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n398), .A2(new_n407), .A3(new_n410), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT6), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(new_n398), .B2(new_n407), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n367), .B(new_n412), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n413), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n311), .A2(new_n222), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n294), .A2(new_n222), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n187), .A2(G224), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(G902), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n429));
  INV_X1    g243(.A(new_n423), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n422), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n405), .A2(KEYINPUT85), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n432), .A2(new_n403), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n403), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n410), .B(KEYINPUT8), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n423), .A2(KEYINPUT86), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n429), .B1(new_n423), .B2(KEYINPUT86), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n431), .B(new_n436), .C1(new_n422), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n413), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n428), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n426), .A2(new_n427), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n427), .B(KEYINPUT87), .Z(new_n445));
  AOI21_X1  g259(.A(new_n424), .B1(new_n416), .B2(new_n418), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n446), .B2(new_n442), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n366), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n449));
  OR2_X1    g263(.A1(KEYINPUT88), .A2(G143), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(G214), .A3(new_n323), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT88), .A2(G143), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G237), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n187), .A3(G214), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n272), .B(new_n451), .C1(new_n453), .C2(new_n456), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n450), .A2(new_n452), .B1(new_n323), .B2(G214), .ZN(new_n458));
  NOR2_X1   g272(.A1(KEYINPUT88), .A2(G143), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G131), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT17), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT17), .B(G131), .C1(new_n458), .C2(new_n460), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n233), .A2(new_n463), .A3(new_n234), .A4(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G113), .B(G122), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(new_n375), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n458), .A2(new_n460), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT18), .A2(G131), .ZN(new_n469));
  OAI211_X1 g283(.A(G146), .B(new_n194), .C1(new_n224), .C2(KEYINPUT73), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n230), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT18), .B(G131), .C1(new_n458), .C2(new_n460), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT89), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n230), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n451), .B(new_n469), .C1(new_n453), .C2(new_n456), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n474), .A2(new_n472), .A3(KEYINPUT89), .A4(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n465), .B(new_n467), .C1(new_n473), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n233), .A2(new_n234), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n463), .A2(new_n464), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n472), .A3(new_n475), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n480), .A2(new_n481), .B1(new_n484), .B2(new_n476), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT92), .B1(new_n485), .B2(new_n467), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n476), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n465), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n489));
  INV_X1    g303(.A(new_n467), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n479), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n449), .B1(new_n492), .B2(G902), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n485), .A2(KEYINPUT92), .A3(new_n467), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n478), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT93), .A3(new_n428), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n493), .A2(new_n497), .A3(G475), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n224), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n198), .B2(new_n500), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n502), .A2(new_n200), .B1(new_n461), .B2(new_n457), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n201), .A3(new_n229), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n467), .B1(new_n504), .B2(new_n487), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n499), .B1(new_n479), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n227), .B(KEYINPUT75), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n507), .A2(new_n503), .B1(new_n484), .B2(new_n476), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT90), .B(new_n478), .C1(new_n508), .C2(new_n467), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n511), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT91), .B1(new_n511), .B2(KEYINPUT20), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n479), .B2(new_n505), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n498), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n280), .A2(G128), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n214), .B2(new_n280), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n277), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n267), .A2(new_n270), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(new_n519), .C1(new_n214), .C2(new_n280), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G122), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(G116), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT94), .B(G122), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(new_n400), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(KEYINPUT94), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G122), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n400), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n529), .B(G107), .C1(new_n530), .C2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n526), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(G107), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n524), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT13), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n519), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n280), .A2(KEYINPUT13), .A3(G128), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n541), .B(new_n542), .C1(new_n214), .C2(new_n280), .ZN(new_n543));
  INV_X1    g357(.A(new_n519), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n288), .A2(new_n289), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(G143), .ZN(new_n546));
  AOI22_X1  g360(.A1(G134), .A2(new_n543), .B1(new_n546), .B2(new_n522), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n529), .A2(G107), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n370), .B(new_n527), .C1(new_n528), .C2(new_n400), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT9), .B(G234), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n552), .A2(new_n248), .A3(G953), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n539), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n539), .B2(new_n551), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n249), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n557), .A2(new_n560), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n518), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT95), .A3(new_n561), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G952), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  INV_X1    g383(.A(G234), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(new_n454), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n187), .B(new_n249), .C1(G234), .C2(G237), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT21), .B(G898), .Z(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT96), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G221), .B1(new_n552), .B2(G902), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G469), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n428), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n187), .A2(G227), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT79), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G140), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n315), .A2(new_n316), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n205), .B1(new_n291), .B2(KEYINPUT1), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n299), .B1(new_n285), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n380), .A3(new_n404), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n405), .A2(new_n294), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(KEYINPUT12), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n587), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n294), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n599), .A2(new_n590), .B1(new_n600), .B2(new_n406), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n385), .A2(new_n390), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n394), .A2(new_n396), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n311), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n598), .B(new_n601), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n586), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n587), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n586), .A2(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n582), .B1(new_n611), .B2(G469), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n597), .A2(new_n605), .A3(new_n607), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n607), .B1(new_n610), .B2(new_n605), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n581), .B(new_n249), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n580), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n448), .A2(new_n517), .A3(new_n578), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n364), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  AOI21_X1  g434(.A(new_n427), .B1(new_n426), .B2(new_n443), .ZN(new_n621));
  INV_X1    g435(.A(new_n427), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n446), .A2(new_n622), .A3(new_n442), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n365), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT97), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n622), .B1(new_n446), .B2(new_n442), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n444), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n365), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n511), .A2(KEYINPUT20), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT91), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n511), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n634), .A3(new_n516), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n493), .A2(new_n497), .A3(G475), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n554), .B2(new_n555), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n521), .A2(new_n523), .B1(new_n536), .B2(new_n537), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n643), .A2(new_n535), .B1(new_n547), .B2(new_n550), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n642), .B1(new_n644), .B2(new_n553), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n555), .A2(KEYINPUT99), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n553), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT33), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n649), .B(new_n639), .C1(new_n554), .C2(new_n555), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n255), .A2(new_n558), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n641), .A2(new_n648), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n556), .A2(new_n558), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n652), .B2(new_n653), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n638), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n641), .A2(new_n648), .A3(new_n650), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(KEYINPUT101), .A3(new_n654), .A4(new_n656), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n637), .A2(new_n662), .A3(new_n576), .ZN(new_n663));
  INV_X1    g477(.A(new_n347), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n330), .A2(KEYINPUT31), .B1(new_n327), .B2(new_n344), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(new_n339), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n346), .A2(new_n249), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(G472), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n261), .A3(new_n616), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n630), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT34), .B(G104), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  AND2_X1   g486(.A1(new_n567), .A2(new_n636), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n506), .A2(new_n509), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n515), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n514), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n673), .A2(new_n677), .A3(new_n576), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n630), .A2(new_n669), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT35), .B(G107), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n667), .A2(G472), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n346), .A2(new_n347), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT25), .B1(new_n257), .B2(new_n249), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n254), .B(new_n255), .C1(new_n243), .C2(new_n246), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n260), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n241), .A2(new_n242), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n251), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n682), .B1(new_n685), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n637), .A2(new_n567), .A3(new_n577), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n444), .A2(new_n447), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n697), .A2(new_n616), .A3(new_n365), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n668), .A2(KEYINPUT102), .A3(new_n693), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT37), .B(G110), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G12));
  AOI21_X1  g516(.A(new_n628), .B1(new_n627), .B2(new_n365), .ZN(new_n703));
  AOI211_X1 g517(.A(KEYINPUT97), .B(new_n366), .C1(new_n444), .C2(new_n626), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n616), .B(new_n693), .C1(new_n358), .C2(new_n359), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n571), .ZN(new_n708));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n708), .B1(new_n572), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n673), .A2(new_n677), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n705), .A2(new_n707), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G128), .ZN(G30));
  XOR2_X1   g529(.A(new_n710), .B(KEYINPUT39), .Z(new_n716));
  NAND2_X1  g530(.A1(new_n616), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT40), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n366), .A3(new_n693), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT104), .Z(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n697), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n444), .A2(new_n447), .A3(new_n721), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n337), .A2(new_n327), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n353), .A2(new_n327), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n428), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n666), .B2(KEYINPUT32), .ZN(new_n730));
  INV_X1    g544(.A(new_n348), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT32), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n684), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n348), .A4(new_n729), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n637), .A2(new_n567), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n719), .A2(new_n725), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G143), .ZN(G45));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n637), .A2(new_n662), .A3(new_n711), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(new_n630), .B2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n637), .A2(new_n662), .A3(new_n711), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n625), .A3(KEYINPUT106), .A4(new_n629), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n707), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G146), .ZN(G48));
  OAI21_X1  g561(.A(new_n249), .B1(new_n613), .B2(new_n614), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G469), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n615), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n580), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n261), .B(new_n751), .C1(new_n358), .C2(new_n359), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n663), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n705), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  INV_X1    g571(.A(new_n678), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n705), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  INV_X1    g574(.A(new_n751), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n703), .A2(new_n704), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n693), .B1(new_n358), .B2(new_n359), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n517), .A2(new_n578), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  NAND3_X1  g581(.A1(new_n738), .A2(new_n625), .A3(new_n629), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n750), .A2(new_n577), .A3(new_n580), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n340), .B1(new_n329), .B2(new_n352), .ZN(new_n771));
  INV_X1    g585(.A(new_n342), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n327), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n264), .B1(new_n335), .B2(new_n320), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n327), .A3(new_n334), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n770), .B(new_n773), .C1(new_n775), .C2(new_n338), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n339), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n770), .B1(new_n331), .B2(new_n773), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n347), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n769), .A2(new_n261), .A3(new_n683), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT108), .B1(new_n768), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n780), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n705), .A3(new_n783), .A4(new_n738), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G122), .ZN(G24));
  NAND3_X1  g600(.A1(new_n779), .A2(new_n683), .A3(new_n693), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n742), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n705), .A2(new_n788), .A3(new_n751), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G125), .ZN(G27));
  INV_X1    g604(.A(new_n360), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n616), .A2(new_n365), .A3(new_n447), .A4(new_n444), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n744), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n792), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n359), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n348), .B(new_n357), .C1(new_n359), .C2(new_n797), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n261), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n796), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n616), .A2(new_n365), .A3(new_n447), .A4(new_n444), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n742), .A2(new_n804), .A3(new_n794), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n688), .B1(new_n252), .B2(new_n247), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n797), .B1(new_n684), .B2(new_n733), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n358), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n808), .B2(new_n798), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT110), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n795), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G131), .ZN(G33));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n712), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n673), .A2(new_n677), .A3(KEYINPUT111), .A4(new_n711), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n791), .A3(new_n792), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G134), .ZN(G36));
  AND2_X1   g631(.A1(new_n658), .A2(new_n661), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT43), .B1(new_n818), .B2(new_n637), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT43), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n517), .A2(new_n820), .A3(new_n662), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(new_n685), .A3(new_n693), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT44), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n444), .A2(new_n365), .A3(new_n447), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n822), .B2(new_n823), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n607), .B1(new_n597), .B2(new_n605), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n608), .A2(new_n610), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT45), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT45), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n610), .A2(new_n605), .A3(new_n607), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n828), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n834), .A3(G469), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT112), .A4(G469), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n582), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(KEYINPUT46), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n615), .B1(new_n839), .B2(KEYINPUT46), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n579), .B(new_n716), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n824), .A2(new_n827), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(new_n268), .ZN(G39));
  NOR2_X1   g658(.A1(new_n358), .A2(new_n359), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n744), .A2(new_n806), .A3(new_n845), .A4(new_n826), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n579), .B1(new_n840), .B2(new_n841), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT47), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(KEYINPUT47), .B(new_n579), .C1(new_n840), .C2(new_n841), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(new_n192), .ZN(G42));
  AOI211_X1 g666(.A(new_n580), .B(new_n366), .C1(new_n750), .C2(KEYINPUT49), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(KEYINPUT49), .B2(new_n750), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n725), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n737), .A2(new_n806), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n517), .A4(new_n662), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n779), .A2(new_n683), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n806), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n819), .A3(new_n708), .A4(new_n821), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n630), .A3(new_n761), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n761), .A2(new_n571), .A3(new_n825), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n637), .A2(new_n662), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n569), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n761), .A2(new_n825), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n819), .A3(new_n708), .A4(new_n821), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n867), .A2(KEYINPUT48), .A3(new_n801), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT48), .B1(new_n867), .B2(new_n801), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n861), .B(new_n865), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n819), .A2(new_n708), .A3(new_n821), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  INV_X1    g686(.A(new_n787), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n866), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT116), .B1(new_n867), .B2(new_n787), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n637), .A2(new_n662), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n856), .A2(new_n862), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n749), .A2(new_n580), .A3(new_n615), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n849), .A2(new_n850), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n860), .A2(new_n825), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n723), .A2(new_n366), .A3(new_n724), .A4(new_n751), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n860), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n860), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT51), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n863), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n891), .A2(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n877), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n870), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n895));
  AND2_X1   g709(.A1(new_n884), .A2(new_n892), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n887), .A2(KEYINPUT115), .A3(new_n888), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT115), .B1(new_n887), .B2(new_n888), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n895), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n788), .A2(new_n792), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n562), .A2(new_n563), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n677), .A2(new_n636), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n616), .A2(new_n711), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n763), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n826), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n816), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n811), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n678), .A2(new_n703), .A3(new_n704), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n911), .A2(new_n753), .B1(new_n762), .B2(new_n765), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n663), .A2(new_n703), .A3(new_n704), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT102), .B1(new_n668), .B2(new_n693), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n617), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n913), .A2(new_n753), .B1(new_n915), .B2(new_n699), .ZN(new_n916));
  INV_X1    g730(.A(new_n903), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n517), .A2(KEYINPUT113), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT113), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n637), .B2(new_n903), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n920), .A3(new_n864), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n448), .A2(new_n576), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n669), .A2(new_n922), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n364), .A2(new_n618), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n785), .A2(new_n912), .A3(new_n916), .A4(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n910), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT52), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n745), .A2(new_n707), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT106), .B1(new_n705), .B2(new_n744), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n905), .A2(new_n693), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n705), .A2(new_n737), .A3(new_n738), .A4(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n714), .A3(new_n789), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n927), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n789), .A2(new_n714), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n746), .A3(KEYINPUT52), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n926), .A2(KEYINPUT53), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT53), .B1(new_n926), .B2(new_n937), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT53), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n934), .A2(new_n936), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n766), .A2(new_n755), .A3(new_n759), .A4(new_n700), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n921), .A2(new_n923), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n619), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n947), .A2(new_n785), .A3(new_n811), .A4(new_n909), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n942), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n926), .A2(KEYINPUT53), .A3(new_n937), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT54), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(KEYINPUT118), .B(new_n901), .C1(new_n941), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n568), .A2(new_n187), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n949), .A2(KEYINPUT54), .A3(new_n950), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT118), .B1(new_n957), .B2(new_n901), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n857), .B1(new_n954), .B2(new_n958), .ZN(G75));
  XNOR2_X1  g773(.A(new_n419), .B(new_n425), .ZN(new_n960));
  XNOR2_X1  g774(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(KEYINPUT56), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n255), .B1(new_n938), .B2(new_n939), .ZN(new_n965));
  INV_X1    g779(.A(new_n445), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n187), .A2(G952), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n249), .B1(new_n949), .B2(new_n950), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT56), .B1(new_n971), .B2(new_n622), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT120), .B1(new_n972), .B2(new_n962), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT56), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n965), .B2(new_n427), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT120), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n976), .A3(new_n963), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n970), .B1(new_n973), .B2(new_n977), .ZN(G51));
  XOR2_X1   g792(.A(new_n582), .B(KEYINPUT57), .Z(new_n979));
  OAI22_X1  g793(.A1(new_n957), .A2(new_n979), .B1(new_n614), .B2(new_n613), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n971), .A2(new_n837), .A3(new_n838), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n968), .B1(new_n980), .B2(new_n981), .ZN(G54));
  AND2_X1   g796(.A1(KEYINPUT58), .A2(G475), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n971), .A2(new_n675), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n675), .B1(new_n971), .B2(new_n983), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(new_n968), .ZN(G60));
  INV_X1    g800(.A(new_n659), .ZN(new_n987));
  NAND2_X1  g801(.A1(G478), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT59), .Z(new_n989));
  OAI21_X1  g803(.A(new_n987), .B1(new_n957), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n989), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n955), .A2(new_n956), .A3(new_n659), .A4(new_n991), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n990), .A2(new_n969), .A3(new_n992), .ZN(G63));
  NAND2_X1  g807(.A1(G217), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT60), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n949), .B2(new_n950), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(new_n257), .ZN(new_n997));
  INV_X1    g811(.A(new_n995), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n691), .B(new_n998), .C1(new_n938), .C2(new_n939), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n997), .A2(KEYINPUT61), .A3(new_n969), .A4(new_n999), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n999), .B(new_n969), .C1(new_n996), .C2(new_n257), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT61), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1000), .A2(new_n1003), .ZN(G66));
  AOI21_X1  g818(.A(new_n187), .B1(new_n575), .B2(G224), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT121), .ZN(new_n1006));
  INV_X1    g820(.A(new_n925), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT122), .Z(new_n1009));
  OAI211_X1 g823(.A(new_n416), .B(new_n418), .C1(G898), .C2(new_n187), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  XNOR2_X1  g825(.A(new_n336), .B(new_n502), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n935), .A2(new_n746), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1013), .A2(new_n1014), .A3(new_n739), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n843), .A2(new_n851), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n792), .A2(new_n716), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1017), .A2(new_n364), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1013), .A2(new_n739), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(KEYINPUT62), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT123), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1022), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1012), .B1(new_n1027), .B2(new_n187), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1012), .B1(new_n709), .B2(new_n187), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n809), .A2(new_n705), .A3(new_n738), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n842), .A2(new_n1030), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n811), .A2(new_n1031), .A3(new_n816), .ZN(new_n1032));
  AND3_X1   g846(.A1(new_n1016), .A2(new_n1032), .A3(new_n1013), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1029), .B1(new_n1033), .B2(new_n187), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT125), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  OR3_X1    g851(.A1(new_n1028), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1037), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  INV_X1    g854(.A(new_n726), .ZN(new_n1041));
  XNOR2_X1  g855(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1041), .A2(new_n350), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1045), .B1(new_n949), .B2(new_n950), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1021), .A2(new_n1025), .A3(new_n1007), .A4(new_n1026), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1041), .B1(new_n1047), .B2(new_n1044), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n1016), .A2(new_n1032), .A3(new_n1007), .A4(new_n1013), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n1049), .A2(new_n1044), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n969), .B1(new_n1050), .B2(new_n350), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT127), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g867(.A(KEYINPUT127), .B(new_n969), .C1(new_n1050), .C2(new_n350), .ZN(new_n1054));
  AOI211_X1 g868(.A(new_n1046), .B(new_n1048), .C1(new_n1053), .C2(new_n1054), .ZN(G57));
endmodule


