//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007;
  NAND2_X1  g000(.A1(G231gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT92), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G1gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT86), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G15gat), .B(G22gat), .Z(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT86), .B1(new_n216), .B2(new_n210), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n207), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n210), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(G8gat), .B1(new_n210), .B2(KEYINPUT86), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(KEYINPUT87), .A3(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n218), .A2(new_n223), .B1(G8gat), .B2(new_n219), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT21), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT9), .ZN(new_n226));
  INV_X1    g025(.A(G64gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G57gat), .ZN(new_n228));
  INV_X1    g027(.A(G57gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G64gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT90), .B1(G71gat), .B2(G78gat), .ZN(new_n232));
  INV_X1    g031(.A(G71gat), .ZN(new_n233));
  INV_X1    g032(.A(G78gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(KEYINPUT90), .A2(G71gat), .A3(G78gat), .ZN(new_n236));
  OR3_X1    g035(.A1(new_n231), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  OR3_X1    g036(.A1(new_n229), .A2(new_n227), .A3(KEYINPUT91), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n227), .B1(new_n229), .B2(KEYINPUT91), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n233), .A2(new_n234), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n226), .A2(G71gat), .A3(G78gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n238), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT93), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT93), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n245), .A3(new_n242), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n225), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n237), .A2(new_n242), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(KEYINPUT21), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n224), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n218), .A2(new_n223), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n219), .A2(G8gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n249), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n206), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G127gat), .B(G155gat), .Z(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  NAND3_X1  g059(.A1(new_n250), .A2(new_n255), .A3(new_n206), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n260), .ZN(new_n263));
  INV_X1    g062(.A(new_n261), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G78gat), .B(G106gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G22gat), .B(G50gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT31), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT79), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n274));
  INV_X1    g073(.A(G141gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G148gat), .ZN(new_n276));
  INV_X1    g075(.A(G148gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G141gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G155gat), .B(G162gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT2), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT73), .A4(new_n282), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n277), .A2(G141gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n275), .A2(G148gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(G155gat), .B2(G162gat), .ZN(new_n290));
  AND2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n285), .A2(new_n286), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n274), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT22), .ZN(new_n300));
  INV_X1    g099(.A(G211gat), .ZN(new_n301));
  INV_X1    g100(.A(G218gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G211gat), .B(G218gat), .Z(new_n305));
  OR2_X1    g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(new_n306), .B2(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n296), .ZN(new_n312));
  AND2_X1   g111(.A1(G228gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n296), .B2(KEYINPUT3), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n285), .A2(new_n295), .A3(KEYINPUT75), .A4(new_n286), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n319), .B(new_n320), .C1(new_n297), .C2(new_n311), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n310), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n316), .A2(new_n317), .B1(new_n322), .B2(new_n314), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n310), .A2(new_n315), .A3(KEYINPUT80), .A4(new_n312), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n273), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n317), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n314), .ZN(new_n327));
  AND4_X1   g126(.A1(new_n273), .A2(new_n326), .A3(new_n327), .A4(new_n324), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n272), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n324), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT79), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(new_n273), .A3(new_n324), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n271), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335));
  INV_X1    g134(.A(G85gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  OR2_X1    g138(.A1(new_n296), .A2(new_n297), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341));
  INV_X1    g140(.A(G120gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G113gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(G113gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G127gat), .ZN(new_n347));
  INV_X1    g146(.A(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G127gat), .A2(G134gat), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n342), .B2(G113gat), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n343), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT1), .B1(new_n349), .B2(new_n350), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n296), .A2(KEYINPUT3), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT4), .B1(new_n296), .B2(new_n360), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n346), .A2(new_n351), .B1(new_n357), .B2(new_n358), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n372), .A2(new_n286), .A3(new_n295), .A4(new_n285), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(KEYINPUT4), .B(new_n360), .C1(new_n319), .C2(new_n320), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  INV_X1    g177(.A(G155gat), .ZN(new_n379));
  INV_X1    g178(.A(G162gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n292), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n381), .A2(new_n281), .A3(new_n290), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n284), .A2(new_n283), .B1(new_n382), .B2(new_n289), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT75), .B1(new_n383), .B2(new_n286), .ZN(new_n384));
  INV_X1    g183(.A(new_n320), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n378), .B(new_n372), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(KEYINPUT78), .A3(new_n371), .A4(new_n374), .ZN(new_n387));
  AOI211_X1 g186(.A(new_n363), .B(new_n367), .C1(new_n377), .C2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n296), .B(new_n372), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT5), .B1(new_n389), .B2(new_n364), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n360), .B1(new_n319), .B2(new_n320), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT76), .B1(new_n391), .B2(new_n378), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n372), .B1(new_n384), .B2(new_n385), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT4), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n363), .A2(new_n365), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n390), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n339), .B1(new_n388), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(new_n390), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n387), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n373), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT77), .B1(new_n373), .B2(KEYINPUT4), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT78), .B1(new_n408), .B2(new_n386), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n362), .B(new_n366), .C1(new_n405), .C2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n339), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n400), .A2(new_n401), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT37), .ZN(new_n414));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT25), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT24), .ZN(new_n422));
  NOR2_X1   g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423));
  OAI22_X1  g222(.A1(new_n419), .A2(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n426), .A2(new_n427), .B1(KEYINPUT24), .B2(new_n421), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n417), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G169gat), .A2(G176gat), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT64), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n421), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT24), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n432), .A2(new_n425), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n423), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT24), .A3(new_n421), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT23), .ZN(new_n438));
  INV_X1    g237(.A(G169gat), .ZN(new_n439));
  INV_X1    g238(.A(G176gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n418), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(KEYINPUT25), .A3(new_n437), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n429), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT66), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT26), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT26), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(new_n439), .A3(new_n440), .A4(KEYINPUT66), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n446), .B(new_n448), .C1(new_n427), .C2(new_n426), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT27), .B(G183gat), .ZN(new_n450));
  INV_X1    g249(.A(G190gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(KEYINPUT28), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n449), .A2(new_n421), .A3(new_n454), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n416), .B1(new_n461), .B2(new_n274), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n459), .A2(new_n454), .A3(new_n421), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n463), .A2(new_n449), .B1(new_n429), .B2(new_n443), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n415), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT69), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n415), .B1(new_n464), .B2(KEYINPUT29), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n308), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n462), .A2(new_n465), .A3(new_n309), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT70), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n461), .A2(new_n416), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n468), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n309), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n471), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n414), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n477), .A3(new_n414), .ZN(new_n481));
  XNOR2_X1  g280(.A(G8gat), .B(G36gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(G92gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT71), .B(G64gat), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND2_X1  g284(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT38), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT6), .B(new_n339), .C1(new_n388), .C2(new_n399), .ZN(new_n488));
  INV_X1    g287(.A(new_n485), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n476), .A2(new_n477), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n308), .B1(new_n474), .B2(new_n475), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n462), .A2(new_n465), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n414), .B1(new_n493), .B2(new_n309), .ZN(new_n494));
  AOI211_X1 g293(.A(KEYINPUT38), .B(new_n489), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(new_n481), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n413), .A2(new_n487), .A3(new_n488), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT81), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n490), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT30), .A4(new_n489), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n489), .B1(new_n472), .B2(new_n479), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n470), .A2(KEYINPUT70), .A3(new_n471), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n478), .B1(new_n476), .B2(new_n477), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n485), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n507), .A2(KEYINPUT81), .A3(new_n500), .A4(new_n501), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n362), .B1(new_n405), .B2(new_n409), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT39), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n365), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n389), .B2(new_n364), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n363), .B1(new_n377), .B2(new_n387), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n364), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n515), .A3(new_n411), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n512), .A2(new_n515), .A3(KEYINPUT40), .A4(new_n411), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n400), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n334), .B(new_n497), .C1(new_n509), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n464), .A2(new_n360), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n461), .A2(new_n372), .ZN(new_n523));
  INV_X1    g322(.A(G227gat), .ZN(new_n524));
  INV_X1    g323(.A(G233gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT32), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G43gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n527), .B(KEYINPUT32), .C1(new_n529), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n523), .ZN(new_n538));
  INV_X1    g337(.A(new_n526), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT34), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT34), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n534), .A2(new_n541), .A3(new_n543), .A4(new_n536), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(KEYINPUT68), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n550), .A3(new_n546), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n537), .A2(KEYINPUT68), .A3(new_n544), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT36), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n413), .A2(new_n488), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n507), .A2(new_n500), .A3(new_n501), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n334), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n521), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n551), .A2(new_n552), .B1(new_n329), .B2(new_n333), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT35), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n334), .A2(new_n547), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n509), .A2(new_n555), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n571));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G134gat), .B(G162gat), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(G29gat), .A2(G36gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT14), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(KEYINPUT82), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n577), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT83), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n581), .A2(new_n582), .B1(G29gat), .B2(G36gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G43gat), .B(G50gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT15), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT15), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT84), .B(G43gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(G50gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT85), .B(G50gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(G43gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n589), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G29gat), .A2(G36gat), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n581), .A2(new_n587), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n585), .A2(new_n588), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(KEYINPUT17), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(KEYINPUT17), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n596), .A2(new_n594), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n587), .B1(new_n583), .B2(new_n584), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n598), .B(KEYINPUT17), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n606));
  XOR2_X1   g405(.A(G99gat), .B(G106gat), .Z(new_n607));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT7), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(G92gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n336), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n607), .A2(new_n608), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI211_X1 g416(.A(new_n608), .B(new_n607), .C1(new_n611), .C2(new_n614), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n606), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n607), .A2(new_n608), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n621), .A2(new_n611), .A3(new_n609), .A4(new_n614), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(KEYINPUT95), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n624), .B2(new_n597), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n576), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n619), .A2(new_n623), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n601), .B2(new_n604), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n631), .A2(new_n575), .A3(new_n627), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n574), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(new_n576), .A3(new_n628), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n575), .B1(new_n631), .B2(new_n627), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n573), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G113gat), .B(G141gat), .ZN(new_n638));
  INV_X1    g437(.A(G197gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT11), .B(G169gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n253), .B1(new_n601), .B2(new_n604), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n224), .A2(new_n597), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(KEYINPUT18), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n224), .B(new_n597), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n648), .B(KEYINPUT13), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n648), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n645), .A2(new_n655), .A3(new_n646), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(KEYINPUT18), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n644), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n647), .A2(new_n648), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT89), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT18), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n656), .A2(KEYINPUT18), .B1(new_n650), .B2(new_n652), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT89), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n643), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n244), .B2(new_n246), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n248), .A2(new_n620), .A3(new_n622), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n243), .B1(new_n617), .B2(new_n618), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n630), .A2(new_n669), .B1(new_n672), .B2(new_n668), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n667), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n668), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n244), .A2(new_n246), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n678), .A2(new_n623), .A3(new_n619), .A4(KEYINPUT10), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(KEYINPUT96), .A3(new_n674), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n672), .B2(new_n674), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT97), .A4(new_n675), .ZN(new_n685));
  XNOR2_X1  g484(.A(G120gat), .B(G148gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G204gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT98), .B(G176gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n685), .B(new_n684), .C1(new_n673), .C2(new_n675), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n682), .A2(new_n692), .B1(new_n693), .B2(new_n689), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n666), .A2(new_n695), .ZN(new_n696));
  AND4_X1   g495(.A1(new_n267), .A2(new_n569), .A3(new_n637), .A4(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n555), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT99), .B(G1gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1324gat));
  INV_X1    g500(.A(new_n509), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G8gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT16), .B(G8gat), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g506(.A(new_n705), .B(KEYINPUT42), .S(new_n707), .Z(G1325gat));
  AOI21_X1  g507(.A(G15gat), .B1(new_n697), .B2(new_n547), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n554), .A2(G15gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n697), .B2(new_n710), .ZN(G1326gat));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n559), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT100), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n714), .A2(KEYINPUT100), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n717), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n715), .A3(new_n712), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1327gat));
  INV_X1    g520(.A(new_n637), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n569), .A2(KEYINPUT44), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n521), .A2(new_n560), .B1(new_n564), .B2(new_n567), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n637), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n694), .B(KEYINPUT101), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n666), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n723), .A2(new_n726), .A3(new_n266), .A4(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n555), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n267), .A2(new_n637), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n555), .A2(G29gat), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n569), .A2(new_n696), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1328gat));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n666), .A3(new_n695), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n732), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n509), .A2(G36gat), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT103), .ZN(new_n745));
  OAI21_X1  g544(.A(G36gat), .B1(new_n730), .B2(new_n509), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n742), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(G1329gat));
  AND2_X1   g547(.A1(new_n549), .A2(new_n553), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n749), .A2(new_n590), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n730), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n741), .A2(new_n547), .A3(new_n732), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n752), .A2(new_n590), .B1(new_n753), .B2(KEYINPUT47), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n751), .B2(new_n754), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(G1330gat));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n759));
  INV_X1    g558(.A(new_n592), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n759), .B(new_n760), .C1(new_n730), .C2(new_n334), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n559), .A2(KEYINPUT106), .A3(new_n592), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n334), .B2(new_n760), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n759), .A3(new_n765), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n742), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n761), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n762), .B1(new_n761), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1331gat));
  NAND2_X1  g569(.A1(new_n658), .A2(new_n665), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n561), .B2(new_n568), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n727), .A2(new_n266), .A3(new_n722), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n555), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(new_n229), .ZN(G1332gat));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n509), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  AND2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n777), .B2(new_n778), .ZN(G1333gat));
  XNOR2_X1  g580(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n772), .A2(new_n547), .A3(new_n773), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(KEYINPUT107), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(KEYINPUT107), .ZN(new_n786));
  AOI21_X1  g585(.A(G71gat), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G71gat), .B1(new_n774), .B2(new_n749), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n786), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n233), .B1(new_n791), .B2(new_n784), .ZN(new_n792));
  INV_X1    g591(.A(new_n782), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n788), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(G1334gat));
  NOR2_X1   g594(.A1(new_n774), .A2(new_n334), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(new_n234), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n771), .A2(new_n694), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n723), .A2(new_n726), .A3(new_n266), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n555), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n772), .B2(new_n732), .ZN(new_n802));
  INV_X1    g601(.A(new_n732), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n771), .A4(new_n803), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n698), .A2(new_n336), .A3(new_n695), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(G1336gat));
  AOI21_X1  g606(.A(new_n556), .B1(new_n488), .B2(new_n413), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n749), .B1(new_n808), .B2(new_n334), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n509), .A2(new_n520), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n497), .A2(new_n334), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n566), .A2(new_n555), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n813), .A2(new_n509), .B1(new_n563), .B2(KEYINPUT35), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n666), .B(new_n732), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT110), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n802), .B2(new_n804), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(KEYINPUT110), .A3(new_n801), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n702), .A2(new_n613), .A3(new_n728), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT109), .Z(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G92gat), .B1(new_n799), .B2(new_n509), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n822), .B(new_n825), .C1(new_n805), .C2(new_n819), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(G1337gat));
  NOR2_X1   g626(.A1(new_n802), .A2(new_n804), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n694), .A2(G99gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n547), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G99gat), .B1(new_n799), .B2(new_n749), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT111), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1338gat));
  NOR3_X1   g635(.A1(new_n727), .A2(G106gat), .A3(new_n334), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n818), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G106gat), .B1(new_n799), .B2(new_n334), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n828), .B2(new_n837), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1339gat));
  AOI21_X1  g643(.A(new_n691), .B1(new_n676), .B2(new_n681), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n673), .B2(new_n675), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT96), .B1(new_n680), .B2(new_n674), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n667), .B(new_n675), .C1(new_n677), .C2(new_n679), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n673), .A2(new_n675), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n690), .B1(new_n851), .B2(new_n846), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n845), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  INV_X1    g655(.A(new_n647), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n655), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n856), .B(new_n655), .C1(new_n645), .C2(new_n646), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n650), .B2(new_n652), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n642), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT55), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n855), .A2(new_n665), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n267), .B1(new_n863), .B2(new_n722), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n665), .A2(new_n695), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n853), .A2(new_n854), .ZN(new_n866));
  INV_X1    g665(.A(new_n845), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n862), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n637), .B(new_n865), .C1(new_n666), .C2(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n267), .A2(new_n637), .A3(new_n694), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n864), .A2(new_n869), .B1(new_n666), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(new_n555), .A3(new_n702), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n562), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n355), .A3(new_n771), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n334), .A2(new_n547), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G113gat), .B1(new_n876), .B2(new_n666), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(G1340gat));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n342), .A3(new_n695), .ZN(new_n879));
  OAI21_X1  g678(.A(G120gat), .B1(new_n876), .B2(new_n727), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1341gat));
  NOR3_X1   g680(.A1(new_n876), .A2(new_n347), .A3(new_n266), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n873), .A2(new_n267), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n347), .B2(new_n883), .ZN(G1342gat));
  NAND3_X1  g683(.A1(new_n873), .A2(new_n348), .A3(new_n722), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n885), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT113), .B1(new_n885), .B2(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n888));
  OAI21_X1  g687(.A(G134gat), .B1(new_n876), .B2(new_n637), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(G1343gat));
  NAND2_X1  g689(.A1(new_n864), .A2(new_n869), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n666), .A2(new_n870), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n559), .ZN(new_n894));
  XOR2_X1   g693(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n871), .A2(new_n334), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n554), .A2(new_n555), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n509), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT114), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n896), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G141gat), .B1(new_n903), .B2(new_n666), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n771), .A2(new_n275), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n897), .A2(new_n907), .A3(new_n900), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n897), .B2(new_n900), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n509), .B(new_n906), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n509), .A3(new_n900), .A4(new_n906), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT116), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(new_n904), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n911), .ZN(G1344gat));
  OR2_X1    g715(.A1(new_n908), .A2(new_n909), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n917), .A2(new_n277), .A3(new_n509), .A4(new_n695), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n666), .B2(new_n870), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n267), .A2(new_n637), .A3(new_n694), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n771), .A2(new_n921), .A3(KEYINPUT118), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n891), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n924), .B2(new_n559), .ZN(new_n925));
  INV_X1    g724(.A(new_n895), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n871), .A2(new_n334), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n902), .A2(new_n695), .ZN(new_n929));
  OAI21_X1  g728(.A(G148gat), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT59), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n277), .A2(KEYINPUT59), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n903), .B2(new_n694), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n930), .B2(KEYINPUT59), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n918), .B1(new_n935), .B2(new_n936), .ZN(G1345gat));
  NOR3_X1   g736(.A1(new_n903), .A2(new_n379), .A3(new_n266), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n267), .A3(new_n509), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n379), .ZN(G1346gat));
  NAND4_X1  g739(.A1(new_n917), .A2(new_n380), .A3(new_n722), .A4(new_n509), .ZN(new_n941));
  OAI21_X1  g740(.A(G162gat), .B1(new_n903), .B2(new_n637), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1347gat));
  AND2_X1   g742(.A1(new_n702), .A2(new_n562), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT120), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n698), .B1(new_n944), .B2(KEYINPUT120), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n945), .A2(new_n893), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n439), .A3(new_n771), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n509), .A2(new_n698), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT121), .B1(new_n949), .B2(new_n547), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(new_n559), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(KEYINPUT121), .A3(new_n547), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n893), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n666), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n948), .A2(new_n954), .ZN(G1348gat));
  NAND3_X1  g754(.A1(new_n947), .A2(new_n440), .A3(new_n695), .ZN(new_n956));
  OAI21_X1  g755(.A(G176gat), .B1(new_n953), .B2(new_n727), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT122), .ZN(G1349gat));
  NAND3_X1  g758(.A1(new_n947), .A2(new_n267), .A3(new_n450), .ZN(new_n960));
  OAI21_X1  g759(.A(G183gat), .B1(new_n953), .B2(new_n266), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n451), .A3(new_n722), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n953), .A2(new_n637), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(G190gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n965), .B2(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1351gat));
  NAND2_X1  g768(.A1(new_n949), .A2(new_n749), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n894), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n639), .A3(new_n771), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT123), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n928), .A2(new_n970), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n771), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n976), .B2(new_n639), .ZN(G1352gat));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n334), .B1(new_n891), .B2(new_n923), .ZN(new_n979));
  OAI22_X1  g778(.A1(new_n894), .A2(new_n926), .B1(new_n979), .B2(KEYINPUT57), .ZN(new_n980));
  INV_X1    g779(.A(new_n970), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n980), .A2(new_n728), .A3(new_n981), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n694), .A2(G204gat), .ZN(new_n986));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n897), .A2(new_n981), .A3(new_n986), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT124), .B1(new_n988), .B2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n978), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n989), .A2(new_n990), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n982), .A2(G204gat), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT125), .A4(new_n987), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n992), .A2(new_n995), .ZN(G1353gat));
  NAND3_X1  g795(.A1(new_n971), .A2(new_n301), .A3(new_n267), .ZN(new_n997));
  OAI211_X1 g796(.A(new_n267), .B(new_n981), .C1(new_n925), .C2(new_n927), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n980), .A2(KEYINPUT126), .A3(new_n267), .A4(new_n981), .ZN(new_n1001));
  AND4_X1   g800(.A1(KEYINPUT63), .A2(new_n1000), .A3(G211gat), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n301), .B1(new_n998), .B2(new_n999), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1003), .B2(new_n1001), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n997), .B1(new_n1002), .B2(new_n1004), .ZN(G1354gat));
  AOI21_X1  g804(.A(G218gat), .B1(new_n971), .B2(new_n722), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n637), .A2(new_n302), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1006), .B1(new_n974), .B2(new_n1007), .ZN(G1355gat));
endmodule


