

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n587, n588, n589, n590, n591, n592, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752;

  AND2_X1 U365 ( .A1(n562), .A2(n561), .ZN(n388) );
  INV_X1 U366 ( .A(n495), .ZN(n702) );
  OR2_X1 U367 ( .A1(n664), .A2(G902), .ZN(n477) );
  BUF_X1 U368 ( .A(G143), .Z(n344) );
  XNOR2_X2 U369 ( .A(n342), .B(KEYINPUT39), .ZN(n606) );
  NAND2_X2 U370 ( .A1(n388), .A2(n389), .ZN(n342) );
  XNOR2_X1 U371 ( .A(n343), .B(n592), .ZN(n594) );
  NAND2_X1 U372 ( .A1(n590), .A2(n591), .ZN(n343) );
  XNOR2_X1 U373 ( .A(G134), .B(G116), .ZN(n418) );
  INV_X1 U374 ( .A(G953), .ZN(n744) );
  XNOR2_X2 U375 ( .A(n552), .B(KEYINPUT1), .ZN(n502) );
  AND2_X2 U376 ( .A1(n608), .A2(n607), .ZN(n610) );
  XNOR2_X2 U377 ( .A(n470), .B(n469), .ZN(n743) );
  INV_X1 U378 ( .A(KEYINPUT32), .ZN(n351) );
  AND2_X1 U379 ( .A1(n692), .A2(n357), .ZN(n370) );
  AND2_X1 U380 ( .A1(n702), .A2(n501), .ZN(n698) );
  XNOR2_X2 U381 ( .A(G113), .B(G116), .ZN(n398) );
  BUF_X1 U382 ( .A(n646), .Z(n662) );
  NAND2_X1 U383 ( .A1(n349), .A2(n350), .ZN(n347) );
  NAND2_X1 U384 ( .A1(n345), .A2(n346), .ZN(n348) );
  NAND2_X1 U385 ( .A1(n347), .A2(n348), .ZN(n508) );
  INV_X1 U386 ( .A(n349), .ZN(n345) );
  INV_X1 U387 ( .A(n350), .ZN(n346) );
  NOR2_X1 U388 ( .A1(n732), .A2(n518), .ZN(n349) );
  XNOR2_X1 U389 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n350) );
  XNOR2_X1 U390 ( .A(n352), .B(n351), .ZN(n657) );
  NOR2_X1 U391 ( .A1(n524), .A2(n496), .ZN(n352) );
  XNOR2_X2 U392 ( .A(n589), .B(n588), .ZN(n654) );
  NAND2_X1 U393 ( .A1(n376), .A2(n368), .ZN(n367) );
  NAND2_X1 U394 ( .A1(n371), .A2(KEYINPUT2), .ZN(n368) );
  XNOR2_X1 U395 ( .A(G902), .B(KEYINPUT15), .ZN(n609) );
  XNOR2_X1 U396 ( .A(G146), .B(G125), .ZN(n436) );
  OR2_X1 U397 ( .A1(n546), .A2(n545), .ZN(n585) );
  XNOR2_X1 U398 ( .A(n360), .B(n359), .ZN(n482) );
  XNOR2_X1 U399 ( .A(KEYINPUT96), .B(KEYINPUT24), .ZN(n360) );
  XNOR2_X1 U400 ( .A(G122), .B(G104), .ZN(n431) );
  XNOR2_X1 U401 ( .A(n344), .B(G113), .ZN(n432) );
  XNOR2_X1 U402 ( .A(G107), .B(G104), .ZN(n402) );
  NAND2_X1 U403 ( .A1(n365), .A2(n363), .ZN(n362) );
  INV_X1 U404 ( .A(KEYINPUT84), .ZN(n374) );
  NOR2_X1 U405 ( .A1(n721), .A2(KEYINPUT47), .ZN(n383) );
  AND2_X1 U406 ( .A1(n381), .A2(n380), .ZN(n379) );
  NOR2_X1 U407 ( .A1(n382), .A2(n680), .ZN(n381) );
  AND2_X1 U408 ( .A1(n721), .A2(KEYINPUT47), .ZN(n382) );
  XNOR2_X1 U409 ( .A(n385), .B(n384), .ZN(n581) );
  INV_X1 U410 ( .A(KEYINPUT73), .ZN(n384) );
  NAND2_X1 U411 ( .A1(n379), .A2(n377), .ZN(n385) );
  NAND2_X1 U412 ( .A1(n378), .A2(n383), .ZN(n377) );
  XNOR2_X1 U413 ( .A(KEYINPUT95), .B(KEYINPUT23), .ZN(n359) );
  AND2_X1 U414 ( .A1(n364), .A2(KEYINPUT65), .ZN(n363) );
  INV_X1 U415 ( .A(KEYINPUT2), .ZN(n364) );
  NAND2_X1 U416 ( .A1(n609), .A2(n371), .ZN(n369) );
  XNOR2_X1 U417 ( .A(n436), .B(n393), .ZN(n396) );
  XNOR2_X1 U418 ( .A(n392), .B(KEYINPUT17), .ZN(n393) );
  INV_X1 U419 ( .A(KEYINPUT76), .ZN(n392) );
  NAND2_X1 U420 ( .A1(n648), .A2(n609), .ZN(n564) );
  INV_X1 U421 ( .A(G902), .ZN(n490) );
  NOR2_X1 U422 ( .A1(G953), .A2(n730), .ZN(n413) );
  XOR2_X1 U423 ( .A(G122), .B(G107), .Z(n419) );
  XOR2_X1 U424 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n421) );
  NAND2_X1 U425 ( .A1(n411), .A2(n356), .ZN(n576) );
  XNOR2_X1 U426 ( .A(n564), .B(n409), .ZN(n411) );
  INV_X1 U427 ( .A(n563), .ZN(n409) );
  XNOR2_X1 U428 ( .A(n576), .B(KEYINPUT19), .ZN(n554) );
  BUF_X1 U429 ( .A(n559), .Z(n707) );
  XNOR2_X1 U430 ( .A(KEYINPUT16), .B(G122), .ZN(n401) );
  XNOR2_X1 U431 ( .A(n489), .B(n488), .ZN(n658) );
  XNOR2_X1 U432 ( .A(n440), .B(n439), .ZN(n635) );
  XNOR2_X1 U433 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U434 ( .A(n743), .B(n474), .ZN(n664) );
  AND2_X1 U435 ( .A1(n615), .A2(G953), .ZN(n667) );
  XNOR2_X1 U436 ( .A(n373), .B(KEYINPUT75), .ZN(n696) );
  NAND2_X1 U437 ( .A1(n612), .A2(n361), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n611), .B(n374), .ZN(n361) );
  XOR2_X1 U439 ( .A(G140), .B(G110), .Z(n353) );
  XOR2_X1 U440 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n354) );
  AND2_X1 U441 ( .A1(n449), .A2(n501), .ZN(n355) );
  NAND2_X1 U442 ( .A1(n410), .A2(G214), .ZN(n356) );
  INV_X1 U443 ( .A(n609), .ZN(n376) );
  AND2_X1 U444 ( .A1(n376), .A2(n371), .ZN(n357) );
  AND2_X1 U445 ( .A1(n369), .A2(n367), .ZN(n358) );
  INV_X1 U446 ( .A(G140), .ZN(n630) );
  NOR2_X2 U447 ( .A1(n651), .A2(n667), .ZN(n653) );
  NOR2_X2 U448 ( .A1(n638), .A2(n667), .ZN(n639) );
  NAND2_X1 U449 ( .A1(n366), .A2(n362), .ZN(n375) );
  AND2_X2 U450 ( .A1(n375), .A2(n372), .ZN(n646) );
  INV_X1 U451 ( .A(n696), .ZN(n372) );
  NOR2_X2 U452 ( .A1(n619), .A2(n741), .ZN(n692) );
  NAND2_X1 U453 ( .A1(n548), .A2(n495), .ZN(n549) );
  XNOR2_X2 U454 ( .A(n494), .B(n386), .ZN(n495) );
  INV_X1 U455 ( .A(n692), .ZN(n365) );
  NOR2_X1 U456 ( .A1(n370), .A2(n358), .ZN(n366) );
  INV_X1 U457 ( .A(KEYINPUT65), .ZN(n371) );
  INV_X1 U458 ( .A(n682), .ZN(n378) );
  NAND2_X1 U459 ( .A1(n682), .A2(KEYINPUT47), .ZN(n380) );
  XOR2_X1 U460 ( .A(n493), .B(n492), .Z(n386) );
  AND2_X1 U461 ( .A1(n507), .A2(n567), .ZN(n387) );
  AND2_X1 U462 ( .A1(n716), .A2(n585), .ZN(n389) );
  XNOR2_X1 U463 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U464 ( .A(n458), .B(n457), .ZN(n463) );
  XNOR2_X1 U465 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U466 ( .A(n444), .B(n443), .ZN(n567) );
  INV_X1 U467 ( .A(n667), .ZN(n616) );
  XNOR2_X2 U468 ( .A(KEYINPUT79), .B(G143), .ZN(n390) );
  XNOR2_X2 U469 ( .A(n390), .B(G128), .ZN(n427) );
  XNOR2_X1 U470 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n391) );
  XNOR2_X2 U471 ( .A(n427), .B(n391), .ZN(n464) );
  NAND2_X1 U472 ( .A1(n744), .A2(G224), .ZN(n394) );
  XNOR2_X1 U473 ( .A(n394), .B(KEYINPUT18), .ZN(n395) );
  XNOR2_X1 U474 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U475 ( .A(n464), .B(n397), .ZN(n406) );
  INV_X1 U476 ( .A(n398), .ZN(n400) );
  XNOR2_X1 U477 ( .A(KEYINPUT3), .B(G119), .ZN(n399) );
  XNOR2_X1 U478 ( .A(n400), .B(n399), .ZN(n461) );
  XNOR2_X1 U479 ( .A(n461), .B(n401), .ZN(n405) );
  XNOR2_X1 U480 ( .A(n402), .B(G110), .ZN(n404) );
  XNOR2_X1 U481 ( .A(G101), .B(KEYINPUT90), .ZN(n403) );
  XNOR2_X1 U482 ( .A(n404), .B(n403), .ZN(n473) );
  XNOR2_X1 U483 ( .A(n405), .B(n473), .ZN(n627) );
  XNOR2_X1 U484 ( .A(n406), .B(n627), .ZN(n648) );
  INV_X1 U485 ( .A(G237), .ZN(n407) );
  NAND2_X1 U486 ( .A1(n490), .A2(n407), .ZN(n410) );
  NAND2_X1 U487 ( .A1(n410), .A2(G210), .ZN(n408) );
  XNOR2_X1 U488 ( .A(n408), .B(KEYINPUT80), .ZN(n563) );
  NAND2_X1 U489 ( .A1(G234), .A2(G237), .ZN(n412) );
  XNOR2_X1 U490 ( .A(n354), .B(n412), .ZN(n414) );
  NAND2_X1 U491 ( .A1(G952), .A2(n414), .ZN(n730) );
  XNOR2_X1 U492 ( .A(n413), .B(KEYINPUT92), .ZN(n546) );
  NAND2_X1 U493 ( .A1(G902), .A2(n414), .ZN(n543) );
  XNOR2_X1 U494 ( .A(G898), .B(KEYINPUT93), .ZN(n623) );
  NAND2_X1 U495 ( .A1(G953), .A2(n623), .ZN(n626) );
  NOR2_X1 U496 ( .A1(n543), .A2(n626), .ZN(n415) );
  OR2_X1 U497 ( .A1(n546), .A2(n415), .ZN(n416) );
  NAND2_X1 U498 ( .A1(n554), .A2(n416), .ZN(n417) );
  XNOR2_X2 U499 ( .A(n417), .B(KEYINPUT0), .ZN(n518) );
  INV_X1 U500 ( .A(n518), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n419), .B(n418), .ZN(n423) );
  XNOR2_X1 U502 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n420) );
  XNOR2_X1 U503 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U504 ( .A(n423), .B(n422), .Z(n426) );
  NAND2_X1 U505 ( .A1(G234), .A2(n744), .ZN(n424) );
  XOR2_X1 U506 ( .A(KEYINPUT8), .B(n424), .Z(n479) );
  NAND2_X1 U507 ( .A1(G217), .A2(n479), .ZN(n425) );
  XNOR2_X1 U508 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U509 ( .A(n427), .B(n428), .ZN(n613) );
  NAND2_X1 U510 ( .A1(n613), .A2(n490), .ZN(n430) );
  INV_X1 U511 ( .A(G478), .ZN(n429) );
  XNOR2_X1 U512 ( .A(n430), .B(n429), .ZN(n566) );
  INV_X1 U513 ( .A(n566), .ZN(n507) );
  XNOR2_X1 U514 ( .A(n630), .B(G131), .ZN(n467) );
  XNOR2_X1 U515 ( .A(n431), .B(n467), .ZN(n435) );
  XOR2_X1 U516 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n433) );
  XNOR2_X1 U517 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U518 ( .A(n435), .B(n434), .Z(n440) );
  XNOR2_X1 U519 ( .A(KEYINPUT10), .B(n436), .ZN(n742) );
  INV_X1 U520 ( .A(n742), .ZN(n438) );
  NOR2_X1 U521 ( .A1(G953), .A2(G237), .ZN(n459) );
  NAND2_X1 U522 ( .A1(G214), .A2(n459), .ZN(n437) );
  NAND2_X1 U523 ( .A1(n635), .A2(n490), .ZN(n444) );
  XOR2_X1 U524 ( .A(KEYINPUT13), .B(KEYINPUT105), .Z(n442) );
  XNOR2_X1 U525 ( .A(KEYINPUT104), .B(G475), .ZN(n441) );
  XOR2_X1 U526 ( .A(n442), .B(n441), .Z(n443) );
  OR2_X1 U527 ( .A1(n507), .A2(n567), .ZN(n719) );
  INV_X1 U528 ( .A(n719), .ZN(n449) );
  NAND2_X1 U529 ( .A1(G234), .A2(n609), .ZN(n445) );
  XNOR2_X1 U530 ( .A(KEYINPUT20), .B(n445), .ZN(n491) );
  NAND2_X1 U531 ( .A1(n491), .A2(G221), .ZN(n447) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n446) );
  XNOR2_X1 U533 ( .A(n447), .B(n446), .ZN(n703) );
  INV_X1 U534 ( .A(KEYINPUT99), .ZN(n448) );
  XNOR2_X1 U535 ( .A(n703), .B(n448), .ZN(n501) );
  NAND2_X1 U536 ( .A1(n450), .A2(n355), .ZN(n452) );
  INV_X1 U537 ( .A(KEYINPUT22), .ZN(n451) );
  XNOR2_X1 U538 ( .A(n452), .B(n451), .ZN(n499) );
  XOR2_X1 U539 ( .A(KEYINPUT5), .B(KEYINPUT101), .Z(n454) );
  XNOR2_X1 U540 ( .A(G146), .B(G131), .ZN(n453) );
  XNOR2_X1 U541 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X1 U542 ( .A(G137), .B(G101), .ZN(n456) );
  INV_X1 U543 ( .A(KEYINPUT74), .ZN(n455) );
  NAND2_X1 U544 ( .A1(n459), .A2(G210), .ZN(n460) );
  XNOR2_X1 U545 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U546 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X2 U547 ( .A(n464), .B(G134), .ZN(n470) );
  XNOR2_X1 U548 ( .A(n470), .B(n465), .ZN(n640) );
  NAND2_X1 U549 ( .A1(n640), .A2(n490), .ZN(n466) );
  XNOR2_X1 U550 ( .A(n466), .B(G472), .ZN(n559) );
  XNOR2_X1 U551 ( .A(n707), .B(KEYINPUT6), .ZN(n572) );
  NAND2_X1 U552 ( .A1(n499), .A2(n572), .ZN(n524) );
  XNOR2_X1 U553 ( .A(KEYINPUT67), .B(G137), .ZN(n486) );
  XNOR2_X1 U554 ( .A(n486), .B(KEYINPUT94), .ZN(n468) );
  XNOR2_X1 U555 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U556 ( .A1(n744), .A2(G227), .ZN(n471) );
  XNOR2_X1 U557 ( .A(n471), .B(G146), .ZN(n472) );
  XNOR2_X1 U558 ( .A(n473), .B(n472), .ZN(n474) );
  INV_X1 U559 ( .A(KEYINPUT71), .ZN(n475) );
  XNOR2_X1 U560 ( .A(n475), .B(G469), .ZN(n476) );
  XNOR2_X2 U561 ( .A(n477), .B(n476), .ZN(n552) );
  INV_X1 U562 ( .A(n502), .ZN(n478) );
  INV_X1 U563 ( .A(n478), .ZN(n699) );
  XNOR2_X1 U564 ( .A(n699), .B(KEYINPUT88), .ZN(n578) );
  NAND2_X1 U565 ( .A1(G221), .A2(n479), .ZN(n484) );
  XNOR2_X1 U566 ( .A(G128), .B(G119), .ZN(n480) );
  XNOR2_X1 U567 ( .A(n353), .B(n480), .ZN(n481) );
  XNOR2_X1 U568 ( .A(n484), .B(n483), .ZN(n489) );
  INV_X1 U569 ( .A(KEYINPUT97), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U571 ( .A(n742), .B(n487), .ZN(n488) );
  NAND2_X1 U572 ( .A1(n658), .A2(n490), .ZN(n494) );
  NAND2_X1 U573 ( .A1(G217), .A2(n491), .ZN(n493) );
  INV_X1 U574 ( .A(KEYINPUT25), .ZN(n492) );
  NAND2_X1 U575 ( .A1(n578), .A2(n495), .ZN(n496) );
  OR2_X1 U576 ( .A1(n707), .A2(n702), .ZN(n497) );
  NOR2_X1 U577 ( .A1(n699), .A2(n497), .ZN(n498) );
  AND2_X1 U578 ( .A1(n499), .A2(n498), .ZN(n676) );
  INV_X1 U579 ( .A(KEYINPUT66), .ZN(n533) );
  NOR2_X1 U580 ( .A1(n676), .A2(n533), .ZN(n500) );
  NAND2_X1 U581 ( .A1(n657), .A2(n500), .ZN(n512) );
  NAND2_X1 U582 ( .A1(n502), .A2(n698), .ZN(n515) );
  INV_X1 U583 ( .A(n515), .ZN(n504) );
  INV_X1 U584 ( .A(n572), .ZN(n503) );
  NAND2_X1 U585 ( .A1(n504), .A2(n503), .ZN(n506) );
  INV_X1 U586 ( .A(KEYINPUT33), .ZN(n505) );
  XNOR2_X2 U587 ( .A(n506), .B(n505), .ZN(n732) );
  NAND2_X1 U588 ( .A1(n508), .A2(n387), .ZN(n511) );
  XNOR2_X1 U589 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n509) );
  XNOR2_X1 U590 ( .A(n509), .B(KEYINPUT77), .ZN(n510) );
  XNOR2_X2 U591 ( .A(n511), .B(n510), .ZN(n656) );
  NOR2_X1 U592 ( .A1(n512), .A2(n656), .ZN(n513) );
  NOR2_X1 U593 ( .A1(n513), .A2(n531), .ZN(n530) );
  INV_X1 U594 ( .A(n707), .ZN(n514) );
  NOR2_X1 U595 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U596 ( .A(n516), .B(KEYINPUT102), .ZN(n713) );
  NAND2_X1 U597 ( .A1(n713), .A2(n450), .ZN(n517) );
  XNOR2_X1 U598 ( .A(n517), .B(KEYINPUT31), .ZN(n688) );
  NAND2_X1 U599 ( .A1(n552), .A2(n698), .ZN(n558) );
  NOR2_X1 U600 ( .A1(n518), .A2(n558), .ZN(n519) );
  XOR2_X1 U601 ( .A(KEYINPUT100), .B(n519), .Z(n520) );
  NOR2_X1 U602 ( .A1(n707), .A2(n520), .ZN(n671) );
  NOR2_X1 U603 ( .A1(n688), .A2(n671), .ZN(n521) );
  XNOR2_X1 U604 ( .A(n521), .B(KEYINPUT103), .ZN(n523) );
  OR2_X1 U605 ( .A1(n567), .A2(n566), .ZN(n677) );
  XNOR2_X1 U606 ( .A(n677), .B(KEYINPUT108), .ZN(n604) );
  AND2_X1 U607 ( .A1(n567), .A2(n566), .ZN(n685) );
  INV_X1 U608 ( .A(n685), .ZN(n681) );
  AND2_X1 U609 ( .A1(n604), .A2(n681), .ZN(n721) );
  INV_X1 U610 ( .A(n721), .ZN(n522) );
  NAND2_X1 U611 ( .A1(n523), .A2(n522), .ZN(n528) );
  INV_X1 U612 ( .A(n524), .ZN(n525) );
  NAND2_X1 U613 ( .A1(n525), .A2(n478), .ZN(n526) );
  XNOR2_X1 U614 ( .A(n526), .B(KEYINPUT87), .ZN(n527) );
  NAND2_X1 U615 ( .A1(n527), .A2(n702), .ZN(n669) );
  NAND2_X1 U616 ( .A1(n528), .A2(n669), .ZN(n529) );
  NOR2_X1 U617 ( .A1(n530), .A2(n529), .ZN(n540) );
  INV_X1 U618 ( .A(KEYINPUT44), .ZN(n531) );
  NAND2_X1 U619 ( .A1(n531), .A2(KEYINPUT66), .ZN(n532) );
  OR2_X2 U620 ( .A1(n656), .A2(n532), .ZN(n535) );
  NAND2_X1 U621 ( .A1(n656), .A2(n533), .ZN(n534) );
  NAND2_X1 U622 ( .A1(n535), .A2(n534), .ZN(n538) );
  INV_X1 U623 ( .A(n676), .ZN(n536) );
  AND2_X1 U624 ( .A1(n657), .A2(n536), .ZN(n537) );
  NAND2_X1 U625 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n542) );
  INV_X1 U627 ( .A(KEYINPUT45), .ZN(n541) );
  XNOR2_X2 U628 ( .A(n542), .B(n541), .ZN(n619) );
  NOR2_X1 U629 ( .A1(G900), .A2(n543), .ZN(n544) );
  AND2_X1 U630 ( .A1(n544), .A2(G953), .ZN(n545) );
  NAND2_X1 U631 ( .A1(n703), .A2(n585), .ZN(n547) );
  XOR2_X1 U632 ( .A(KEYINPUT70), .B(n547), .Z(n548) );
  XNOR2_X1 U633 ( .A(n549), .B(KEYINPUT69), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n571), .A2(n559), .ZN(n551) );
  XNOR2_X1 U635 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n550) );
  XNOR2_X1 U636 ( .A(n551), .B(n550), .ZN(n553) );
  NAND2_X1 U637 ( .A1(n553), .A2(n552), .ZN(n583) );
  INV_X1 U638 ( .A(n583), .ZN(n555) );
  NAND2_X1 U639 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X2 U640 ( .A(n556), .B(KEYINPUT78), .ZN(n682) );
  INV_X1 U641 ( .A(KEYINPUT110), .ZN(n557) );
  XNOR2_X1 U642 ( .A(n558), .B(n557), .ZN(n562) );
  AND2_X1 U643 ( .A1(n559), .A2(n356), .ZN(n560) );
  XNOR2_X1 U644 ( .A(n560), .B(KEYINPUT30), .ZN(n561) );
  XNOR2_X1 U645 ( .A(n564), .B(n563), .ZN(n602) );
  INV_X1 U646 ( .A(n585), .ZN(n565) );
  NOR2_X1 U647 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U649 ( .A1(n602), .A2(n569), .ZN(n570) );
  AND2_X1 U650 ( .A1(n388), .A2(n570), .ZN(n680) );
  NOR2_X1 U651 ( .A1(n572), .A2(n681), .ZN(n573) );
  NAND2_X1 U652 ( .A1(n571), .A2(n573), .ZN(n574) );
  XNOR2_X1 U653 ( .A(KEYINPUT109), .B(n574), .ZN(n599) );
  INV_X1 U654 ( .A(n599), .ZN(n575) );
  NOR2_X1 U655 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U656 ( .A(n577), .B(KEYINPUT36), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n691) );
  INV_X1 U658 ( .A(n691), .ZN(n580) );
  NOR2_X1 U659 ( .A1(n581), .A2(n580), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n602), .B(KEYINPUT38), .ZN(n716) );
  NAND2_X1 U661 ( .A1(n716), .A2(n356), .ZN(n720) );
  NOR2_X1 U662 ( .A1(n720), .A2(n719), .ZN(n582) );
  XNOR2_X1 U663 ( .A(n582), .B(KEYINPUT41), .ZN(n731) );
  NOR2_X1 U664 ( .A1(n731), .A2(n583), .ZN(n584) );
  XNOR2_X1 U665 ( .A(n584), .B(KEYINPUT42), .ZN(n752) );
  INV_X1 U666 ( .A(n752), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n606), .A2(n685), .ZN(n589) );
  INV_X1 U668 ( .A(KEYINPUT112), .ZN(n587) );
  XNOR2_X1 U669 ( .A(n587), .B(KEYINPUT40), .ZN(n588) );
  INV_X1 U670 ( .A(n654), .ZN(n590) );
  INV_X1 U671 ( .A(KEYINPUT46), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n598) );
  INV_X1 U673 ( .A(KEYINPUT68), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT48), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n598), .B(n597), .ZN(n608) );
  AND2_X1 U676 ( .A1(n599), .A2(n356), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n600), .A2(n478), .ZN(n601) );
  XNOR2_X1 U678 ( .A(n601), .B(KEYINPUT43), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n631) );
  INV_X1 U680 ( .A(n604), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n618) );
  AND2_X1 U682 ( .A1(n631), .A2(n618), .ZN(n607) );
  XNOR2_X2 U683 ( .A(n610), .B(KEYINPUT83), .ZN(n741) );
  NAND2_X1 U684 ( .A1(n610), .A2(KEYINPUT2), .ZN(n611) );
  INV_X1 U685 ( .A(n619), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n662), .A2(G478), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(n617) );
  INV_X1 U688 ( .A(G952), .ZN(n615) );
  AND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(G63) );
  XNOR2_X1 U690 ( .A(n618), .B(G134), .ZN(G36) );
  NOR2_X1 U691 ( .A1(n619), .A2(G953), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G224), .A2(G953), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n620), .B(KEYINPUT61), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT125), .ZN(n622) );
  NOR2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n629), .B(n628), .ZN(G69) );
  XNOR2_X1 U699 ( .A(n631), .B(G140), .ZN(G42) );
  NAND2_X1 U700 ( .A1(n646), .A2(G475), .ZN(n637) );
  XOR2_X1 U701 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n633) );
  XNOR2_X1 U702 ( .A(KEYINPUT89), .B(KEYINPUT123), .ZN(n632) );
  XOR2_X1 U703 ( .A(n633), .B(n632), .Z(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n639), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U707 ( .A1(n646), .A2(G472), .ZN(n642) );
  XOR2_X1 U708 ( .A(KEYINPUT62), .B(n640), .Z(n641) );
  XNOR2_X1 U709 ( .A(n642), .B(n641), .ZN(n643) );
  NOR2_X2 U710 ( .A1(n643), .A2(n667), .ZN(n645) );
  XNOR2_X1 U711 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(G57) );
  NAND2_X1 U713 ( .A1(n646), .A2(G210), .ZN(n650) );
  XNOR2_X1 U714 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U717 ( .A(KEYINPUT86), .B(KEYINPUT56), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n653), .B(n652), .ZN(G51) );
  XNOR2_X1 U719 ( .A(G131), .B(KEYINPUT127), .ZN(n655) );
  XNOR2_X1 U720 ( .A(n654), .B(n655), .ZN(G33) );
  XOR2_X1 U721 ( .A(n656), .B(G122), .Z(G24) );
  XNOR2_X1 U722 ( .A(n657), .B(G119), .ZN(G21) );
  NAND2_X1 U723 ( .A1(n662), .A2(G217), .ZN(n660) );
  XOR2_X1 U724 ( .A(KEYINPUT124), .B(n658), .Z(n659) );
  XNOR2_X1 U725 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n661), .A2(n667), .ZN(G66) );
  NAND2_X1 U727 ( .A1(n662), .A2(G469), .ZN(n666) );
  XOR2_X1 U728 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n663) );
  XNOR2_X1 U729 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n666), .B(n665), .ZN(n668) );
  NOR2_X1 U731 ( .A1(n668), .A2(n667), .ZN(G54) );
  XNOR2_X1 U732 ( .A(G101), .B(n669), .ZN(G3) );
  NAND2_X1 U733 ( .A1(n671), .A2(n685), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n670), .B(G104), .ZN(G6) );
  XNOR2_X1 U735 ( .A(G107), .B(KEYINPUT114), .ZN(n675) );
  XOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n673) );
  INV_X1 U737 ( .A(n677), .ZN(n687) );
  NAND2_X1 U738 ( .A1(n671), .A2(n687), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U740 ( .A(n675), .B(n674), .ZN(G9) );
  XOR2_X1 U741 ( .A(G110), .B(n676), .Z(G12) );
  NOR2_X1 U742 ( .A1(n682), .A2(n677), .ZN(n679) );
  XNOR2_X1 U743 ( .A(G128), .B(KEYINPUT29), .ZN(n678) );
  XNOR2_X1 U744 ( .A(n679), .B(n678), .ZN(G30) );
  XOR2_X1 U745 ( .A(n344), .B(n680), .Z(G45) );
  NOR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n684) );
  XNOR2_X1 U747 ( .A(G146), .B(KEYINPUT115), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n684), .B(n683), .ZN(G48) );
  NAND2_X1 U749 ( .A1(n688), .A2(n685), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n686), .B(G113), .ZN(G15) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U752 ( .A(n689), .B(G116), .ZN(G18) );
  XOR2_X1 U753 ( .A(G125), .B(KEYINPUT37), .Z(n690) );
  XNOR2_X1 U754 ( .A(n691), .B(n690), .ZN(G27) );
  BUF_X1 U755 ( .A(n692), .Z(n694) );
  XNOR2_X1 U756 ( .A(KEYINPUT82), .B(KEYINPUT2), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U758 ( .A(KEYINPUT81), .B(n695), .Z(n697) );
  NOR2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n739) );
  NOR2_X1 U760 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U761 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n700) );
  XNOR2_X1 U762 ( .A(n701), .B(n700), .ZN(n710) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U764 ( .A(KEYINPUT116), .B(n704), .Z(n705) );
  XNOR2_X1 U765 ( .A(n705), .B(KEYINPUT49), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U767 ( .A(n708), .B(KEYINPUT117), .ZN(n709) );
  NOR2_X1 U768 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U769 ( .A(KEYINPUT119), .B(n711), .Z(n712) );
  NOR2_X1 U770 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U771 ( .A(KEYINPUT51), .B(n714), .Z(n715) );
  NOR2_X1 U772 ( .A1(n731), .A2(n715), .ZN(n726) );
  NOR2_X1 U773 ( .A1(n716), .A2(n356), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n717), .B(KEYINPUT120), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U777 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n724), .A2(n732), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U780 ( .A(KEYINPUT121), .B(n727), .Z(n728) );
  XNOR2_X1 U781 ( .A(n728), .B(KEYINPUT52), .ZN(n729) );
  NOR2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n737) );
  INV_X1 U783 ( .A(n731), .ZN(n734) );
  INV_X1 U784 ( .A(n732), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(n744), .ZN(n736) );
  OR2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U788 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U789 ( .A(n740), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U790 ( .A(n743), .B(n742), .ZN(n747) );
  XNOR2_X1 U791 ( .A(n741), .B(n747), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U793 ( .A(n746), .B(KEYINPUT126), .ZN(n751) );
  XNOR2_X1 U794 ( .A(n747), .B(G227), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U798 ( .A(G137), .B(n752), .Z(G39) );
endmodule

