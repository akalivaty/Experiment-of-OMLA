//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR3_X1   g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n209), .A2(new_n216), .A3(new_n220), .ZN(G361));
  XOR2_X1   g0021(.A(G238), .B(G244), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(G232), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT2), .B(G226), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(G264), .B(G270), .Z(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n225), .B(new_n228), .ZN(G358));
  XOR2_X1   g0029(.A(G87), .B(G97), .Z(new_n230));
  XOR2_X1   g0030(.A(G107), .B(G116), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G58), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G351));
  INV_X1    g0036(.A(KEYINPUT9), .ZN(new_n237));
  OAI21_X1  g0037(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n238));
  INV_X1    g0038(.A(G150), .ZN(new_n239));
  NOR2_X1   g0039(.A1(G20), .A2(G33), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT8), .B(G58), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n218), .A2(G33), .ZN(new_n243));
  OAI221_X1 g0043(.A(new_n238), .B1(new_n239), .B2(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n219), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(KEYINPUT67), .A3(new_n219), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n252), .A2(new_n218), .A3(G1), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n244), .A2(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n249), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT67), .B1(new_n245), .B2(new_n219), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n252), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n257), .A2(G50), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n237), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n254), .A2(new_n237), .A3(new_n262), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G222), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT66), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n269), .A2(KEYINPUT66), .A3(G222), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n270), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n281), .A2(G223), .B1(G77), .B2(new_n280), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n268), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G41), .A2(G45), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT65), .B1(new_n284), .B2(G1), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT65), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n286), .B(new_n260), .C1(G41), .C2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(new_n266), .B2(new_n267), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(G41), .A2(G45), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n292), .A2(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G226), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n283), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n264), .A2(new_n265), .B1(G190), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT69), .ZN(new_n298));
  OAI21_X1  g0098(.A(G200), .B1(new_n283), .B2(new_n295), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT10), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(new_n265), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n301), .B(new_n299), .C1(new_n302), .C2(new_n263), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n254), .A2(new_n262), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n308), .B(new_n309), .C1(G169), .C2(new_n296), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n300), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n253), .A2(new_n246), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(G68), .A3(new_n261), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT70), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G68), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n240), .A2(G50), .B1(G20), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G77), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n243), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n250), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(KEYINPUT11), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n253), .A2(new_n316), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(KEYINPUT11), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n315), .A2(new_n321), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n269), .A2(G232), .A3(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n269), .A2(G226), .A3(new_n270), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n268), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n288), .A2(new_n290), .B1(new_n293), .B2(G238), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(G179), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(KEYINPUT71), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n334), .B2(new_n336), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n337), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n336), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n335), .B1(new_n331), .B2(new_n332), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n342), .B(new_n339), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n325), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n325), .ZN(new_n349));
  OAI21_X1  g0149(.A(G200), .B1(new_n344), .B2(new_n345), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n334), .A2(G190), .A3(new_n336), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n281), .A2(G238), .B1(G107), .B2(new_n280), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n269), .A2(G232), .A3(new_n270), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n330), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n288), .A2(new_n290), .B1(new_n293), .B2(G244), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n338), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n312), .A2(G77), .A3(new_n261), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G77), .B2(new_n259), .ZN(new_n363));
  INV_X1    g0163(.A(new_n242), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n240), .B1(G20), .B2(G77), .ZN(new_n365));
  INV_X1    g0165(.A(G87), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT68), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT68), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n365), .B1(new_n373), .B2(new_n243), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n363), .B1(new_n374), .B2(new_n246), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n358), .A2(new_n307), .A3(new_n359), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n361), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n358), .B2(new_n359), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n375), .B1(new_n360), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n311), .A2(new_n354), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n280), .B2(new_n218), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n386), .B(G20), .C1(new_n277), .C2(new_n279), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G58), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n316), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n390), .B2(new_n201), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n240), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n386), .B1(new_n269), .B2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n316), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n396), .B1(new_n399), .B2(new_n393), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n395), .A2(new_n400), .A3(new_n246), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n248), .A2(new_n259), .A3(new_n249), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n364), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n389), .A2(KEYINPUT8), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n389), .A2(KEYINPUT8), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n261), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n259), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT72), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(KEYINPUT72), .A3(new_n407), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT73), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n395), .A2(new_n400), .A3(new_n246), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  AOI221_X4 g0214(.A(new_n414), .B1(new_n406), .B2(new_n259), .C1(new_n402), .C2(new_n364), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n408), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT73), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n277), .A2(new_n279), .A3(G226), .A4(G1698), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n277), .A2(new_n279), .A3(G223), .A4(new_n270), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n330), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n288), .A2(new_n290), .B1(new_n293), .B2(G232), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G169), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n307), .B2(new_n425), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n412), .A2(new_n418), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT18), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n412), .A2(new_n430), .A3(new_n418), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n379), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n381), .A2(KEYINPUT74), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n381), .A2(KEYINPUT74), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n423), .A2(new_n424), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n413), .A3(new_n416), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n437), .A2(new_n413), .A3(new_n416), .A4(KEYINPUT17), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n429), .A2(new_n431), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n384), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G257), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G1698), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(G250), .B2(G1698), .ZN(new_n447));
  INV_X1    g0247(.A(G294), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n447), .A2(new_n280), .B1(new_n276), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n260), .A2(G45), .ZN(new_n450));
  OR2_X1    g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n449), .A2(new_n330), .B1(new_n290), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  INV_X1    g0256(.A(new_n452), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(G264), .A3(new_n268), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n338), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n453), .A2(new_n290), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G250), .A2(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n445), .B2(G1698), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(new_n269), .B1(G33), .B2(G294), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n460), .B(new_n462), .C1(new_n465), .C2(new_n268), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n307), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT81), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(G169), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n470), .C1(new_n307), .C2(new_n466), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n277), .A2(new_n279), .A3(new_n218), .A4(G87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n269), .A2(new_n475), .A3(new_n218), .A4(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n276), .A2(new_n479), .A3(G20), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n218), .B2(G107), .ZN(new_n482));
  INV_X1    g0282(.A(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(KEYINPUT23), .A3(G20), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n477), .A2(new_n478), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n478), .B1(new_n477), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n246), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n253), .A2(new_n483), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT25), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n260), .A2(G33), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n248), .A2(new_n259), .A3(new_n249), .A4(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n483), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT82), .B1(new_n472), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n488), .A2(new_n494), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(new_n468), .A3(new_n498), .A4(new_n471), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n454), .A2(G190), .A3(new_n460), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n466), .A2(G200), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n488), .A2(new_n500), .A3(new_n494), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n259), .A2(G97), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n241), .A2(new_n318), .ZN(new_n505));
  XNOR2_X1  g0305(.A(G97), .B(G107), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(KEYINPUT6), .A2(G97), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n505), .B1(new_n512), .B2(G20), .ZN(new_n513));
  OAI21_X1  g0313(.A(G107), .B1(new_n385), .B2(new_n387), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n504), .B1(new_n515), .B2(new_n246), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n492), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n459), .A2(G257), .A3(new_n268), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n462), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT76), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n277), .A2(new_n279), .A3(G244), .A4(new_n270), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G250), .A2(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT4), .A2(G244), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(G1698), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n269), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n330), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n519), .A2(new_n462), .A3(KEYINPUT76), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n522), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n516), .A2(new_n518), .B1(new_n338), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n268), .B1(new_n525), .B2(new_n531), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT75), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT77), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n522), .A2(new_n307), .A3(new_n534), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n537), .B(KEYINPUT75), .ZN(new_n543));
  INV_X1    g0343(.A(new_n534), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT76), .B1(new_n519), .B2(new_n462), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n544), .A2(new_n545), .A3(G179), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT77), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n536), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n246), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n277), .A2(new_n279), .A3(new_n218), .A4(G68), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n218), .A2(G33), .A3(G97), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT19), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n366), .A2(new_n517), .A3(new_n483), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n328), .B1(new_n553), .B2(new_n555), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(G20), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n549), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n492), .A2(new_n373), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n259), .B1(new_n369), .B2(new_n372), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G238), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(G1698), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n277), .A3(new_n279), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT78), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n269), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n277), .A2(new_n279), .A3(G244), .A4(G1698), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(KEYINPUT79), .B1(G33), .B2(G116), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT79), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n269), .A2(new_n575), .A3(G244), .A4(G1698), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n330), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n290), .A2(new_n456), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n268), .A2(G250), .A3(new_n450), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n565), .B1(new_n583), .B2(new_n338), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n577), .B2(new_n330), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n307), .ZN(new_n586));
  INV_X1    g0386(.A(new_n564), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n257), .A2(G87), .A3(new_n259), .A4(new_n491), .ZN(new_n588));
  XNOR2_X1  g0388(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n218), .B1(new_n589), .B2(new_n328), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n557), .B1(new_n590), .B2(new_n559), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n587), .B(new_n588), .C1(new_n591), .C2(new_n549), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(G190), .B2(new_n585), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n583), .A2(G200), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n584), .A2(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n218), .A2(G116), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n258), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n312), .A2(G116), .A3(new_n491), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n219), .B2(new_n245), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n526), .B(new_n218), .C1(G33), .C2(new_n517), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT20), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n596), .ZN(new_n602));
  AND4_X1   g0402(.A1(KEYINPUT20), .A2(new_n600), .A3(new_n602), .A4(new_n246), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n597), .B(new_n598), .C1(new_n601), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G303), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n280), .A2(new_n605), .ZN(new_n606));
  MUX2_X1   g0406(.A(G257), .B(G264), .S(G1698), .Z(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n330), .C1(new_n280), .C2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n459), .A2(G270), .A3(new_n268), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n462), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n610), .A3(G169), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n604), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(G200), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n614), .B(new_n615), .C1(new_n435), .C2(new_n610), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n610), .A2(new_n307), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n604), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n604), .A2(new_n610), .A3(KEYINPUT21), .A4(G169), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n613), .A2(new_n616), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n544), .A2(new_n545), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n543), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G200), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n535), .A2(new_n381), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n483), .B1(new_n397), .B2(new_n398), .ZN(new_n625));
  INV_X1    g0425(.A(new_n505), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n510), .B1(new_n506), .B2(new_n507), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n218), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n246), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n504), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n518), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n623), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n548), .A2(new_n595), .A3(new_n620), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n444), .A2(new_n503), .A3(new_n634), .ZN(G372));
  NAND2_X1  g0435(.A1(new_n413), .A2(new_n416), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n430), .A3(new_n427), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n430), .B1(new_n636), .B2(new_n427), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n348), .A2(new_n378), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n440), .A2(new_n441), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n352), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n300), .A2(new_n306), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n310), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n578), .A2(G190), .A3(new_n582), .ZN(new_n650));
  INV_X1    g0450(.A(new_n592), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n650), .B(new_n651), .C1(new_n379), .C2(new_n585), .ZN(new_n652));
  AND4_X1   g0452(.A1(G244), .A2(new_n277), .A3(new_n279), .A4(G1698), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n569), .A2(new_n571), .B1(new_n653), .B2(new_n575), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n268), .B1(new_n654), .B2(new_n574), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n338), .B1(new_n655), .B2(new_n581), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n586), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n649), .B1(new_n548), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n535), .A2(new_n338), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n631), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n543), .A2(new_n546), .A3(KEYINPUT77), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n595), .A2(new_n665), .A3(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n652), .A2(new_n658), .A3(new_n502), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n613), .A2(new_n618), .A3(new_n619), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n469), .B1(new_n307), .B2(new_n466), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n497), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n668), .A2(new_n673), .A3(new_n548), .A4(new_n633), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n658), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n648), .B1(new_n444), .B2(new_n676), .ZN(G369));
  NAND2_X1  g0477(.A1(new_n258), .A2(new_n218), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n679), .A2(new_n680), .A3(G213), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G343), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n620), .B1(new_n614), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n669), .A2(new_n604), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n686), .A2(KEYINPUT83), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(KEYINPUT83), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT84), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT84), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n687), .B2(new_n688), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n503), .B1(new_n497), .B2(new_n684), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n472), .A2(new_n495), .A3(new_n682), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(G330), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n669), .A2(new_n682), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n503), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n672), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n682), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  NOR2_X1   g0502(.A1(new_n559), .A2(G116), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G1), .ZN(new_n704));
  INV_X1    g0504(.A(new_n207), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  MUX2_X1   g0506(.A(new_n704), .B(new_n217), .S(new_n706), .Z(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  NAND2_X1  g0508(.A1(new_n675), .A2(new_n682), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT89), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n379), .B1(new_n543), .B2(new_n621), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n713), .A2(new_n631), .A3(new_n624), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT88), .B1(new_n714), .B2(new_n665), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n496), .A2(new_n499), .A3(new_n670), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT88), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n548), .A2(new_n633), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n715), .A2(new_n716), .A3(new_n668), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n658), .B(KEYINPUT87), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n660), .B2(new_n666), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT29), .A3(new_n682), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n711), .A2(new_n712), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n684), .B1(new_n719), .B2(new_n721), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT86), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n610), .A2(new_n307), .A3(new_n466), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n622), .A2(new_n583), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n535), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n460), .B1(new_n465), .B2(new_n268), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n610), .A2(new_n732), .A3(new_n307), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(new_n733), .A3(KEYINPUT30), .A4(new_n585), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n731), .A2(new_n585), .A3(new_n733), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n730), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT31), .B1(new_n737), .B2(new_n684), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n728), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR3_X1    g0541(.A1(new_n634), .A2(new_n503), .A3(new_n684), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n737), .A2(new_n684), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT86), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n727), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT90), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n727), .A2(KEYINPUT90), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n708), .B1(new_n753), .B2(G1), .ZN(G364));
  NOR2_X1   g0554(.A1(new_n252), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n260), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n706), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n219), .B1(G20), .B2(new_n338), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n762));
  NOR2_X1   g0562(.A1(new_n218), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n381), .A3(new_n379), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT94), .B(G159), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n435), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n218), .A2(new_n307), .A3(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n766), .B1(new_n366), .B2(new_n767), .C1(new_n770), .C2(new_n389), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n763), .A2(new_n381), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G107), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n269), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n381), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n218), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n517), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n771), .A2(new_n775), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n769), .A2(new_n381), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(KEYINPUT92), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(KEYINPUT92), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n218), .A2(new_n307), .A3(new_n379), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT93), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT93), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(new_n768), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n785), .A2(G77), .B1(G50), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n787), .A2(new_n381), .A3(new_n788), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n780), .B(new_n791), .C1(new_n316), .C2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n280), .B1(new_n777), .B2(new_n448), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n770), .A2(new_n796), .B1(new_n797), .B2(new_n781), .ZN(new_n798));
  INV_X1    g0598(.A(new_n767), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n795), .B(new_n798), .C1(G303), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  INV_X1    g0601(.A(G329), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n772), .A2(new_n801), .B1(new_n764), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n790), .A2(G326), .B1(KEYINPUT96), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(KEYINPUT96), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n792), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n800), .A2(new_n804), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n761), .B1(new_n794), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n760), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT91), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n280), .B1(new_n814), .B2(G355), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n207), .B(new_n815), .C1(new_n814), .C2(G355), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n705), .A2(new_n269), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G45), .B2(new_n217), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n235), .A2(new_n455), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n816), .B1(G116), .B2(new_n207), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n759), .B(new_n809), .C1(new_n813), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n689), .ZN(new_n822));
  INV_X1    g0622(.A(new_n812), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n693), .A2(G330), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n759), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n693), .A2(G330), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(G396));
  NOR2_X1   g0628(.A1(new_n760), .A2(new_n810), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n759), .B1(new_n318), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n784), .A2(new_n479), .B1(new_n605), .B2(new_n789), .ZN(new_n831));
  INV_X1    g0631(.A(new_n764), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n269), .B(new_n778), .C1(G311), .C2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n770), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n834), .A2(G294), .B1(G107), .B2(new_n799), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(new_n366), .C2(new_n772), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n831), .B(new_n836), .C1(G283), .C2(new_n792), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n792), .A2(G150), .B1(new_n834), .B2(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n789), .C1(new_n784), .C2(new_n765), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT34), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n269), .B1(new_n764), .B2(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n251), .A2(new_n767), .B1(new_n772), .B2(new_n316), .ZN(new_n844));
  INV_X1    g0644(.A(new_n777), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n843), .B(new_n844), .C1(G58), .C2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n837), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n382), .A2(new_n380), .B1(new_n375), .B2(new_n682), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n378), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n361), .A2(new_n376), .A3(new_n377), .A4(new_n682), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n830), .B1(new_n847), .B2(new_n761), .C1(new_n811), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n851), .B(KEYINPUT97), .ZN(new_n854));
  INV_X1    g0654(.A(new_n658), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n660), .B2(new_n666), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n684), .B1(new_n856), .B2(new_n674), .ZN(new_n857));
  OR3_X1    g0657(.A1(new_n854), .A2(new_n857), .A3(KEYINPUT98), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT98), .B1(new_n854), .B2(new_n857), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(new_n709), .C2(new_n851), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n759), .B1(new_n860), .B2(new_n748), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT99), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n748), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n861), .B2(new_n862), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n853), .B1(new_n863), .B2(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n739), .A2(new_n740), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n742), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n325), .A2(new_n684), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n348), .A2(new_n353), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT14), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n346), .A3(new_n337), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n325), .B(new_n684), .C1(new_n873), .C2(new_n352), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n851), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n395), .A2(new_n400), .A3(new_n250), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n681), .B1(new_n878), .B2(new_n411), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n643), .B1(KEYINPUT18), .B2(new_n428), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n880), .B2(new_n431), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n412), .A2(new_n418), .A3(new_n681), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n438), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n428), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n427), .B1(new_n878), .B2(new_n411), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n879), .A2(new_n886), .A3(new_n438), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n877), .B1(new_n881), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT100), .ZN(new_n892));
  INV_X1    g0692(.A(new_n879), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n443), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n892), .B1(new_n891), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n876), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  AOI221_X4 g0701(.A(new_n877), .B1(new_n885), .B2(new_n888), .C1(new_n443), .C2(new_n893), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n417), .B1(new_n413), .B2(new_n416), .ZN(new_n904));
  INV_X1    g0704(.A(new_n681), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT102), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n440), .A2(new_n907), .A3(new_n441), .ZN(new_n908));
  INV_X1    g0708(.A(new_n639), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n637), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n907), .B1(new_n440), .B2(new_n441), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n636), .A2(new_n427), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n438), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n885), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT38), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n901), .B1(new_n902), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n643), .A2(KEYINPUT102), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n640), .A3(new_n908), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n920), .A2(new_n906), .B1(new_n915), .B2(new_n885), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n895), .B(KEYINPUT103), .C1(KEYINPUT38), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n745), .A2(new_n738), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n634), .A2(new_n503), .A3(new_n684), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n875), .B(KEYINPUT40), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n918), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n900), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n444), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n868), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n930), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(G330), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT104), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n902), .B2(new_n917), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n873), .A2(new_n325), .A3(new_n682), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT101), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT101), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n873), .A2(new_n941), .A3(new_n325), .A4(new_n682), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n894), .B2(new_n889), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT100), .B1(new_n902), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n870), .A2(new_n874), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n684), .B(new_n851), .C1(new_n856), .C2(new_n674), .ZN(new_n950));
  INV_X1    g0750(.A(new_n850), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n641), .A2(new_n905), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n944), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n444), .B1(new_n724), .B2(new_n726), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n647), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n934), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n934), .A2(new_n959), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n260), .C2(new_n755), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n219), .A2(new_n218), .A3(new_n479), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  OAI21_X1  g0767(.A(G77), .B1(new_n389), .B2(new_n316), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n217), .A2(new_n968), .B1(G50), .B2(new_n316), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n252), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT105), .ZN(G367));
  AOI21_X1  g0772(.A(new_n696), .B1(new_n669), .B2(new_n682), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(new_n699), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n825), .B(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n631), .A2(new_n684), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n715), .A2(new_n718), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n665), .A2(new_n684), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n701), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT45), .Z(new_n982));
  NOR2_X1   g0782(.A1(new_n701), .A2(new_n980), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT44), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n697), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(new_n984), .ZN(new_n986));
  INV_X1    g0786(.A(new_n697), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n976), .A2(new_n753), .A3(new_n985), .A4(new_n988), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n989), .A2(new_n753), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n706), .B(KEYINPUT41), .Z(new_n991));
  OAI21_X1  g0791(.A(new_n756), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n980), .A2(new_n699), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT106), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n496), .A2(new_n499), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n978), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n684), .B1(new_n997), .B2(new_n548), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n994), .B2(KEYINPUT42), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n595), .B1(new_n651), .B2(new_n682), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n855), .A2(new_n592), .A3(new_n684), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1003), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT43), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1005), .A2(new_n1008), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n987), .A2(new_n980), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1012), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1007), .A2(new_n812), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n817), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n813), .B1(new_n207), .B2(new_n373), .C1(new_n1017), .C2(new_n228), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n758), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT107), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n280), .B1(new_n764), .B2(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n770), .A2(new_n605), .B1(new_n517), .B2(new_n772), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G107), .C2(new_n845), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n767), .A2(new_n479), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT46), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT108), .Z(new_n1027));
  OAI211_X1 g0827(.A(new_n1024), .B(new_n1027), .C1(KEYINPUT46), .C2(new_n1025), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G311), .A2(new_n790), .B1(new_n792), .B2(G294), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n801), .B2(new_n784), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n834), .A2(G150), .B1(G68), .B2(new_n845), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n280), .B1(new_n773), .B2(G77), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n784), .C2(new_n251), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n764), .A2(new_n839), .B1(new_n767), .B2(new_n389), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT109), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n790), .A2(G143), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n765), .C2(new_n793), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1028), .A2(new_n1030), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT47), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n761), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1020), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n992), .A2(new_n1015), .B1(new_n1016), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(G387));
  INV_X1    g0844(.A(new_n706), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n976), .B2(new_n753), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n975), .A2(new_n751), .A3(new_n752), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n225), .A2(new_n455), .A3(new_n269), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(G50), .B2(new_n242), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n455), .C1(new_n316), .C2(new_n318), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1050), .A2(G50), .A3(new_n242), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n280), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n703), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n705), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n813), .B1(new_n207), .B2(new_n483), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n781), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n792), .A2(new_n364), .B1(new_n1058), .B2(G68), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT112), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n373), .A2(new_n777), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G50), .B2(new_n834), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT111), .ZN(new_n1063));
  INV_X1    g0863(.A(G159), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n789), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n280), .B1(new_n832), .B2(G150), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n799), .A2(G77), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n517), .C2(new_n772), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n790), .A2(G322), .B1(new_n834), .B2(G317), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n605), .B2(new_n784), .C1(new_n797), .C2(new_n793), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n845), .A2(G283), .B1(new_n799), .B2(G294), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT49), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n772), .A2(new_n479), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n269), .B(new_n1078), .C1(G326), .C2(new_n832), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1069), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n758), .B1(new_n1056), .B2(new_n1057), .C1(new_n1080), .C2(new_n761), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n696), .C2(new_n823), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n975), .B2(new_n756), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1048), .A2(new_n1087), .ZN(G393));
  NAND3_X1  g0888(.A1(new_n988), .A2(KEYINPUT114), .A3(new_n985), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n986), .A2(new_n1090), .A3(new_n987), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n757), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n817), .A2(new_n232), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n813), .B1(new_n207), .B2(new_n517), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n758), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n793), .A2(new_n251), .B1(new_n777), .B2(new_n318), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n785), .B2(new_n364), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n280), .B1(new_n832), .B2(G143), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n316), .B2(new_n767), .C1(new_n366), .C2(new_n772), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT116), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n789), .A2(new_n239), .B1(new_n770), .B2(new_n1064), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1103));
  XNOR2_X1  g0903(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1098), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n789), .A2(new_n1021), .B1(new_n770), .B2(new_n797), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT52), .Z(new_n1107));
  OAI22_X1  g0907(.A1(new_n781), .A2(new_n448), .B1(new_n767), .B2(new_n801), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n774), .B(new_n280), .C1(new_n796), .C2(new_n764), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(G116), .C2(new_n845), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n605), .B2(new_n793), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1105), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1096), .B1(new_n1112), .B2(new_n760), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n980), .B2(new_n823), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n989), .A2(new_n706), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n975), .B1(new_n751), .B2(new_n752), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n1092), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1093), .B(new_n1114), .C1(new_n1115), .C2(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n951), .B1(new_n857), .B2(new_n852), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n949), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n943), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n938), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n849), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n684), .B(new_n1123), .C1(new_n719), .C2(new_n721), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n949), .B1(new_n1124), .B2(new_n951), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT117), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n940), .A2(new_n1126), .A3(new_n942), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n940), .B2(new_n942), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1125), .A2(new_n918), .A3(new_n922), .A4(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n747), .A2(G330), .A3(new_n852), .A4(new_n949), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1122), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n918), .A2(new_n922), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n722), .A2(new_n682), .A3(new_n849), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n850), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1136), .B2(new_n949), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1133), .A2(new_n1137), .B1(new_n938), .B2(new_n1121), .ZN(new_n1138));
  INV_X1    g0938(.A(G330), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n742), .B2(new_n867), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n875), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1132), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n938), .A2(new_n810), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n829), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n758), .B1(new_n364), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G283), .A2(new_n790), .B1(new_n792), .B2(G107), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n517), .B2(new_n784), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n280), .B1(new_n764), .B2(new_n448), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G87), .B2(new_n799), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n845), .A2(G77), .B1(new_n773), .B2(G68), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n479), .C2(new_n770), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n767), .A2(new_n239), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT53), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1154), .B1(new_n1155), .B2(new_n789), .C1(new_n784), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n792), .A2(G137), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n834), .A2(G132), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n280), .B1(new_n832), .B2(G125), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n845), .A2(G159), .B1(new_n773), .B2(G50), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1148), .A2(new_n1152), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1146), .B1(new_n1163), .B2(new_n760), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1143), .A2(new_n757), .B1(new_n1144), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1140), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n444), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n957), .A2(new_n647), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n868), .A2(G330), .A3(new_n854), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1120), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n951), .B1(new_n725), .B2(new_n849), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n1131), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n747), .A2(G330), .A3(new_n852), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1173), .A2(new_n1120), .B1(new_n875), .B2(new_n1140), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1174), .B2(new_n1119), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1045), .B1(new_n1142), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1141), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1129), .B1(new_n1171), .B2(new_n1120), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n918), .A2(new_n922), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n943), .A2(new_n952), .B1(new_n936), .B2(new_n937), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1178), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1183), .A2(new_n1132), .A3(new_n1168), .A4(new_n1175), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1177), .A2(KEYINPUT118), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT118), .B1(new_n1177), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1165), .B1(new_n1185), .B2(new_n1186), .ZN(G378));
  NAND2_X1  g0987(.A1(new_n1173), .A2(new_n1120), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1119), .B1(new_n1188), .B2(new_n1141), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1170), .A2(new_n1171), .A3(new_n1131), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1168), .B1(new_n1142), .B2(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n944), .A2(new_n954), .A3(new_n955), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n311), .A2(new_n309), .A3(new_n681), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n309), .A2(new_n681), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n300), .A2(new_n306), .A3(new_n310), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1194), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n927), .A2(G330), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n900), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT40), .B1(new_n948), .B2(new_n876), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n927), .A2(G330), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT121), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1201), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1198), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1200), .A2(KEYINPUT121), .A3(new_n1201), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1205), .A2(new_n1206), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1193), .B1(new_n1204), .B2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1201), .B(new_n1200), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1203), .A2(new_n900), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1217), .A3(new_n956), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1192), .A2(new_n1214), .A3(KEYINPUT57), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT122), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1192), .A2(new_n1214), .A3(new_n1218), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1184), .B2(new_n1168), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1225), .A2(KEYINPUT122), .A3(new_n1214), .A4(new_n1218), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1221), .A2(new_n1224), .A3(new_n1226), .A4(new_n706), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1212), .A2(new_n810), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n758), .B1(G50), .B2(new_n1145), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1067), .B1(new_n389), .B2(new_n772), .C1(new_n770), .C2(new_n483), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n373), .A2(new_n781), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n269), .A2(G41), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n764), .B2(new_n801), .C1(new_n316), .C2(new_n777), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n517), .B2(new_n793), .C1(new_n479), .C2(new_n789), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT58), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n251), .B1(G33), .B2(G41), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n1236), .A2(new_n1237), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1237), .B2(new_n1236), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G137), .A2(new_n1058), .B1(new_n845), .B2(G150), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n793), .B2(new_n842), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n770), .A2(new_n1155), .B1(new_n767), .B2(new_n1156), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT119), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(G125), .C2(new_n790), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT59), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT120), .ZN(new_n1247));
  AOI211_X1 g1047(.A(G33), .B(G41), .C1(new_n832), .C2(G124), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n765), .C2(new_n772), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1246), .A2(KEYINPUT120), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1240), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1230), .B1(new_n1251), .B2(new_n760), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1228), .A2(new_n757), .B1(new_n1229), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1227), .A2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n1120), .A2(new_n810), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n758), .B1(G68), .B2(new_n1145), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT124), .Z(new_n1257));
  OAI22_X1  g1057(.A1(new_n793), .A2(new_n479), .B1(new_n448), .B2(new_n789), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G107), .B2(new_n785), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n280), .B1(new_n772), .B2(new_n318), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT125), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n770), .A2(new_n801), .B1(new_n605), .B2(new_n764), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1061), .B(new_n1262), .C1(G97), .C2(new_n799), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1259), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n834), .A2(G137), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n842), .B2(new_n789), .C1(new_n793), .C2(new_n1156), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n781), .A2(new_n239), .B1(new_n767), .B2(new_n1064), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n269), .B1(new_n764), .B2(new_n1155), .C1(new_n389), .C2(new_n772), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(G50), .C2(new_n845), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1264), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1257), .B1(new_n1274), .B2(new_n760), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1175), .A2(new_n757), .B1(new_n1255), .B2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n991), .B(KEYINPUT123), .Z(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1176), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1276), .B1(new_n1279), .B2(new_n1280), .ZN(G381));
  XOR2_X1   g1081(.A(G375), .B(KEYINPUT127), .Z(new_n1282));
  NOR3_X1   g1082(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1283));
  INV_X1    g1083(.A(G396), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1048), .A2(new_n1284), .A3(new_n1087), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1177), .A2(new_n1184), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1165), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1282), .A2(new_n1043), .A3(new_n1283), .A4(new_n1288), .ZN(G407));
  INV_X1    g1089(.A(new_n1287), .ZN(new_n1290));
  INV_X1    g1090(.A(G343), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(G213), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1282), .A2(new_n1290), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(G407), .A2(G213), .A3(new_n1294), .ZN(G409));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1284), .B1(new_n1048), .B2(new_n1087), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1285), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1297), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(G390), .A3(new_n1285), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1299), .A2(new_n1043), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1043), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1227), .A2(G378), .A3(new_n1253), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1228), .A2(new_n1192), .A3(new_n1278), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1253), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1290), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1292), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1167), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n648), .B(new_n1311), .C1(new_n727), .C2(new_n444), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1191), .A2(KEYINPUT60), .A3(new_n1312), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1313), .A2(new_n706), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1314), .B1(new_n1280), .B2(new_n1315), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1316), .A2(G384), .A3(new_n1276), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1316), .B2(new_n1276), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G2897), .B(new_n1293), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1318), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1316), .A2(G384), .A3(new_n1276), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1293), .A2(G2897), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1310), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1326), .B1(new_n1310), .B2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1293), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1327), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1304), .A2(new_n1325), .A3(new_n1329), .A4(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1330), .A2(new_n1333), .A3(new_n1327), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1335), .B1(new_n1330), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1330), .B2(new_n1327), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1334), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1332), .B1(new_n1339), .B2(new_n1304), .ZN(G405));
  NAND2_X1  g1140(.A1(G375), .A2(new_n1290), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1305), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1327), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1328), .A3(new_n1305), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1345), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1304), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(G402));
endmodule


