//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n608, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n468), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n466), .A2(new_n468), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n482), .A3(new_n464), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n477), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(new_n482), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n464), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(G124), .B2(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n466), .A2(new_n468), .A3(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n490), .B1(G114), .B2(G2104), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n491), .A2(new_n464), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n466), .A2(new_n468), .A3(new_n495), .A4(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n492), .A2(new_n493), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n481), .B2(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n496), .A2(new_n497), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n464), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n499), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT72), .A3(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(G88), .B1(G50), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(G166));
  NAND2_X1  g102(.A1(new_n523), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n522), .A2(new_n535), .B1(new_n524), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT74), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n540), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n522), .A2(new_n546), .B1(new_n524), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n523), .A2(G91), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT75), .Z(new_n558));
  XNOR2_X1  g133(.A(new_n516), .B(KEYINPUT76), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n562), .A2(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n558), .A2(new_n566), .ZN(G299));
  XOR2_X1   g142(.A(new_n533), .B(KEYINPUT77), .Z(G286));
  NAND2_X1  g143(.A1(new_n520), .A2(new_n526), .ZN(G303));
  NAND2_X1  g144(.A1(new_n523), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n525), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n523), .A2(G86), .B1(G48), .B2(new_n525), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n516), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT78), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n577), .A2(new_n580), .A3(G651), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n540), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n522), .A2(new_n585), .B1(new_n524), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n524), .B(KEYINPUT79), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G54), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n512), .A2(G92), .A3(new_n521), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n559), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n592), .B(new_n594), .C1(new_n540), .C2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G286), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G280));
  NOR2_X1   g182(.A1(new_n599), .A2(G559), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G860), .B2(new_n600), .ZN(G148));
  NAND2_X1  g184(.A1(new_n549), .A2(new_n603), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n608), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n487), .A2(G123), .ZN(new_n613));
  INV_X1    g188(.A(new_n483), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G135), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n618), .B(new_n619), .C1(G111), .C2(new_n464), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n613), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT82), .B(G2096), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2100), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT84), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  AND2_X1   g217(.A1(new_n642), .A2(G14), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI211_X1 g225(.A(KEYINPUT17), .B(new_n645), .C1(new_n648), .C2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n647), .B2(new_n649), .ZN(new_n653));
  OAI221_X1 g228(.A(new_n651), .B1(new_n647), .B2(new_n649), .C1(new_n653), .C2(new_n645), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n647), .A2(new_n644), .A3(new_n649), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2096), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT86), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n661), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1986), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n674), .B(new_n678), .Z(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n680), .A2(G26), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n487), .A2(G128), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n614), .A2(G140), .ZN(new_n683));
  OAI21_X1  g258(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n464), .A2(G116), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n681), .B1(new_n686), .B2(G29), .ZN(new_n687));
  MUX2_X1   g262(.A(new_n681), .B(new_n687), .S(KEYINPUT28), .Z(new_n688));
  INV_X1    g263(.A(G2067), .ZN(new_n689));
  INV_X1    g264(.A(G27), .ZN(new_n690));
  OAI21_X1  g265(.A(KEYINPUT95), .B1(new_n690), .B2(G29), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n690), .A2(KEYINPUT95), .A3(G29), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n691), .B(new_n692), .C1(G164), .C2(new_n680), .ZN(new_n693));
  OAI22_X1  g268(.A1(new_n688), .A2(new_n689), .B1(G2078), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT97), .ZN(new_n695));
  NAND2_X1  g270(.A1(G162), .A2(G29), .ZN(new_n696));
  OR2_X1    g271(.A1(G29), .A2(G35), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n695), .B1(new_n703), .B2(G2090), .ZN(new_n704));
  INV_X1    g279(.A(G2090), .ZN(new_n705));
  OAI211_X1 g280(.A(KEYINPUT97), .B(new_n705), .C1(new_n701), .C2(new_n702), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n694), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(G299), .A2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n709), .A2(KEYINPUT23), .A3(G20), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT23), .ZN(new_n711));
  INV_X1    g286(.A(G20), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n708), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1956), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n550), .A2(new_n709), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n709), .B2(G19), .ZN(new_n717));
  INV_X1    g292(.A(G1341), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(KEYINPUT24), .A2(G34), .ZN(new_n720));
  NAND2_X1  g295(.A1(KEYINPUT24), .A2(G34), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n680), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G160), .B2(new_n680), .ZN(new_n723));
  OAI22_X1  g298(.A1(new_n717), .A2(new_n718), .B1(G2084), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n715), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n688), .A2(new_n689), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n707), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT90), .B1(G4), .B2(G16), .ZN(new_n728));
  OR3_X1    g303(.A1(KEYINPUT90), .A2(G4), .A3(G16), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(new_n599), .C2(new_n709), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1348), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  OR2_X1    g307(.A1(KEYINPUT30), .A2(G28), .ZN(new_n733));
  NAND2_X1  g308(.A1(KEYINPUT30), .A2(G28), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n621), .A2(new_n680), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n735), .B(new_n736), .C1(G2084), .C2(new_n723), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n731), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT25), .Z(new_n740));
  INV_X1    g315(.A(G139), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n483), .B2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT91), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  INV_X1    g321(.A(G127), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n478), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G2105), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G29), .B2(G33), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT92), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n753), .A2(new_n754), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n703), .A2(G2090), .ZN(new_n758));
  NAND2_X1  g333(.A1(G171), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G5), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n693), .A2(G2078), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n757), .A2(new_n758), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n727), .A2(new_n738), .A3(new_n756), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G21), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G168), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT94), .B(G1966), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n709), .A2(G22), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G166), .B2(new_n709), .ZN(new_n771));
  MUX2_X1   g346(.A(new_n770), .B(new_n771), .S(KEYINPUT87), .Z(new_n772));
  INV_X1    g347(.A(G1971), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G23), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT33), .B(G1976), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n709), .A2(G6), .ZN(new_n780));
  INV_X1    g355(.A(G305), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n709), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT32), .B(G1981), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n774), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n709), .A2(G24), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n588), .B2(new_n709), .ZN(new_n788));
  INV_X1    g363(.A(G1986), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n774), .A2(new_n791), .A3(new_n779), .A4(new_n784), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n487), .A2(G119), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n614), .A2(G131), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n464), .A2(G107), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G25), .B(new_n797), .S(G29), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT35), .B(G1991), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n798), .B(new_n799), .Z(new_n800));
  NAND4_X1  g375(.A1(new_n786), .A2(new_n790), .A3(new_n792), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT89), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n801), .A2(new_n804), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n765), .B(new_n769), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n614), .A2(G141), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n811));
  NAND3_X1  g386(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT26), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n811), .B(new_n813), .C1(new_n487), .C2(G129), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G29), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G29), .B2(G32), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT27), .B(G1996), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n760), .A2(new_n761), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n807), .A2(new_n820), .A3(new_n821), .ZN(G311));
  INV_X1    g397(.A(new_n807), .ZN(new_n823));
  INV_X1    g398(.A(new_n820), .ZN(new_n824));
  INV_X1    g399(.A(new_n821), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(G150));
  AOI22_X1  g401(.A1(new_n523), .A2(G93), .B1(G55), .B2(new_n525), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n540), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n600), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n829), .B(new_n549), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT39), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n832), .B1(new_n837), .B2(G860), .ZN(G145));
  XNOR2_X1  g413(.A(new_n621), .B(G160), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G162), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n797), .B(new_n625), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G118), .B2(new_n464), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT99), .B1(new_n614), .B2(G142), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n614), .A2(KEYINPUT99), .A3(G142), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n487), .A2(G130), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n850));
  OAI221_X1 g425(.A(new_n845), .B1(new_n846), .B2(new_n847), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n842), .B(new_n851), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n816), .A2(new_n750), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n751), .A2(new_n815), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n494), .A2(new_n498), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n686), .B(new_n855), .Z(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n853), .B2(new_n854), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n852), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n853), .A2(new_n854), .ZN(new_n861));
  INV_X1    g436(.A(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n842), .B(new_n851), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n857), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n841), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n865), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n840), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n863), .A2(new_n857), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n870), .B2(new_n852), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n866), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT101), .B(G37), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(KEYINPUT103), .A3(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT103), .B1(new_n873), .B2(new_n875), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT102), .B1(new_n860), .B2(new_n865), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n883), .A2(new_n871), .A3(new_n840), .ZN(new_n884));
  NOR4_X1   g459(.A1(new_n884), .A2(new_n877), .A3(new_n874), .A4(new_n866), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT40), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n886), .ZN(G395));
  NAND2_X1  g462(.A1(new_n829), .A2(new_n603), .ZN(new_n888));
  INV_X1    g463(.A(new_n835), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n608), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G299), .B(new_n596), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n596), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G299), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n892), .B1(new_n898), .B2(new_n890), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n776), .B(G303), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G305), .ZN(new_n901));
  XNOR2_X1  g476(.A(G303), .B(G288), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n781), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n588), .B(KEYINPUT104), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n904), .B1(new_n901), .B2(new_n903), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n906), .A2(KEYINPUT42), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  INV_X1    g485(.A(new_n907), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT105), .A3(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n908), .B1(new_n913), .B2(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n899), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n888), .B1(new_n915), .B2(new_n603), .ZN(G295));
  OAI21_X1  g491(.A(new_n888), .B1(new_n915), .B2(new_n603), .ZN(G331));
  INV_X1    g492(.A(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(G171), .A2(G286), .ZN(new_n919));
  NAND2_X1  g494(.A1(G301), .A2(G168), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n835), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n889), .A3(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n896), .B2(new_n897), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n891), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n918), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n922), .A2(new_n923), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n898), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n913), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n927), .A2(new_n930), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n896), .A2(KEYINPUT107), .A3(new_n897), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n895), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n936), .A2(new_n924), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n918), .B1(new_n938), .B2(new_n926), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n874), .B1(new_n929), .B2(new_n913), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n933), .A2(new_n934), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n935), .A2(KEYINPUT44), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n927), .A2(new_n932), .A3(new_n930), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n939), .A2(new_n940), .A3(new_n931), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n944), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(new_n471), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n472), .A2(new_n473), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n464), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n954), .A3(G40), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n494), .B2(new_n498), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n960), .A2(G1996), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n816), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n686), .B(new_n689), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT111), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n816), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n960), .A2(new_n964), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n969), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n967), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n797), .B(new_n799), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n588), .B(new_n789), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n499), .A2(new_n961), .A3(new_n506), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n981), .A2(KEYINPUT50), .B1(new_n957), .B2(new_n958), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n961), .B(new_n984), .C1(new_n494), .C2(new_n498), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT113), .ZN(new_n986));
  AOI21_X1  g561(.A(G1961), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n963), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n502), .B2(new_n505), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n959), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n991), .A2(G2078), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n499), .A2(new_n506), .A3(KEYINPUT45), .A4(new_n961), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n957), .A2(new_n958), .B1(new_n962), .B2(new_n963), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n959), .A2(new_n997), .A3(new_n964), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n993), .A2(G2078), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n994), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1966), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n998), .B2(new_n999), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT117), .B(G2084), .Z(new_n1006));
  NAND3_X1  g581(.A1(new_n982), .A2(new_n986), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(G168), .A3(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(KEYINPUT125), .A2(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1008), .A2(KEYINPUT51), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(G8), .A3(new_n533), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(KEYINPUT124), .A3(new_n533), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1012), .A2(new_n1013), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT62), .ZN(new_n1022));
  OAI211_X1 g597(.A(G171), .B(new_n1003), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n982), .A2(new_n986), .A3(new_n705), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n982), .A2(new_n986), .A3(KEYINPUT114), .A4(new_n705), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n991), .A2(new_n773), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT55), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1029), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n499), .A2(new_n506), .A3(new_n1034), .A4(new_n961), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n962), .A2(new_n983), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(new_n959), .A3(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n773), .A2(new_n991), .B1(new_n1037), .B2(new_n705), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1031), .B1(new_n1038), .B2(new_n1018), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n1040));
  INV_X1    g615(.A(G40), .ZN(new_n1041));
  NOR4_X1   g616(.A1(new_n471), .A2(new_n474), .A3(new_n956), .A4(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n989), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n570), .A2(new_n571), .A3(G1976), .A4(new_n572), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(G8), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n776), .A2(G1976), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1043), .A2(G8), .A3(new_n1045), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT115), .B1(new_n1050), .B2(new_n1044), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1048), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1044), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1049), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G305), .A2(G1981), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n781), .A2(new_n676), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(new_n1056), .A3(KEYINPUT49), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1043), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1018), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1039), .A2(new_n1054), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT126), .B1(new_n1033), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1029), .A2(G8), .A3(new_n1032), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1050), .A2(KEYINPUT115), .A3(new_n1044), .A4(new_n1052), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1043), .A2(G8), .A3(new_n1045), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1047), .B1(new_n1069), .B2(KEYINPUT52), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1064), .B(new_n1068), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT126), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1067), .A2(new_n1073), .A3(new_n1074), .A4(new_n1039), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n1022), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT127), .B1(new_n1023), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1021), .A2(new_n1022), .B1(new_n1066), .B2(new_n1075), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT127), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1019), .A2(KEYINPUT124), .A3(new_n533), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT124), .B1(new_n1019), .B2(new_n533), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1008), .A2(KEYINPUT51), .A3(new_n1009), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT51), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1084), .A2(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G301), .B1(new_n1088), .B2(KEYINPUT62), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1082), .A2(new_n1083), .A3(new_n1003), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1018), .B(G286), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1067), .A2(new_n1073), .A3(new_n1039), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT118), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1019), .A2(new_n605), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1029), .A2(G8), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1031), .A2(KEYINPUT119), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT63), .A4(new_n1073), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1093), .A2(new_n1103), .A3(new_n1094), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1096), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1976), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1064), .A2(new_n1106), .A3(new_n776), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1060), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1033), .A2(new_n1073), .B1(new_n1063), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT120), .B1(new_n565), .B2(new_n564), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT121), .B1(new_n1110), .B2(KEYINPUT57), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1110), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n1113));
  OAI21_X1  g688(.A(G299), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(new_n566), .A3(new_n558), .A4(new_n1111), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT123), .ZN(new_n1118));
  INV_X1    g693(.A(new_n991), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1037), .A2(G1956), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1114), .A2(new_n1124), .A3(new_n1116), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1118), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n982), .B2(new_n986), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1062), .A2(new_n689), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT122), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1117), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n893), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1126), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n596), .B1(new_n1134), .B2(KEYINPUT60), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1139), .B(new_n893), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1138), .A2(new_n1140), .B1(KEYINPUT60), .B2(new_n1134), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1126), .A2(KEYINPUT61), .A3(new_n1135), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1135), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1117), .B1(new_n1122), .B2(new_n1121), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT58), .B(G1341), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n991), .A2(G1996), .B1(new_n1062), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n550), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT59), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1142), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1137), .B1(new_n1141), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(G301), .B(KEYINPUT54), .Z(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n964), .A2(new_n990), .A3(new_n1001), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n955), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1003), .A2(new_n1154), .B1(new_n1157), .B2(new_n994), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1076), .A2(new_n1088), .A3(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1105), .B(new_n1109), .C1(new_n1152), .C2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n980), .B1(new_n1091), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n971), .A2(new_n789), .A3(new_n588), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT48), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n977), .A2(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n797), .A2(new_n799), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n975), .A2(new_n1165), .B1(G2067), .B2(new_n686), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n971), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT46), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n966), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n966), .A2(new_n1168), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n972), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT47), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1164), .A2(new_n1167), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1161), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g749(.A(G229), .ZN(new_n1176));
  NAND3_X1  g750(.A1(new_n948), .A2(G319), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g751(.A1(G401), .A2(G227), .ZN(new_n1178));
  OAI21_X1  g752(.A(new_n1178), .B1(new_n882), .B2(new_n885), .ZN(new_n1179));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1179), .ZN(G308));
  NAND2_X1  g754(.A1(new_n878), .A2(new_n880), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n462), .B1(new_n946), .B2(new_n947), .ZN(new_n1182));
  NAND4_X1  g756(.A1(new_n1181), .A2(new_n1176), .A3(new_n1182), .A4(new_n1178), .ZN(G225));
endmodule


