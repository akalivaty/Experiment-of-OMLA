

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n390), .B(n312), .ZN(n313) );
  XNOR2_X1 U322 ( .A(n470), .B(KEYINPUT37), .ZN(n471) );
  INV_X1 U323 ( .A(KEYINPUT104), .ZN(n470) );
  XOR2_X1 U324 ( .A(G36GAT), .B(G218GAT), .Z(n395) );
  XNOR2_X1 U325 ( .A(n319), .B(n318), .ZN(n323) );
  XNOR2_X1 U326 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U327 ( .A(n485), .B(KEYINPUT125), .ZN(n577) );
  INV_X1 U328 ( .A(n577), .ZN(n582) );
  XNOR2_X1 U329 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n289) );
  AND2_X1 U330 ( .A1(G226GAT), .A2(G233GAT), .ZN(n290) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U332 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n401) );
  XNOR2_X1 U333 ( .A(n405), .B(n311), .ZN(n312) );
  XNOR2_X1 U334 ( .A(n374), .B(n291), .ZN(n375) );
  XNOR2_X1 U335 ( .A(n395), .B(n290), .ZN(n396) );
  XNOR2_X1 U336 ( .A(n376), .B(n375), .ZN(n381) );
  XNOR2_X1 U337 ( .A(n397), .B(n396), .ZN(n399) );
  XNOR2_X1 U338 ( .A(n472), .B(n471), .ZN(n528) );
  INV_X1 U339 ( .A(G218GAT), .ZN(n487) );
  XNOR2_X1 U340 ( .A(n340), .B(n339), .ZN(n572) );
  INV_X1 U341 ( .A(G29GAT), .ZN(n474) );
  XNOR2_X1 U342 ( .A(n487), .B(KEYINPUT62), .ZN(n488) );
  XNOR2_X1 U343 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U344 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U345 ( .A(n489), .B(n488), .ZN(G1355GAT) );
  XNOR2_X1 U346 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n477), .B(n476), .ZN(G1328GAT) );
  INV_X1 U348 ( .A(KEYINPUT121), .ZN(n446) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(G176GAT), .ZN(n298) );
  XOR2_X1 U350 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n293) );
  XNOR2_X1 U351 ( .A(KEYINPUT18), .B(KEYINPUT83), .ZN(n292) );
  XNOR2_X1 U352 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U353 ( .A(n294), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U354 ( .A(G190GAT), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U356 ( .A(n298), .B(n297), .Z(n398) );
  XOR2_X1 U357 ( .A(G43GAT), .B(G134GAT), .Z(n367) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G71GAT), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n299), .B(G120GAT), .ZN(n321) );
  XOR2_X1 U360 ( .A(n367), .B(n321), .Z(n301) );
  NAND2_X1 U361 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U362 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U363 ( .A(KEYINPUT82), .B(KEYINPUT85), .Z(n303) );
  XNOR2_X1 U364 ( .A(KEYINPUT20), .B(KEYINPUT86), .ZN(n302) );
  XNOR2_X1 U365 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U366 ( .A(n305), .B(n304), .Z(n307) );
  XOR2_X1 U367 ( .A(G113GAT), .B(G15GAT), .Z(n335) );
  XOR2_X1 U368 ( .A(KEYINPUT0), .B(G127GAT), .Z(n406) );
  XNOR2_X1 U369 ( .A(n335), .B(n406), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U371 ( .A(n398), .B(n308), .ZN(n541) );
  INV_X1 U372 ( .A(n541), .ZN(n509) );
  XOR2_X1 U373 ( .A(G64GAT), .B(KEYINPUT73), .Z(n310) );
  XNOR2_X1 U374 ( .A(G204GAT), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n390) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G57GAT), .Z(n405) );
  NAND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XOR2_X1 U378 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n344) );
  XNOR2_X1 U379 ( .A(n313), .B(n344), .ZN(n319) );
  XOR2_X1 U380 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n315) );
  XNOR2_X1 U381 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n314) );
  XNOR2_X1 U382 ( .A(n315), .B(n314), .ZN(n317) );
  XNOR2_X1 U383 ( .A(G176GAT), .B(G106GAT), .ZN(n316) );
  XNOR2_X1 U384 ( .A(G78GAT), .B(KEYINPUT71), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n320), .B(G148GAT), .ZN(n430) );
  XOR2_X1 U386 ( .A(n321), .B(n430), .Z(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n576) );
  XNOR2_X1 U388 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n576), .B(n324), .ZN(n561) );
  XOR2_X1 U390 ( .A(G141GAT), .B(G197GAT), .Z(n326) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G50GAT), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n326), .B(n325), .ZN(n340) );
  XOR2_X1 U393 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n328) );
  NAND2_X1 U394 ( .A1(G229GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U396 ( .A(n329), .B(KEYINPUT29), .Z(n334) );
  XOR2_X1 U397 ( .A(G29GAT), .B(KEYINPUT8), .Z(n331) );
  XNOR2_X1 U398 ( .A(KEYINPUT68), .B(KEYINPUT7), .ZN(n330) );
  XNOR2_X1 U399 ( .A(n331), .B(n330), .ZN(n379) );
  XNOR2_X1 U400 ( .A(G22GAT), .B(G1GAT), .ZN(n332) );
  XNOR2_X1 U401 ( .A(n332), .B(G8GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n379), .B(n345), .ZN(n333) );
  XNOR2_X1 U403 ( .A(n334), .B(n333), .ZN(n336) );
  XOR2_X1 U404 ( .A(n336), .B(n335), .Z(n338) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(G43GAT), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n339) );
  NAND2_X1 U407 ( .A1(n561), .A2(n572), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n341), .B(KEYINPUT46), .ZN(n363) );
  XOR2_X1 U409 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n343) );
  XNOR2_X1 U410 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n343), .B(n342), .ZN(n349) );
  XOR2_X1 U412 ( .A(n344), .B(G183GAT), .Z(n347) );
  XNOR2_X1 U413 ( .A(n345), .B(G15GAT), .ZN(n346) );
  XNOR2_X1 U414 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n362) );
  XOR2_X1 U416 ( .A(G78GAT), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U417 ( .A(G127GAT), .B(G71GAT), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U419 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n353) );
  XNOR2_X1 U420 ( .A(G155GAT), .B(G57GAT), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U422 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U423 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n357) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U426 ( .A(G64GAT), .B(n358), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n490) );
  NAND2_X1 U429 ( .A1(n363), .A2(n490), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n364), .B(KEYINPUT113), .ZN(n382) );
  XOR2_X1 U431 ( .A(KEYINPUT67), .B(KEYINPUT75), .Z(n366) );
  XNOR2_X1 U432 ( .A(G99GAT), .B(G92GAT), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U434 ( .A(KEYINPUT11), .B(n395), .Z(n369) );
  XNOR2_X1 U435 ( .A(n367), .B(G85GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U438 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n373) );
  XNOR2_X1 U439 ( .A(G190GAT), .B(KEYINPUT76), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U441 ( .A(G106GAT), .B(G162GAT), .Z(n378) );
  XNOR2_X1 U442 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n439) );
  XNOR2_X1 U444 ( .A(n379), .B(n439), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n478) );
  NAND2_X1 U446 ( .A1(n382), .A2(n478), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n383), .B(KEYINPUT47), .ZN(n388) );
  XNOR2_X1 U448 ( .A(KEYINPUT36), .B(n478), .ZN(n486) );
  NOR2_X1 U449 ( .A1(n486), .A2(n490), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n384), .B(n289), .ZN(n385) );
  NAND2_X1 U451 ( .A1(n385), .A2(n576), .ZN(n386) );
  NOR2_X1 U452 ( .A1(n572), .A2(n386), .ZN(n387) );
  NOR2_X1 U453 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U454 ( .A(KEYINPUT48), .B(n389), .ZN(n539) );
  XOR2_X1 U455 ( .A(KEYINPUT94), .B(n390), .Z(n394) );
  XOR2_X1 U456 ( .A(G211GAT), .B(KEYINPUT21), .Z(n392) );
  XNOR2_X1 U457 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n437) );
  XNOR2_X1 U459 ( .A(G8GAT), .B(n437), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n454) );
  XNOR2_X1 U462 ( .A(n454), .B(KEYINPUT119), .ZN(n400) );
  NOR2_X1 U463 ( .A1(n539), .A2(n400), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n425) );
  XOR2_X1 U465 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n404) );
  XNOR2_X1 U466 ( .A(KEYINPUT92), .B(KEYINPUT1), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n410) );
  XOR2_X1 U468 ( .A(n405), .B(G134GAT), .Z(n408) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(n406), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U471 ( .A(n410), .B(n409), .Z(n412) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U474 ( .A(G148GAT), .B(G162GAT), .Z(n414) );
  XNOR2_X1 U475 ( .A(G113GAT), .B(G120GAT), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U477 ( .A(n416), .B(n415), .Z(n424) );
  XOR2_X1 U478 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n418) );
  XNOR2_X1 U479 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(G141GAT), .B(n419), .Z(n440) );
  XOR2_X1 U482 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n421) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n440), .B(n422), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n496) );
  NAND2_X1 U487 ( .A1(n425), .A2(n496), .ZN(n427) );
  INV_X1 U488 ( .A(KEYINPUT65), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n483) );
  XOR2_X1 U490 ( .A(G218GAT), .B(G204GAT), .Z(n429) );
  XNOR2_X1 U491 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U493 ( .A(n431), .B(n430), .Z(n436) );
  XOR2_X1 U494 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n433) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U497 ( .A(KEYINPUT24), .B(n434), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U499 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n462) );
  NOR2_X1 U502 ( .A1(n483), .A2(n462), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n443), .B(KEYINPUT55), .ZN(n444) );
  NOR2_X1 U504 ( .A1(n509), .A2(n444), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n569) );
  NAND2_X1 U506 ( .A1(n569), .A2(n561), .ZN(n450) );
  XOR2_X1 U507 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n448) );
  XNOR2_X1 U508 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n452) );
  NAND2_X1 U512 ( .A1(n462), .A2(n509), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n484) );
  XNOR2_X1 U514 ( .A(n454), .B(KEYINPUT95), .ZN(n453) );
  XNOR2_X1 U515 ( .A(n453), .B(KEYINPUT27), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n484), .A2(n461), .ZN(n555) );
  NAND2_X1 U517 ( .A1(n541), .A2(n454), .ZN(n455) );
  XOR2_X1 U518 ( .A(KEYINPUT98), .B(n455), .Z(n456) );
  NOR2_X1 U519 ( .A1(n462), .A2(n456), .ZN(n457) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n457), .Z(n458) );
  NOR2_X1 U521 ( .A1(n555), .A2(n458), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n459), .B(KEYINPUT99), .ZN(n460) );
  NAND2_X1 U523 ( .A1(n460), .A2(n496), .ZN(n467) );
  NOR2_X1 U524 ( .A1(n496), .A2(n461), .ZN(n463) );
  XOR2_X1 U525 ( .A(n462), .B(KEYINPUT28), .Z(n514) );
  NAND2_X1 U526 ( .A1(n463), .A2(n514), .ZN(n540) );
  XNOR2_X1 U527 ( .A(KEYINPUT87), .B(n509), .ZN(n464) );
  NOR2_X1 U528 ( .A1(n540), .A2(n464), .ZN(n465) );
  XOR2_X1 U529 ( .A(KEYINPUT96), .B(n465), .Z(n466) );
  NAND2_X1 U530 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U531 ( .A(KEYINPUT100), .B(n468), .ZN(n492) );
  INV_X1 U532 ( .A(n490), .ZN(n581) );
  NOR2_X1 U533 ( .A1(n486), .A2(n581), .ZN(n469) );
  NAND2_X1 U534 ( .A1(n492), .A2(n469), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n576), .A2(n572), .ZN(n495) );
  NOR2_X1 U536 ( .A1(n528), .A2(n495), .ZN(n473) );
  XOR2_X1 U537 ( .A(KEYINPUT38), .B(n473), .Z(n513) );
  NOR2_X1 U538 ( .A1(n496), .A2(n513), .ZN(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT39), .B(KEYINPUT105), .ZN(n475) );
  INV_X1 U540 ( .A(n478), .ZN(n566) );
  NAND2_X1 U541 ( .A1(n569), .A2(n566), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n480) );
  INV_X1 U543 ( .A(G190GAT), .ZN(n479) );
  NOR2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n486), .A2(n577), .ZN(n489) );
  NOR2_X1 U546 ( .A1(n490), .A2(n566), .ZN(n491) );
  XNOR2_X1 U547 ( .A(KEYINPUT16), .B(n491), .ZN(n493) );
  NAND2_X1 U548 ( .A1(n493), .A2(n492), .ZN(n494) );
  XOR2_X1 U549 ( .A(KEYINPUT101), .B(n494), .Z(n518) );
  NOR2_X1 U550 ( .A1(n495), .A2(n518), .ZN(n504) );
  INV_X1 U551 ( .A(n496), .ZN(n554) );
  NAND2_X1 U552 ( .A1(n504), .A2(n554), .ZN(n497) );
  XNOR2_X1 U553 ( .A(n497), .B(KEYINPUT34), .ZN(n498) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n504), .A2(n454), .ZN(n499) );
  XNOR2_X1 U556 ( .A(n499), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n501) );
  NAND2_X1 U558 ( .A1(n504), .A2(n541), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(n503) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT102), .Z(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  INV_X1 U562 ( .A(n514), .ZN(n535) );
  NAND2_X1 U563 ( .A1(n504), .A2(n535), .ZN(n505) );
  XNOR2_X1 U564 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  INV_X1 U565 ( .A(n454), .ZN(n506) );
  NOR2_X1 U566 ( .A1(n513), .A2(n506), .ZN(n507) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(n507), .Z(n508) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n508), .ZN(G1329GAT) );
  NOR2_X1 U569 ( .A1(n513), .A2(n509), .ZN(n511) );
  XNOR2_X1 U570 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U574 ( .A(KEYINPUT108), .B(n515), .Z(n516) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(n516), .ZN(G1331GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n520) );
  INV_X1 U577 ( .A(n572), .ZN(n517) );
  NAND2_X1 U578 ( .A1(n517), .A2(n561), .ZN(n527) );
  NOR2_X1 U579 ( .A1(n518), .A2(n527), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n524), .A2(n554), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n524), .A2(n454), .ZN(n522) );
  XNOR2_X1 U584 ( .A(n522), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n524), .A2(n541), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .Z(n526) );
  NAND2_X1 U588 ( .A1(n524), .A2(n535), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n534), .A2(n554), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n529), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n534), .A2(n454), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n534), .A2(n541), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n533) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT110), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1339GAT) );
  XOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT115), .Z(n545) );
  NOR2_X1 U604 ( .A1(n539), .A2(n540), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT114), .B(n543), .Z(n551) );
  NAND2_X1 U607 ( .A1(n551), .A2(n572), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U610 ( .A1(n561), .A2(n551), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n549) );
  NAND2_X1 U613 ( .A1(n551), .A2(n581), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n550), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n566), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U620 ( .A1(n539), .A2(n556), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n572), .A2(n565), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n559) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT117), .B(n560), .Z(n563) );
  NAND2_X1 U627 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n581), .A2(n565), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n572), .A2(n569), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT123), .Z(n571) );
  NAND2_X1 U636 ( .A1(n569), .A2(n581), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  NAND2_X1 U639 ( .A1(n582), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n579) );
  OR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1354GAT) );
endmodule

