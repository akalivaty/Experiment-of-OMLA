

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588;

  AND2_X1 U321 ( .A1(n567), .A2(n553), .ZN(n325) );
  XNOR2_X1 U322 ( .A(n300), .B(G85GAT), .ZN(n351) );
  NOR2_X1 U323 ( .A1(n564), .A2(n368), .ZN(n369) );
  XNOR2_X1 U324 ( .A(n479), .B(KEYINPUT104), .ZN(n480) );
  OR2_X1 U325 ( .A1(n291), .A2(n569), .ZN(n571) );
  XNOR2_X1 U326 ( .A(n388), .B(n387), .ZN(n524) );
  XNOR2_X1 U327 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n289) );
  XOR2_X1 U328 ( .A(G190GAT), .B(G218GAT), .Z(n290) );
  NAND2_X1 U329 ( .A1(n568), .A2(n567), .ZN(n291) );
  XNOR2_X1 U330 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n365) );
  XNOR2_X1 U331 ( .A(n366), .B(n365), .ZN(n367) );
  INV_X1 U332 ( .A(G99GAT), .ZN(n300) );
  AND2_X1 U333 ( .A1(n362), .A2(n361), .ZN(n363) );
  XNOR2_X1 U334 ( .A(n432), .B(n289), .ZN(n298) );
  INV_X1 U335 ( .A(n380), .ZN(n381) );
  XNOR2_X1 U336 ( .A(n299), .B(n298), .ZN(n302) );
  XNOR2_X1 U337 ( .A(n354), .B(n290), .ZN(n355) );
  INV_X1 U338 ( .A(KEYINPUT37), .ZN(n479) );
  XNOR2_X1 U339 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U340 ( .A(n417), .B(n416), .ZN(n458) );
  XNOR2_X1 U341 ( .A(n356), .B(n355), .ZN(n358) );
  XNOR2_X1 U342 ( .A(n384), .B(n383), .ZN(n386) );
  XNOR2_X1 U343 ( .A(n481), .B(n480), .ZN(n521) );
  NOR2_X1 U344 ( .A1(n569), .A2(n526), .ZN(n563) );
  XNOR2_X1 U345 ( .A(n360), .B(n359), .ZN(n560) );
  INV_X1 U346 ( .A(G43GAT), .ZN(n483) );
  XNOR2_X1 U347 ( .A(n460), .B(G218GAT), .ZN(n461) );
  XNOR2_X1 U348 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U349 ( .A(n483), .B(KEYINPUT40), .ZN(n484) );
  XNOR2_X1 U350 ( .A(n462), .B(n461), .ZN(G1355GAT) );
  XNOR2_X1 U351 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n485), .B(n484), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(G92GAT), .B(G64GAT), .Z(n293) );
  XNOR2_X1 U354 ( .A(G176GAT), .B(G204GAT), .ZN(n292) );
  XNOR2_X1 U355 ( .A(n293), .B(n292), .ZN(n295) );
  INV_X1 U356 ( .A(KEYINPUT74), .ZN(n294) );
  XNOR2_X1 U357 ( .A(n295), .B(n294), .ZN(n378) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G71GAT), .Z(n443) );
  XNOR2_X1 U359 ( .A(n378), .B(n443), .ZN(n299) );
  XOR2_X1 U360 ( .A(KEYINPUT73), .B(G78GAT), .Z(n297) );
  XNOR2_X1 U361 ( .A(G148GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U362 ( .A(n297), .B(n296), .ZN(n432) );
  XOR2_X1 U363 ( .A(G57GAT), .B(KEYINPUT13), .Z(n332) );
  XNOR2_X1 U364 ( .A(n351), .B(n332), .ZN(n301) );
  XOR2_X1 U365 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U366 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n304) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U369 ( .A(KEYINPUT71), .B(n305), .Z(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n582) );
  XNOR2_X1 U371 ( .A(KEYINPUT41), .B(n582), .ZN(n567) );
  XOR2_X1 U372 ( .A(G1GAT), .B(G15GAT), .Z(n329) );
  XOR2_X1 U373 ( .A(G141GAT), .B(G22GAT), .Z(n421) );
  XOR2_X1 U374 ( .A(n329), .B(n421), .Z(n309) );
  NAND2_X1 U375 ( .A1(G229GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U376 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U377 ( .A(G169GAT), .B(G8GAT), .Z(n379) );
  XOR2_X1 U378 ( .A(n310), .B(n379), .Z(n318) );
  XOR2_X1 U379 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n312) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(G197GAT), .ZN(n311) );
  XNOR2_X1 U381 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U382 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n314) );
  XNOR2_X1 U383 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n313) );
  XNOR2_X1 U384 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U385 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U386 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U387 ( .A(G29GAT), .B(KEYINPUT7), .Z(n320) );
  XNOR2_X1 U388 ( .A(G43GAT), .B(G36GAT), .ZN(n319) );
  XNOR2_X1 U389 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U390 ( .A(G50GAT), .B(KEYINPUT8), .Z(n321) );
  XNOR2_X1 U391 ( .A(n322), .B(n321), .ZN(n346) );
  XOR2_X1 U392 ( .A(n323), .B(n346), .Z(n577) );
  INV_X1 U393 ( .A(n577), .ZN(n553) );
  XNOR2_X1 U394 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n324) );
  XNOR2_X1 U395 ( .A(n325), .B(n324), .ZN(n362) );
  XOR2_X1 U396 ( .A(KEYINPUT78), .B(G211GAT), .Z(n327) );
  XNOR2_X1 U397 ( .A(G127GAT), .B(G155GAT), .ZN(n326) );
  XNOR2_X1 U398 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U399 ( .A(n328), .B(G64GAT), .Z(n331) );
  XNOR2_X1 U400 ( .A(G8GAT), .B(n329), .ZN(n330) );
  XNOR2_X1 U401 ( .A(n331), .B(n330), .ZN(n345) );
  XOR2_X1 U402 ( .A(n332), .B(G78GAT), .Z(n334) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U404 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U405 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n336) );
  XNOR2_X1 U406 ( .A(G71GAT), .B(KEYINPUT15), .ZN(n335) );
  XNOR2_X1 U407 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U408 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U409 ( .A(G183GAT), .B(KEYINPUT76), .Z(n380) );
  XOR2_X1 U410 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n340) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(KEYINPUT14), .ZN(n339) );
  XNOR2_X1 U412 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U413 ( .A(n380), .B(n341), .ZN(n342) );
  XNOR2_X1 U414 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U415 ( .A(n345), .B(n344), .Z(n587) );
  INV_X1 U416 ( .A(n587), .ZN(n574) );
  INV_X1 U417 ( .A(n346), .ZN(n350) );
  XOR2_X1 U418 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n348) );
  XNOR2_X1 U419 ( .A(G92GAT), .B(KEYINPUT65), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U421 ( .A(n350), .B(n349), .ZN(n360) );
  XOR2_X1 U422 ( .A(KEYINPUT10), .B(n351), .Z(n356) );
  XOR2_X1 U423 ( .A(G106GAT), .B(KEYINPUT9), .Z(n353) );
  XNOR2_X1 U424 ( .A(G134GAT), .B(G162GAT), .ZN(n352) );
  XNOR2_X1 U425 ( .A(n353), .B(n352), .ZN(n354) );
  NAND2_X1 U426 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n359) );
  NOR2_X1 U428 ( .A1(n574), .A2(n560), .ZN(n361) );
  XOR2_X1 U429 ( .A(KEYINPUT47), .B(n363), .Z(n371) );
  XNOR2_X1 U430 ( .A(KEYINPUT70), .B(n553), .ZN(n564) );
  INV_X1 U431 ( .A(KEYINPUT36), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n364), .B(n560), .ZN(n477) );
  NOR2_X1 U433 ( .A1(n587), .A2(n477), .ZN(n366) );
  NAND2_X1 U434 ( .A1(n367), .A2(n582), .ZN(n368) );
  XOR2_X1 U435 ( .A(KEYINPUT113), .B(n369), .Z(n370) );
  NOR2_X1 U436 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U437 ( .A(KEYINPUT48), .B(n372), .ZN(n548) );
  XOR2_X1 U438 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n374) );
  XNOR2_X1 U439 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n448) );
  XOR2_X1 U441 ( .A(G211GAT), .B(KEYINPUT21), .Z(n376) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(G218GAT), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n433) );
  XNOR2_X1 U444 ( .A(n448), .B(n433), .ZN(n388) );
  INV_X1 U445 ( .A(KEYINPUT97), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n384) );
  XNOR2_X1 U447 ( .A(G36GAT), .B(n379), .ZN(n382) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n387) );
  NOR2_X1 U450 ( .A1(n548), .A2(n524), .ZN(n390) );
  XNOR2_X1 U451 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n415) );
  XOR2_X1 U453 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n392) );
  XNOR2_X1 U454 ( .A(G113GAT), .B(G127GAT), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U456 ( .A(G134GAT), .B(KEYINPUT0), .Z(n393) );
  XOR2_X1 U457 ( .A(n394), .B(n393), .Z(n453) );
  XOR2_X1 U458 ( .A(G155GAT), .B(KEYINPUT3), .Z(n396) );
  XNOR2_X1 U459 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n425) );
  XNOR2_X1 U461 ( .A(G1GAT), .B(n425), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n397), .B(G57GAT), .ZN(n401) );
  XOR2_X1 U463 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n399) );
  XNOR2_X1 U464 ( .A(G141GAT), .B(KEYINPUT96), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U467 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n403) );
  XNOR2_X1 U468 ( .A(G120GAT), .B(KEYINPUT94), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n453), .B(n406), .ZN(n414) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n412) );
  XOR2_X1 U473 ( .A(G148GAT), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n407) );
  XNOR2_X1 U475 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U476 ( .A(G29GAT), .B(G85GAT), .Z(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n522) );
  NAND2_X1 U480 ( .A1(n415), .A2(n522), .ZN(n417) );
  INV_X1 U481 ( .A(KEYINPUT64), .ZN(n416) );
  XOR2_X1 U482 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n419) );
  XNOR2_X1 U483 ( .A(G50GAT), .B(G204GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U485 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U488 ( .A(n424), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U489 ( .A(n425), .B(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n429) );
  XNOR2_X1 U492 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n467) );
  NAND2_X1 U497 ( .A1(n458), .A2(n467), .ZN(n437) );
  INV_X1 U498 ( .A(KEYINPUT55), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n569) );
  XOR2_X1 U500 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n439) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(G15GAT), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n452) );
  XOR2_X1 U503 ( .A(G176GAT), .B(G183GAT), .Z(n441) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G99GAT), .ZN(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n445) );
  AND2_X1 U507 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n447) );
  INV_X1 U509 ( .A(KEYINPUT86), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n448), .B(KEYINPUT20), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n568) );
  INV_X1 U515 ( .A(n568), .ZN(n526) );
  NAND2_X1 U516 ( .A1(n563), .A2(n560), .ZN(n456) );
  NOR2_X1 U517 ( .A1(n467), .A2(n568), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT26), .ZN(n551) );
  NAND2_X1 U519 ( .A1(n551), .A2(n458), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT124), .ZN(n586) );
  NOR2_X1 U521 ( .A1(n477), .A2(n586), .ZN(n462) );
  XNOR2_X1 U522 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n460) );
  NAND2_X1 U523 ( .A1(n582), .A2(n564), .ZN(n491) );
  INV_X1 U524 ( .A(KEYINPUT27), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n524), .B(n463), .ZN(n469) );
  INV_X1 U526 ( .A(n469), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n464), .A2(n522), .ZN(n465) );
  XOR2_X1 U528 ( .A(KEYINPUT98), .B(n465), .Z(n549) );
  XOR2_X1 U529 ( .A(n467), .B(KEYINPUT28), .Z(n500) );
  NOR2_X1 U530 ( .A1(n549), .A2(n500), .ZN(n534) );
  NAND2_X1 U531 ( .A1(n534), .A2(n526), .ZN(n475) );
  OR2_X1 U532 ( .A1(n526), .A2(n524), .ZN(n466) );
  NAND2_X1 U533 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U534 ( .A(KEYINPUT25), .B(n468), .Z(n471) );
  NAND2_X1 U535 ( .A1(n469), .A2(n551), .ZN(n470) );
  AND2_X1 U536 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(n472), .ZN(n473) );
  NAND2_X1 U538 ( .A1(n473), .A2(n522), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U540 ( .A(KEYINPUT100), .B(n476), .ZN(n489) );
  NOR2_X1 U541 ( .A1(n574), .A2(n477), .ZN(n478) );
  NAND2_X1 U542 ( .A1(n489), .A2(n478), .ZN(n481) );
  NOR2_X1 U543 ( .A1(n491), .A2(n521), .ZN(n482) );
  XOR2_X1 U544 ( .A(KEYINPUT38), .B(n482), .Z(n506) );
  NOR2_X1 U545 ( .A1(n506), .A2(n526), .ZN(n485) );
  INV_X1 U546 ( .A(n560), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n574), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT16), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT81), .B(n488), .ZN(n490) );
  NAND2_X1 U550 ( .A1(n490), .A2(n489), .ZN(n510) );
  OR2_X1 U551 ( .A1(n491), .A2(n510), .ZN(n501) );
  NOR2_X1 U552 ( .A1(n522), .A2(n501), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT34), .B(n492), .Z(n493) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U555 ( .A1(n524), .A2(n501), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1325GAT) );
  NOR2_X1 U558 ( .A1(n501), .A2(n526), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n497) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1326GAT) );
  INV_X1 U563 ( .A(n500), .ZN(n531) );
  NOR2_X1 U564 ( .A1(n531), .A2(n501), .ZN(n502) );
  XOR2_X1 U565 ( .A(G22GAT), .B(n502), .Z(G1327GAT) );
  NOR2_X1 U566 ( .A1(n506), .A2(n522), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n524), .A2(n506), .ZN(n505) );
  XOR2_X1 U570 ( .A(G36GAT), .B(n505), .Z(G1329GAT) );
  NOR2_X1 U571 ( .A1(n506), .A2(n531), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  NAND2_X1 U574 ( .A1(n567), .A2(n577), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(KEYINPUT106), .ZN(n520) );
  OR2_X1 U576 ( .A1(n520), .A2(n510), .ZN(n516) );
  NOR2_X1 U577 ( .A1(n522), .A2(n516), .ZN(n512) );
  XNOR2_X1 U578 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n524), .A2(n516), .ZN(n514) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n514), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n526), .A2(n516), .ZN(n515) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n515), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n531), .A2(n516), .ZN(n518) );
  XNOR2_X1 U586 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U589 ( .A1(n521), .A2(n520), .ZN(n530) );
  NOR2_X1 U590 ( .A1(n522), .A2(n530), .ZN(n523) );
  XOR2_X1 U591 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U592 ( .A1(n524), .A2(n530), .ZN(n525) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n530), .ZN(n527) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n529) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(n533) );
  NOR2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U600 ( .A(n533), .B(n532), .Z(G1339GAT) );
  NAND2_X1 U601 ( .A1(n568), .A2(n534), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n535), .A2(n548), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT114), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n544), .A2(n564), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U607 ( .A1(n544), .A2(n567), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U609 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U611 ( .A1(n544), .A2(n574), .ZN(n541) );
  XNOR2_X1 U612 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U613 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U615 ( .A1(n560), .A2(n544), .ZN(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NOR2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(n552), .Z(n561) );
  NAND2_X1 U621 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U624 ( .A1(n561), .A2(n567), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n574), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U632 ( .A(G169GAT), .B(KEYINPUT121), .Z(n566) );
  NAND2_X1 U633 ( .A1(n563), .A2(n564), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XNOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n573) );
  XOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT56), .Z(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  XOR2_X1 U639 ( .A(G183GAT), .B(KEYINPUT123), .Z(n576) );
  NAND2_X1 U640 ( .A1(n563), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n586), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XNOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n584) );
  NOR2_X1 U648 ( .A1(n586), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G204GAT), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n588), .Z(G1354GAT) );
endmodule

