//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT67), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(G116), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(KEYINPUT5), .A3(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G119), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT5), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G116), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(G113), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G113), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G113), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n196), .A2(new_n198), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G104), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(G107), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n210), .B2(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n211), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n220), .A2(new_n222), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n203), .A2(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT84), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n191), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n196), .A2(KEYINPUT5), .A3(new_n198), .ZN(new_n230));
  OAI21_X1  g044(.A(G113), .B1(new_n196), .B2(KEYINPUT5), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n209), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n221), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n203), .A2(new_n209), .A3(new_n221), .A4(new_n226), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(KEYINPUT84), .A3(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n229), .A2(new_n236), .A3(KEYINPUT85), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT85), .B1(new_n229), .B2(new_n236), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n232), .B2(new_n233), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n226), .A2(new_n221), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n242), .A2(KEYINPUT80), .A3(new_n209), .A4(new_n203), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n216), .B1(new_n217), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n220), .B1(new_n211), .B2(new_n212), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n196), .A2(new_n198), .ZN(new_n249));
  INV_X1    g063(.A(new_n208), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n209), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(G101), .C1(new_n245), .C2(new_n246), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n241), .A2(new_n243), .A3(new_n255), .A4(new_n189), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT64), .B1(new_n259), .B2(G143), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT64), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n257), .A3(G146), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n263), .A2(new_n264), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G125), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(KEYINPUT1), .C1(new_n257), .C2(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G128), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n265), .B2(KEYINPUT1), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n267), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n260), .A2(new_n262), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n279), .A3(G128), .A4(new_n265), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n280), .A3(new_n271), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT81), .B(G224), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G953), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n283), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n272), .A2(new_n281), .A3(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n288), .A2(KEYINPUT86), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(KEYINPUT86), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n256), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n188), .B1(new_n239), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n241), .A2(new_n243), .A3(new_n255), .ZN(new_n293));
  INV_X1    g107(.A(new_n189), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT6), .A3(new_n256), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n282), .B(new_n285), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n293), .A2(new_n298), .A3(new_n294), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n296), .A2(KEYINPUT82), .A3(new_n297), .A4(new_n299), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n292), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G210), .B1(G237), .B2(G902), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n187), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n303), .ZN(new_n307));
  INV_X1    g121(.A(new_n292), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n305), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G214), .B1(G237), .B2(G902), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n187), .A3(new_n310), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT88), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n312), .A2(new_n317), .A3(new_n313), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G217), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(G234), .B2(new_n188), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n200), .B2(G128), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n193), .A2(new_n195), .A3(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n326));
  INV_X1    g140(.A(G128), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n194), .A2(G119), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n192), .A2(KEYINPUT67), .ZN(new_n329));
  OAI211_X1 g143(.A(KEYINPUT75), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G110), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n192), .A2(G128), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT23), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n200), .B2(G128), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  OR2_X1    g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n271), .A2(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(G146), .B(new_n342), .C1(new_n345), .C2(new_n340), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n259), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n342), .B1(new_n345), .B2(new_n340), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n259), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n351), .A2(new_n346), .B1(new_n336), .B2(new_n337), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g169(.A(KEYINPUT76), .B(new_n332), .C1(new_n331), .C2(new_n334), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G137), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n359), .A2(G221), .A3(G234), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n361), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n349), .B(new_n363), .C1(new_n355), .C2(new_n356), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n188), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n364), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n322), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n362), .A2(new_n364), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n370), .A2(G902), .A3(new_n321), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT69), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n277), .A2(new_n280), .ZN(new_n375));
  INV_X1    g189(.A(G137), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT65), .A3(G134), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT65), .ZN(new_n378));
  INV_X1    g192(.A(G134), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(G137), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n376), .A2(G134), .ZN(new_n381));
  OAI211_X1 g195(.A(G131), .B(new_n377), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT11), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n379), .B2(G137), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n376), .A2(KEYINPUT11), .A3(G134), .ZN(new_n385));
  INV_X1    g199(.A(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n379), .A2(G137), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G131), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n388), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n375), .A2(new_n390), .B1(new_n393), .B2(new_n270), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n196), .A2(new_n198), .A3(new_n208), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n208), .B1(new_n196), .B2(new_n198), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n374), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n375), .A2(new_n390), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n270), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT68), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n395), .B2(new_n396), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n251), .A2(KEYINPUT68), .A3(new_n209), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n399), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n393), .A2(new_n270), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n389), .B1(new_n280), .B2(new_n277), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT69), .B(new_n252), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n398), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n409));
  NOR2_X1   g223(.A1(G237), .A2(G953), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G210), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G101), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n402), .A2(new_n403), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n416), .A2(KEYINPUT69), .B1(new_n417), .B2(new_n394), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n415), .B1(new_n418), .B2(new_n398), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n404), .A2(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT70), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n409), .B(new_n414), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n408), .A2(KEYINPUT28), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n421), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n414), .A4(new_n409), .ZN(new_n428));
  INV_X1    g242(.A(new_n404), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT30), .B1(new_n405), .B2(new_n406), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n399), .A2(new_n431), .A3(new_n400), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n429), .B1(new_n433), .B2(new_n252), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(new_n414), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT29), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n424), .A2(new_n428), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n399), .A2(new_n400), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n402), .A2(new_n403), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT73), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n404), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(KEYINPUT73), .A3(new_n439), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(KEYINPUT28), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n414), .A2(KEYINPUT29), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n420), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT74), .B1(new_n446), .B2(new_n188), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(KEYINPUT74), .A3(new_n188), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G472), .B1(new_n437), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n452));
  INV_X1    g266(.A(new_n414), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n408), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n408), .A2(KEYINPUT28), .B1(KEYINPUT70), .B2(new_n420), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT30), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n431), .B1(new_n399), .B2(new_n400), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n252), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n414), .A3(new_n404), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT31), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n434), .A2(KEYINPUT31), .A3(new_n414), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(G472), .A2(G902), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n452), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT32), .ZN(new_n468));
  INV_X1    g282(.A(new_n466), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n468), .B(new_n469), .C1(new_n456), .C2(new_n464), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n373), .B1(new_n451), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT17), .ZN(new_n473));
  INV_X1    g287(.A(G237), .ZN(new_n474));
  AND4_X1   g288(.A1(G143), .A2(new_n474), .A3(new_n359), .A4(G214), .ZN(new_n475));
  AOI21_X1  g289(.A(G143), .B1(new_n410), .B2(G214), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n359), .A3(G214), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n257), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n410), .A2(G143), .A3(G214), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(G131), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n473), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n351), .A2(new_n346), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT91), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n482), .B2(G131), .ZN(new_n488));
  AOI211_X1 g302(.A(KEYINPUT90), .B(new_n386), .C1(new_n480), .C2(new_n481), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT17), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n351), .A2(new_n346), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n480), .A2(new_n386), .A3(new_n481), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n478), .A2(new_n484), .A3(new_n473), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(KEYINPUT18), .A2(G131), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n345), .A2(G146), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n482), .A2(new_n497), .B1(new_n498), .B2(new_n347), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n482), .A2(new_n497), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n215), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n496), .A2(new_n506), .A3(new_n503), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n188), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G475), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n478), .A2(new_n484), .A3(new_n494), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n345), .B(KEYINPUT19), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n346), .C1(G146), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n503), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n509), .B2(new_n517), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(KEYINPUT20), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n518), .A2(new_n521), .A3(new_n524), .A4(new_n519), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G952), .ZN(new_n527));
  AOI211_X1 g341(.A(G953), .B(new_n527), .C1(G234), .C2(G237), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n188), .B(new_n359), .C1(G234), .C2(G237), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT21), .B(G898), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G478), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT9), .B(G234), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n535), .A2(new_n320), .A3(G953), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n327), .A2(G143), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n379), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n257), .A2(G128), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n538), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n540), .B(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G122), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT93), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G122), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n197), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n544), .A2(G116), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT94), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n551));
  INV_X1    g365(.A(new_n549), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT93), .B(G122), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n197), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G107), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n210), .A3(new_n554), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n543), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT95), .B1(new_n541), .B2(new_n538), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n541), .A2(new_n538), .A3(KEYINPUT95), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n379), .A3(new_n561), .ZN(new_n562));
  OR3_X1    g376(.A1(new_n544), .A2(KEYINPUT14), .A3(G116), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT14), .B1(new_n544), .B2(G116), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G107), .B1(new_n565), .B2(new_n548), .ZN(new_n566));
  INV_X1    g380(.A(new_n561), .ZN(new_n567));
  OAI21_X1  g381(.A(G134), .B1(new_n567), .B2(new_n559), .ZN(new_n568));
  AND4_X1   g382(.A1(new_n557), .A2(new_n562), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n537), .B1(new_n558), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n543), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n550), .A2(new_n210), .A3(new_n554), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n210), .B1(new_n550), .B2(new_n554), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n557), .A2(new_n562), .A3(new_n566), .A4(new_n568), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n536), .ZN(new_n576));
  AOI21_X1  g390(.A(G902), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n534), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n574), .A2(new_n575), .A3(new_n536), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n536), .B1(new_n574), .B2(new_n575), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n188), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT96), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n578), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n579), .B1(new_n585), .B2(new_n534), .ZN(new_n586));
  AND4_X1   g400(.A1(new_n512), .A2(new_n526), .A3(new_n532), .A4(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G221), .B1(new_n535), .B2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n254), .A2(new_n270), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n279), .A2(G128), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n591), .B(new_n258), .C1(new_n260), .C2(new_n262), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n278), .A2(new_n265), .B1(new_n593), .B2(G128), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n221), .B(new_n226), .C1(new_n592), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n248), .A2(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT79), .ZN(new_n598));
  INV_X1    g412(.A(new_n393), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n242), .A2(KEYINPUT10), .A3(new_n375), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n597), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n595), .A2(new_n596), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n210), .A2(G104), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n216), .B2(new_n217), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n219), .B1(new_n605), .B2(new_n214), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n270), .B(new_n254), .C1(new_n603), .C2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n602), .A2(new_n599), .A3(new_n600), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n233), .A2(new_n280), .A3(new_n277), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n599), .B1(new_n611), .B2(new_n595), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(G110), .B(G140), .ZN(new_n615));
  INV_X1    g429(.A(G227), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(G953), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n615), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n601), .B2(new_n609), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n597), .A2(new_n600), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n393), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n614), .A2(new_n618), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(G469), .B1(new_n622), .B2(G902), .ZN(new_n623));
  INV_X1    g437(.A(G469), .ZN(new_n624));
  INV_X1    g438(.A(new_n618), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n610), .A2(new_n625), .A3(new_n613), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n610), .B2(new_n621), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n624), .B(new_n188), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n589), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n587), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n319), .A2(new_n472), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  NAND2_X1  g446(.A1(new_n622), .A2(G469), .ZN(new_n633));
  NAND2_X1  g447(.A1(G469), .A2(G902), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n635), .A2(new_n372), .A3(new_n588), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n465), .B2(new_n188), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n469), .B1(new_n456), .B2(new_n464), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n304), .B2(new_n305), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n311), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n309), .A2(new_n642), .A3(new_n310), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n313), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n523), .A2(new_n525), .B1(G475), .B2(new_n511), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT98), .B(G478), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n577), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n570), .A2(new_n576), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT33), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n188), .A2(G478), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n648), .A2(new_n531), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n641), .A2(new_n647), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  AOI21_X1  g472(.A(new_n524), .B1(new_n518), .B2(new_n519), .ZN(new_n659));
  INV_X1    g473(.A(new_n519), .ZN(new_n660));
  AOI211_X1 g474(.A(KEYINPUT20), .B(new_n660), .C1(new_n509), .C2(new_n517), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n508), .B2(new_n509), .ZN(new_n662));
  INV_X1    g476(.A(G475), .ZN(new_n663));
  OAI22_X1  g477(.A1(new_n659), .A2(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n664), .A2(new_n586), .A3(new_n531), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n647), .A2(new_n641), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n367), .A2(new_n368), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n321), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n361), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n357), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n321), .A2(G902), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n670), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n675), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT99), .B1(new_n369), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n679), .A2(new_n640), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n319), .A2(new_n630), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT100), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT37), .B(G110), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n528), .B1(new_n529), .B2(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n664), .A2(new_n586), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n671), .B1(new_n670), .B2(new_n675), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n369), .A2(new_n677), .A3(KEYINPUT99), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n629), .B(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n446), .A2(KEYINPUT74), .A3(new_n188), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n447), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n424), .A2(new_n428), .A3(new_n436), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n637), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n414), .B1(new_n426), .B2(new_n409), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT31), .B1(new_n434), .B2(new_n414), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n397), .B1(new_n430), .B2(new_n432), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n697), .A2(new_n461), .A3(new_n429), .A4(new_n453), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g513(.A(KEYINPUT32), .B(new_n466), .C1(new_n695), .C2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n639), .B2(new_n452), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n646), .A2(new_n690), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n327), .ZN(G30));
  XOR2_X1   g518(.A(new_n686), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n629), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT101), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n312), .A2(new_n314), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT38), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n712));
  INV_X1    g526(.A(new_n679), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n648), .A2(new_n586), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n313), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n460), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n442), .A2(new_n453), .A3(new_n443), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n188), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n701), .B1(G472), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n709), .A2(new_n711), .A3(new_n712), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT102), .B(G143), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G45));
  NAND2_X1  g537(.A1(new_n451), .A2(new_n471), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n648), .A2(new_n654), .A3(new_n686), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n629), .A3(new_n679), .A4(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT103), .B1(new_n726), .B2(new_n646), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n679), .A3(new_n629), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n702), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n647), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NAND4_X1  g547(.A1(new_n644), .A2(new_n655), .A3(new_n313), .A4(new_n645), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n610), .A2(new_n621), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n735), .A2(new_n618), .B1(new_n619), .B2(new_n613), .ZN(new_n736));
  OAI21_X1  g550(.A(G469), .B1(new_n736), .B2(G902), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n737), .A2(new_n588), .A3(new_n628), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(new_n372), .C1(new_n694), .C2(new_n701), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT41), .B(G113), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND4_X1  g556(.A1(new_n644), .A2(new_n313), .A3(new_n645), .A4(new_n665), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n739), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n197), .ZN(G18));
  OAI211_X1 g559(.A(new_n587), .B(new_n679), .C1(new_n701), .C2(new_n694), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n644), .A2(new_n313), .A3(new_n645), .A4(new_n738), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n192), .ZN(G21));
  NAND4_X1  g563(.A1(new_n644), .A2(new_n313), .A3(new_n645), .A4(new_n714), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n444), .A2(new_n420), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n453), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n469), .B1(new_n464), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n638), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n738), .A3(new_n372), .A4(new_n532), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n544), .ZN(G24));
  NAND3_X1  g571(.A1(new_n725), .A2(new_n679), .A3(new_n754), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n747), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n271), .ZN(G27));
  INV_X1    g574(.A(new_n313), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n312), .B2(new_n314), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(new_n472), .A3(new_n629), .A4(new_n725), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n639), .A2(KEYINPUT32), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n470), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n373), .B1(new_n451), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n762), .A4(new_n629), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  AND4_X1   g586(.A1(new_n472), .A2(new_n762), .A3(new_n629), .A4(new_n687), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n379), .ZN(G36));
  OR2_X1    g588(.A1(new_n622), .A2(KEYINPUT45), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n622), .A2(KEYINPUT45), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(G469), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n634), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n634), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(KEYINPUT105), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(KEYINPUT105), .ZN(new_n781));
  OAI221_X1 g595(.A(new_n628), .B1(KEYINPUT46), .B2(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n588), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n705), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n654), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n648), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT43), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n789), .A2(new_n640), .A3(new_n713), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT107), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n762), .B1(new_n790), .B2(new_n791), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n786), .B(new_n795), .C1(KEYINPUT107), .C2(new_n792), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  XNOR2_X1  g611(.A(new_n783), .B(KEYINPUT47), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n702), .A2(new_n373), .A3(new_n725), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n762), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NOR2_X1   g615(.A1(new_n703), .A2(new_n759), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n369), .A2(new_n677), .A3(new_n686), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n629), .A2(new_n803), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n750), .A2(new_n719), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n730), .B1(new_n729), .B2(new_n647), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n646), .A2(new_n728), .A3(KEYINPUT103), .A4(new_n702), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n802), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n732), .A2(KEYINPUT52), .A3(new_n802), .A4(new_n805), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(KEYINPUT109), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n773), .B1(new_n765), .B2(new_n770), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n577), .A2(new_n578), .ZN(new_n814));
  AOI211_X1 g628(.A(KEYINPUT96), .B(G902), .C1(new_n570), .C2(new_n576), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n534), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n579), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n526), .A2(new_n512), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n648), .B2(new_n654), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n636), .A2(new_n820), .A3(new_n532), .A4(new_n640), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n316), .B2(new_n318), .ZN(new_n822));
  OAI22_X1  g636(.A1(new_n747), .A2(new_n746), .B1(new_n750), .B2(new_n755), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n739), .B1(new_n734), .B2(new_n743), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n710), .A2(new_n313), .A3(new_n629), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n758), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n664), .A2(new_n818), .A3(new_n686), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n724), .A2(new_n629), .A3(new_n679), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n710), .A2(new_n313), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n679), .A2(new_n629), .A3(new_n829), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(KEYINPUT108), .A3(new_n762), .A4(new_n724), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n827), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n319), .B(new_n630), .C1(new_n680), .C2(new_n472), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n813), .A2(new_n825), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT109), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n808), .A2(new_n839), .A3(new_n809), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n812), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n810), .A2(new_n811), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT110), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n844), .A2(new_n838), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n842), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n813), .A2(new_n825), .A3(new_n836), .A4(new_n837), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n842), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n812), .A3(new_n840), .ZN(new_n854));
  XOR2_X1   g668(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n855));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT110), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n846), .A2(new_n857), .A3(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n849), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n528), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n789), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n372), .A3(new_n754), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n831), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n737), .A2(new_n628), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n588), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n798), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n738), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n862), .A2(new_n711), .A3(new_n313), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n869));
  AND2_X1   g683(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n831), .A2(new_n867), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n861), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n679), .A2(new_n754), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n868), .A2(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n372), .A3(new_n528), .A4(new_n719), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT113), .Z(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n648), .A3(new_n654), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n866), .A2(new_n871), .A3(new_n875), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n873), .A2(new_n768), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT48), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n862), .A2(new_n747), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n527), .B(G953), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n884), .B(new_n887), .C1(new_n886), .C2(new_n885), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n648), .A2(new_n654), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n877), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n859), .A2(new_n881), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n864), .A2(KEYINPUT49), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n864), .A2(KEYINPUT49), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n372), .A2(new_n313), .A3(new_n588), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n788), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n719), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n892), .A2(new_n893), .B1(new_n711), .B2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n188), .B1(new_n851), .B2(new_n854), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n296), .A2(new_n299), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n297), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT115), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n359), .A2(G952), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n901), .A2(new_n904), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n851), .A2(new_n854), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(new_n855), .Z(new_n911));
  XOR2_X1   g725(.A(new_n634), .B(KEYINPUT57), .Z(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n736), .B(KEYINPUT116), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n900), .A2(G469), .A3(new_n776), .A4(new_n775), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  INV_X1    g732(.A(new_n518), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n907), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(KEYINPUT117), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(KEYINPUT117), .B2(new_n921), .ZN(G60));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n652), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n907), .B1(new_n911), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n859), .A2(new_n927), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n924), .B(new_n929), .C1(new_n930), .C2(new_n652), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n652), .B1(new_n859), .B2(new_n927), .ZN(new_n932));
  INV_X1    g746(.A(new_n929), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT118), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT119), .B1(new_n910), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n940), .B(new_n937), .C1(new_n851), .C2(new_n854), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n673), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n853), .A2(new_n840), .A3(new_n812), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n844), .B2(new_n838), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n940), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n910), .A2(KEYINPUT119), .A3(new_n938), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n370), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n907), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n942), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n939), .A2(new_n941), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n370), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n946), .A2(new_n953), .A3(new_n370), .A4(new_n947), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n942), .A2(KEYINPUT61), .A3(new_n949), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT121), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n948), .A2(KEYINPUT120), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n956), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT121), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n952), .B1(new_n961), .B2(new_n965), .ZN(G66));
  NAND2_X1  g780(.A1(new_n825), .A2(new_n837), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n359), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT122), .Z(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n284), .B2(new_n530), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT123), .ZN(new_n972));
  INV_X1    g786(.A(G898), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n902), .B1(new_n973), .B2(G953), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  XNOR2_X1  g789(.A(new_n433), .B(new_n514), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n786), .A2(new_n647), .A3(new_n714), .A4(new_n768), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n796), .A2(new_n977), .A3(new_n800), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n732), .A2(new_n802), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT124), .Z(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n813), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n359), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n616), .A2(G900), .A3(G953), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n721), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n707), .A2(new_n472), .A3(new_n762), .A4(new_n820), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n800), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n987), .A2(new_n989), .A3(new_n796), .A4(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n985), .B1(new_n991), .B2(G953), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n984), .B1(new_n976), .B2(new_n992), .ZN(G72));
  NOR3_X1   g807(.A1(new_n978), .A2(new_n967), .A3(new_n981), .ZN(new_n994));
  XNOR2_X1  g808(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT126), .Z(new_n998));
  NOR2_X1   g812(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n434), .B(KEYINPUT127), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n999), .A2(new_n414), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n414), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n991), .A2(new_n967), .ZN(new_n1003));
  INV_X1    g817(.A(new_n998), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n997), .B1(new_n435), .B2(new_n716), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n847), .A2(new_n1006), .ZN(new_n1007));
  NOR4_X1   g821(.A1(new_n1001), .A2(new_n1005), .A3(new_n907), .A4(new_n1007), .ZN(G57));
endmodule


