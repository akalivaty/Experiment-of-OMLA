//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  AND2_X1   g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n203));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OR3_X1    g006(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT99), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n209), .B2(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G43gat), .B(G50gat), .Z(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n212), .B(KEYINPUT100), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(new_n206), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI22_X1  g020(.A1(new_n213), .A2(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT105), .A2(G85gat), .A3(G92gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  NAND2_X1  g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230));
  INV_X1    g029(.A(G85gat), .ZN(new_n231));
  INV_X1    g030(.A(G92gat), .ZN(new_n232));
  AOI22_X1  g031(.A1(KEYINPUT8), .A2(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G99gat), .B(G106gat), .Z(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(new_n225), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT106), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n236), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n222), .A2(new_n240), .B1(KEYINPUT41), .B2(new_n202), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G134gat), .B(G162gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n245), .A3(new_n241), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n205), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n205), .A3(new_n246), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G8gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(G15gat), .B(G22gat), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n252), .A2(G1gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT101), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT16), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n252), .B1(new_n256), .B2(G1gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n258), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT103), .ZN(new_n263));
  INV_X1    g062(.A(G64gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G57gat), .ZN(new_n265));
  INV_X1    g064(.A(G57gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G64gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G71gat), .B(G78gat), .Z(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT104), .B(G57gat), .Z(new_n272));
  OAI21_X1  g071(.A(new_n265), .B1(new_n272), .B2(new_n264), .ZN(new_n273));
  INV_X1    g072(.A(new_n270), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n263), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n261), .B1(KEYINPUT21), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G183gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n279));
  NAND2_X1  g078(.A1(G231gat), .A2(G233gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n278), .B(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n276), .A2(KEYINPUT21), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G155gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n282), .A2(new_n287), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n250), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n240), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT107), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n271), .A2(new_n275), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(new_n236), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n293), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n276), .A2(new_n240), .A3(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G230gat), .A2(G233gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n297), .A2(new_n302), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(G176gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(G204gat), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT108), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n308), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n292), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT109), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n224), .A2(new_n259), .A3(new_n260), .A4(new_n225), .ZN(new_n319));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n222), .A2(new_n261), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n319), .A2(KEYINPUT18), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT102), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT18), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n222), .B(new_n261), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n320), .B(KEYINPUT13), .Z(new_n328));
  AOI22_X1  g127(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G169gat), .B(G197gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G141gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT98), .B(KEYINPUT11), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT12), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n324), .A2(new_n329), .A3(new_n336), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G120gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G120gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(G113gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n347));
  INV_X1    g146(.A(G113gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G120gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n343), .A2(new_n345), .A3(new_n350), .A4(G113gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n342), .A2(G113gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT71), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n363));
  AOI211_X1 g162(.A(new_n363), .B(new_n360), .C1(new_n352), .C2(new_n356), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT24), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n366), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  INV_X1    g166(.A(G183gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G183gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n367), .B1(new_n372), .B2(KEYINPUT24), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT64), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT65), .ZN(new_n375));
  INV_X1    g174(.A(G169gat), .ZN(new_n376));
  INV_X1    g175(.A(G176gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT23), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(G169gat), .B2(G176gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n373), .A2(new_n374), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n366), .A2(G183gat), .A3(G190gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G183gat), .B(G190gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n366), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT25), .B1(new_n386), .B2(KEYINPUT64), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n382), .A2(new_n375), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(KEYINPUT68), .A2(G169gat), .A3(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n390), .A2(new_n391), .B1(G169gat), .B2(G176gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT26), .B1(new_n393), .B2(KEYINPUT68), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n392), .A2(new_n394), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n368), .A2(KEYINPUT27), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT27), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G183gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n398), .A3(new_n370), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT66), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT67), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(KEYINPUT67), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT28), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT67), .B1(new_n399), .B2(KEYINPUT66), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n395), .B(new_n403), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT25), .B1(new_n386), .B2(new_n382), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n389), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT72), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n365), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n357), .A2(KEYINPUT71), .A3(new_n361), .ZN(new_n412));
  INV_X1    g211(.A(new_n349), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n346), .B2(KEYINPUT70), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n355), .B1(new_n414), .B2(new_n351), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n363), .B1(new_n415), .B2(new_n360), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n389), .A2(new_n407), .A3(new_n408), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT72), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n411), .A2(new_n419), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT74), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n422), .B2(new_n423), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT32), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n419), .A3(new_n421), .ZN(new_n429));
  INV_X1    g228(.A(new_n420), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT33), .B1(new_n429), .B2(new_n430), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT73), .B(G71gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(G99gat), .ZN(new_n434));
  XOR2_X1   g233(.A(G15gat), .B(G43gat), .Z(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  AOI221_X4 g237(.A(new_n428), .B1(KEYINPUT33), .B2(new_n436), .C1(new_n429), .C2(new_n430), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n427), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT78), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n431), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n429), .A2(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n446), .A3(new_n436), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(new_n437), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(KEYINPUT78), .A3(new_n427), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n425), .A2(new_n426), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n451), .A3(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT77), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT77), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n447), .A2(new_n451), .A3(new_n454), .A4(new_n448), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n442), .A2(new_n450), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OR2_X1    g255(.A1(G197gat), .A2(G204gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(G197gat), .A2(G204gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT22), .ZN(new_n459));
  NAND2_X1  g258(.A1(G211gat), .A2(G218gat), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n457), .A2(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G218gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n286), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n460), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(KEYINPUT79), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(KEYINPUT79), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT79), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n468), .A3(new_n460), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n469), .A3(new_n461), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G226gat), .ZN(new_n472));
  INV_X1    g271(.A(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n418), .A2(KEYINPUT80), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n389), .A2(new_n407), .A3(new_n477), .A4(new_n408), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n474), .A2(KEYINPUT29), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n409), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n471), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n409), .A2(new_n474), .ZN(new_n484));
  INV_X1    g283(.A(new_n471), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n478), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n481), .ZN(new_n487));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G92gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT81), .B(G64gat), .ZN(new_n490));
  XOR2_X1   g289(.A(new_n489), .B(new_n490), .Z(new_n491));
  NAND4_X1  g290(.A1(new_n483), .A2(new_n487), .A3(KEYINPUT30), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n487), .ZN(new_n493));
  INV_X1    g292(.A(new_n491), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n492), .A2(KEYINPUT82), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n483), .A2(new_n487), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT30), .A4(new_n491), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n487), .A3(new_n491), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n503));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n506));
  NAND2_X1  g305(.A1(G155gat), .A2(G162gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(G155gat), .A2(G162gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(KEYINPUT2), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT84), .ZN(new_n512));
  XNOR2_X1  g311(.A(G141gat), .B(G148gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G155gat), .B(G162gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n507), .B2(KEYINPUT2), .ZN(new_n517));
  INV_X1    g316(.A(G148gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(G141gat), .ZN(new_n519));
  INV_X1    g318(.A(G141gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(G148gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n515), .B(new_n517), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n506), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n357), .B2(new_n361), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT85), .B(KEYINPUT3), .Z(new_n525));
  NAND3_X1  g324(.A1(new_n514), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n514), .A2(new_n522), .A3(new_n528), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI211_X1 g329(.A(KEYINPUT5), .B(new_n505), .C1(new_n524), .C2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n514), .A2(new_n522), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n412), .A2(new_n416), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n357), .A2(new_n361), .A3(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n530), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n532), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n504), .A3(new_n542), .ZN(new_n543));
  AND4_X1   g342(.A1(KEYINPUT4), .A2(new_n412), .A3(new_n416), .A4(new_n533), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n505), .B1(new_n524), .B2(new_n530), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n412), .A2(new_n416), .A3(KEYINPUT4), .A4(new_n533), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT87), .A4(new_n542), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n514), .A2(new_n522), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n415), .B2(new_n360), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n505), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT5), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n504), .B1(new_n535), .B2(new_n551), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT5), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT88), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n539), .B1(new_n549), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561));
  XNOR2_X1  g360(.A(G1gat), .B(G29gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT0), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n266), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(new_n231), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(G57gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G85gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n561), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(G85gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n231), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT93), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n503), .B1(new_n560), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n545), .A2(new_n548), .B1(new_n558), .B2(new_n555), .ZN(new_n575));
  OAI211_X1 g374(.A(KEYINPUT96), .B(new_n572), .C1(new_n575), .C2(new_n539), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n549), .A2(new_n559), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT89), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n569), .A2(new_n570), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n538), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT89), .B1(new_n575), .B2(new_n582), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n577), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n560), .A2(new_n581), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT6), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n502), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT92), .B(G22gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G228gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT29), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n471), .B1(new_n530), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n466), .A2(new_n470), .A3(new_n595), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n533), .B1(new_n597), .B2(new_n525), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n506), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n594), .B1(new_n600), .B2(new_n550), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT29), .B1(new_n527), .B2(new_n529), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(new_n471), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n599), .A2(KEYINPUT91), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT91), .B1(new_n599), .B2(new_n603), .ZN(new_n605));
  XNOR2_X1  g404(.A(G78gat), .B(G106gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT31), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(G50gat), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  AND4_X1   g409(.A1(KEYINPUT91), .A2(new_n599), .A3(new_n603), .A4(new_n609), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n593), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(new_n609), .ZN(new_n613));
  INV_X1    g412(.A(new_n604), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n592), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n456), .A2(new_n591), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT35), .ZN(new_n620));
  INV_X1    g419(.A(new_n590), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n589), .B1(new_n622), .B2(KEYINPUT90), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT90), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n584), .A2(new_n585), .A3(new_n624), .A4(new_n586), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT83), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT83), .B1(new_n495), .B2(new_n498), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n501), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n438), .A2(new_n439), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n631), .A2(new_n451), .B1(new_n617), .B2(new_n612), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n440), .A2(KEYINPUT76), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT76), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n449), .A2(new_n634), .A3(new_n427), .ZN(new_n635));
  AND4_X1   g434(.A1(KEYINPUT35), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n619), .A2(new_n620), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n633), .A2(KEYINPUT36), .A3(new_n452), .A4(new_n635), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n456), .B2(KEYINPUT36), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n552), .B2(new_n505), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n535), .A2(new_n551), .A3(KEYINPUT94), .A4(new_n504), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(KEYINPUT39), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n537), .A2(new_n541), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n505), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n641), .A2(KEYINPUT95), .A3(KEYINPUT39), .A4(new_n642), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n504), .B1(new_n537), .B2(new_n541), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n572), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n649), .A2(new_n652), .A3(KEYINPUT40), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT40), .B1(new_n649), .B2(new_n652), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n502), .A2(new_n655), .A3(new_n577), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n656), .A2(new_n618), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT37), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n658), .B(new_n494), .C1(new_n496), .C2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n483), .B2(new_n487), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT97), .B1(new_n661), .B2(new_n491), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n496), .A2(new_n659), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT38), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n485), .B1(new_n479), .B2(new_n482), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n484), .B(new_n471), .C1(new_n486), .C2(new_n481), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(KEYINPUT37), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n491), .A2(KEYINPUT38), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n670), .A2(new_n499), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n665), .A2(new_n588), .A3(new_n671), .A4(new_n590), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n618), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n626), .B2(new_n629), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n639), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n341), .B1(new_n637), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n318), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n626), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n502), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(G8gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n684), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n685), .A2(KEYINPUT110), .A3(new_n686), .A4(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1325gat));
  INV_X1    g491(.A(new_n639), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n456), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n694), .A2(G15gat), .B1(new_n678), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT111), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n674), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(new_n316), .ZN(new_n702));
  INV_X1    g501(.A(new_n250), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n702), .A2(new_n290), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n677), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n626), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n705), .A2(G29gat), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT45), .Z(new_n708));
  NOR3_X1   g507(.A1(new_n702), .A2(new_n341), .A3(new_n290), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n637), .A2(new_n676), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n250), .ZN(new_n712));
  AOI211_X1 g511(.A(KEYINPUT44), .B(new_n703), .C1(new_n637), .C2(new_n676), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n706), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n708), .A2(new_n715), .ZN(G1328gat));
  INV_X1    g515(.A(new_n502), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n705), .A2(G36gat), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(G36gat), .B1(new_n714), .B2(new_n717), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1329gat));
  OAI21_X1  g520(.A(G43gat), .B1(new_n714), .B2(new_n639), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n695), .A2(G43gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n705), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g524(.A(G50gat), .B1(new_n714), .B2(new_n618), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n618), .A2(G50gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n705), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g528(.A1(new_n292), .A2(new_n341), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n316), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n626), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(new_n272), .ZN(G1332gat));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n717), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  NOR3_X1   g539(.A1(new_n732), .A2(G71gat), .A3(new_n695), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n733), .A2(new_n693), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(G71gat), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n733), .A2(new_n674), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g545(.A(new_n703), .B1(new_n637), .B2(new_n676), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n340), .A2(new_n290), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(KEYINPUT51), .A3(new_n748), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n316), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n231), .A3(new_n626), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n316), .A2(new_n340), .A3(new_n290), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n712), .B2(new_n713), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT112), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n758), .B(new_n755), .C1(new_n712), .C2(new_n713), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n757), .A2(new_n626), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n754), .B1(new_n760), .B2(new_n231), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n756), .B2(new_n717), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n751), .A2(new_n752), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n316), .A2(G92gat), .A3(new_n717), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n764), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n757), .A2(new_n502), .A3(new_n759), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n770), .A2(KEYINPUT114), .A3(G92gat), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT114), .B1(new_n770), .B2(G92gat), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n773));
  AND2_X1   g572(.A1(new_n749), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n752), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n766), .B(KEYINPUT115), .Z(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n771), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n769), .B1(new_n779), .B2(new_n768), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n757), .A2(new_n693), .A3(new_n759), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G99gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n316), .A2(new_n695), .A3(G99gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT117), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1338gat));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(G106gat), .B1(new_n756), .B2(new_n618), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n618), .A2(G106gat), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n753), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n753), .B2(new_n790), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n787), .B(new_n788), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n757), .A2(new_n674), .A3(new_n759), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n702), .B(new_n790), .C1(new_n774), .C2(new_n775), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n795), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n793), .B1(new_n800), .B2(new_n787), .ZN(G1339gat));
  NAND4_X1  g600(.A1(new_n299), .A2(G230gat), .A3(G233gat), .A4(new_n300), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n303), .A2(KEYINPUT54), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n301), .A2(new_n804), .A3(new_n302), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n803), .A2(KEYINPUT55), .A3(new_n308), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n309), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n803), .A2(new_n308), .A3(new_n805), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n309), .A3(KEYINPUT120), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n809), .A2(new_n340), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n327), .A2(new_n328), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n335), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n339), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n314), .A2(new_n315), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n250), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n250), .A2(new_n818), .ZN(new_n821));
  INV_X1    g620(.A(new_n809), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n813), .A2(new_n812), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n291), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n702), .B2(new_n730), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n695), .A2(new_n674), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n706), .A2(new_n502), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n348), .A3(new_n341), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n828), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n340), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n834), .B2(new_n348), .ZN(G1340gat));
  NAND4_X1  g634(.A1(new_n833), .A2(new_n343), .A3(new_n345), .A4(new_n702), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n829), .B2(new_n316), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n839), .A3(new_n290), .ZN(new_n840));
  OAI21_X1  g639(.A(G127gat), .B1(new_n829), .B2(new_n291), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1342gat));
  INV_X1    g641(.A(G134gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n833), .A2(new_n843), .A3(new_n250), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n829), .B2(new_n703), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n826), .A2(new_n674), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n828), .A2(new_n639), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n520), .A3(new_n340), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n849), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n340), .A2(new_n812), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n819), .B1(new_n807), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n703), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n290), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n730), .A2(new_n702), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n674), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n852), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n341), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n856), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n858), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n870), .B(new_n856), .C1(new_n857), .C2(new_n849), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n518), .A3(new_n702), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n318), .A2(new_n341), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n859), .B(new_n674), .C1(new_n877), .C2(new_n865), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n850), .A2(KEYINPUT57), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n702), .A3(new_n853), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n860), .A2(new_n868), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT59), .B(new_n518), .C1(new_n883), .C2(new_n702), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n875), .B1(new_n882), .B2(new_n884), .ZN(G1345gat));
  NAND2_X1  g684(.A1(new_n290), .A2(G155gat), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT122), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(G155gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n854), .B2(new_n291), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n888), .A2(KEYINPUT123), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n869), .B2(new_n703), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n703), .A2(G162gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n854), .B2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n626), .A2(new_n717), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n814), .A2(new_n819), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n703), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n290), .B1(new_n901), .B2(new_n864), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n827), .B(new_n899), .C1(new_n902), .C2(new_n866), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n826), .A2(new_n905), .A3(new_n827), .A4(new_n899), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(new_n376), .A3(new_n341), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n826), .A2(new_n899), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n832), .ZN(new_n910));
  AOI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n340), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n908), .A2(new_n911), .ZN(G1348gat));
  OAI21_X1  g711(.A(G176gat), .B1(new_n907), .B2(new_n316), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n377), .A3(new_n702), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  NAND3_X1  g714(.A1(new_n904), .A2(new_n290), .A3(new_n906), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n290), .A2(new_n396), .A3(new_n398), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n916), .A2(G183gat), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n370), .A3(new_n250), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n250), .A3(new_n906), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(G190gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n924), .B2(G190gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT126), .B(new_n923), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1351gat));
  NAND2_X1  g731(.A1(new_n639), .A2(new_n899), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n850), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n340), .ZN(new_n935));
  INV_X1    g734(.A(new_n933), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n878), .A2(new_n879), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n340), .A2(G197gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  XOR2_X1   g739(.A(KEYINPUT127), .B(G204gat), .Z(new_n941));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n702), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT62), .Z(new_n943));
  AND3_X1   g742(.A1(new_n880), .A2(new_n702), .A3(new_n936), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n941), .B2(new_n944), .ZN(G1353gat));
  NAND3_X1  g744(.A1(new_n934), .A2(new_n286), .A3(new_n290), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n938), .A2(new_n290), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n948));
  OAI211_X1 g747(.A(KEYINPUT63), .B(G211gat), .C1(new_n937), .C2(new_n291), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n948), .B2(new_n950), .ZN(G1354gat));
  AOI21_X1  g750(.A(G218gat), .B1(new_n934), .B2(new_n250), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n703), .A2(new_n463), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n938), .B2(new_n953), .ZN(G1355gat));
endmodule


