//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n206), .C1(new_n202), .C2(new_n203), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT15), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT96), .B1(new_n209), .B2(G50gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n207), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n212), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n208), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT17), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n220), .B(KEYINPUT98), .C1(G1gat), .C2(new_n218), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G8gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT99), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G8gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n221), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT99), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT97), .B(KEYINPUT17), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n217), .A2(new_n224), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n216), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n222), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n233), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n216), .B(new_n226), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n231), .B(KEYINPUT13), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT95), .ZN(new_n242));
  XOR2_X1   g041(.A(G113gat), .B(G141gat), .Z(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT94), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n245));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n244), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(KEYINPUT95), .A3(new_n249), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT23), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n255), .A2(G169gat), .A3(G176gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G169gat), .ZN(new_n260));
  INV_X1    g059(.A(G176gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT23), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(KEYINPUT65), .A3(new_n257), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT25), .B1(new_n265), .B2(KEYINPUT23), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT24), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT24), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(G183gat), .A3(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G183gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n266), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n264), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n275), .A2(new_n273), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n255), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n262), .A2(new_n287), .A3(new_n257), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n280), .A2(new_n282), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n265), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n257), .B1(new_n293), .B2(KEYINPUT26), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n267), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n275), .A2(KEYINPUT27), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n274), .B(new_n276), .C1(new_n299), .C2(KEYINPUT68), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n275), .A2(KEYINPUT27), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n298), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n274), .A2(new_n276), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n307), .A2(KEYINPUT28), .A3(new_n303), .A4(new_n304), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n297), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n292), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G197gat), .B(G204gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT22), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n289), .B1(new_n279), .B2(KEYINPUT67), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n309), .B1(new_n321), .B2(new_n282), .ZN(new_n322));
  INV_X1    g121(.A(new_n292), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT29), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n311), .B(new_n320), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n264), .A2(new_n278), .A3(new_n281), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n281), .B1(new_n264), .B2(new_n278), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n328), .A2(new_n329), .A3(new_n289), .ZN(new_n330));
  OAI22_X1  g129(.A1(new_n330), .A2(new_n309), .B1(KEYINPUT29), .B2(new_n323), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n331), .A2(KEYINPUT76), .A3(new_n320), .A4(new_n311), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n311), .B1(new_n322), .B2(new_n324), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n319), .B(KEYINPUT75), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G8gat), .B(G36gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(G64gat), .ZN(new_n337));
  INV_X1    g136(.A(G92gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n327), .A2(new_n332), .A3(new_n335), .A4(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n325), .A2(new_n326), .B1(new_n333), .B2(new_n334), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n343), .A2(KEYINPUT30), .A3(new_n332), .A4(new_n339), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n332), .A3(new_n335), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(KEYINPUT77), .A3(new_n332), .ZN(new_n350));
  INV_X1    g149(.A(new_n339), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n353));
  AND2_X1   g152(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n354));
  AND2_X1   g153(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n356));
  OAI22_X1  g155(.A1(new_n353), .A2(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT2), .ZN(new_n358));
  INV_X1    g157(.A(G141gat), .ZN(new_n359));
  INV_X1    g158(.A(G148gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G162gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G155gat), .ZN(new_n363));
  INV_X1    g162(.A(G155gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G162gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n361), .A2(new_n363), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n361), .A3(new_n366), .ZN(new_n372));
  XNOR2_X1  g171(.A(G155gat), .B(G162gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n369), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n367), .B1(KEYINPUT2), .B2(new_n357), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n361), .A2(new_n366), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n378), .B2(new_n371), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G113gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT69), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G113gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n384), .A3(G120gat), .ZN(new_n385));
  INV_X1    g184(.A(G120gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G113gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G134gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G127gat), .ZN(new_n390));
  INV_X1    g189(.A(G127gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G134gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n392), .ZN(new_n397));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(KEYINPUT1), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n376), .A2(new_n380), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n369), .A2(new_n375), .A3(new_n396), .A4(new_n399), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT70), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n394), .B1(new_n387), .B2(new_n385), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n381), .A2(G120gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n408), .A2(new_n393), .B1(new_n390), .B2(new_n392), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n405), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n358), .A2(new_n368), .B1(new_n372), .B2(new_n374), .ZN(new_n411));
  INV_X1    g210(.A(new_n387), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT69), .B(G113gat), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(G120gat), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT70), .B(new_n399), .C1(new_n414), .C2(new_n394), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT4), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n401), .A2(new_n404), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  OAI22_X1  g217(.A1(new_n377), .A2(new_n379), .B1(new_n406), .B2(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n417), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT81), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n423), .B(new_n417), .C1(new_n402), .C2(new_n419), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT5), .B(new_n418), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G57gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G85gat), .ZN(new_n429));
  INV_X1    g228(.A(G57gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n427), .B(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G85gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n410), .A2(new_n411), .A3(new_n403), .A4(new_n415), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n417), .A4(new_n401), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n435), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n441), .A2(KEYINPUT83), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT83), .B1(new_n441), .B2(new_n442), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n435), .B1(new_n425), .B2(new_n440), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n440), .ZN(new_n447));
  INV_X1    g246(.A(new_n442), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n434), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(KEYINPUT84), .A3(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n346), .B(new_n352), .C1(new_n446), .C2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT31), .ZN(new_n456));
  INV_X1    g255(.A(G50gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT85), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n376), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n334), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n370), .B1(new_n319), .B2(KEYINPUT29), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n369), .A2(new_n375), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n462), .A2(G228gat), .A3(G233gat), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n319), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G228gat), .ZN(new_n469));
  INV_X1    g268(.A(G233gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT86), .B(G22gat), .Z(new_n472));
  AND3_X1   g271(.A1(new_n466), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n466), .B2(new_n471), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n459), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n466), .A2(new_n471), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G22gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n466), .A2(new_n471), .A3(new_n478), .A4(new_n472), .ZN(new_n479));
  INV_X1    g278(.A(new_n458), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n473), .A2(new_n478), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n454), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n410), .A2(new_n415), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n330), .A2(new_n488), .A3(new_n309), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n291), .B2(new_n310), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G227gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(new_n470), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT34), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n495));
  OAI221_X1 g294(.A(new_n495), .B1(new_n492), .B2(new_n470), .C1(new_n489), .C2(new_n490), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G99gat), .ZN(new_n498));
  XOR2_X1   g297(.A(G15gat), .B(G43gat), .Z(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n500));
  INV_X1    g299(.A(G71gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G43gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n500), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n498), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n500), .A2(new_n504), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G71gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(G99gat), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n511), .A3(KEYINPUT72), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(KEYINPUT33), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n511), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n488), .B1(new_n330), .B2(new_n309), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n322), .A2(new_n487), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n493), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n517), .A2(KEYINPUT32), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT32), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT33), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n514), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n497), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n524), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n522), .B1(new_n513), .B2(new_n516), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n520), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n526), .A2(new_n528), .B1(new_n494), .B2(new_n496), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n486), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n494), .A2(new_n496), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n528), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(KEYINPUT73), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n523), .ZN(new_n536));
  INV_X1    g335(.A(new_n514), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n536), .A2(new_n537), .B1(new_n527), .B2(new_n520), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n538), .A2(new_n497), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT36), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(KEYINPUT74), .B(new_n486), .C1(new_n525), .C2(new_n529), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n532), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n334), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n331), .A2(new_n311), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n320), .B1(new_n331), .B2(new_n311), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(KEYINPUT89), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n333), .A2(KEYINPUT89), .A3(new_n319), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT37), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT38), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n327), .A2(new_n552), .A3(new_n335), .A4(new_n332), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n351), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT90), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n553), .A2(new_n351), .ZN(new_n556));
  AOI211_X1 g355(.A(new_n323), .B(new_n309), .C1(new_n321), .C2(new_n282), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n324), .B1(new_n291), .B2(new_n310), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n319), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n548), .A3(new_n545), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT38), .B1(new_n562), .B2(KEYINPUT37), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n555), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n349), .A2(KEYINPUT37), .A3(new_n350), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n551), .B1(new_n567), .B2(new_n556), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT91), .ZN(new_n569));
  AND4_X1   g368(.A1(KEYINPUT84), .A2(new_n447), .A3(new_n448), .A4(new_n434), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT84), .B1(new_n445), .B2(new_n448), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n451), .A2(KEYINPUT91), .A3(new_n452), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n441), .A2(new_n442), .ZN(new_n574));
  INV_X1    g373(.A(new_n445), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n327), .A2(new_n332), .A3(new_n335), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n339), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n566), .A2(new_n568), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n347), .A2(new_n348), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT77), .B1(new_n343), .B2(new_n332), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n345), .B1(new_n582), .B2(new_n351), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n417), .B1(new_n438), .B2(new_n401), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT39), .B1(new_n420), .B2(new_n421), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n589), .B2(new_n435), .ZN(new_n590));
  AOI211_X1 g389(.A(KEYINPUT88), .B(new_n434), .C1(new_n584), .C2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g393(.A(KEYINPUT40), .B(new_n586), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n575), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n483), .B1(new_n583), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n485), .B(new_n543), .C1(new_n579), .C2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n346), .A2(new_n483), .A3(new_n352), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n525), .B2(new_n529), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n534), .A2(new_n497), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n533), .A2(new_n538), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT92), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT35), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n574), .A2(new_n575), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n572), .A2(new_n573), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n599), .A2(new_n605), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n483), .B1(new_n535), .B2(new_n540), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT35), .B1(new_n454), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n253), .B1(new_n598), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT102), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n430), .A2(G64gat), .ZN(new_n622));
  INV_X1    g421(.A(G64gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(G57gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n625), .B2(KEYINPUT100), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(KEYINPUT100), .B2(new_n625), .ZN(new_n627));
  XOR2_X1   g426(.A(G71gat), .B(G78gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n624), .A2(KEYINPUT101), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(KEYINPUT101), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n622), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n628), .A2(new_n621), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n629), .A2(new_n634), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n226), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT103), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n644), .A3(new_n226), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n639), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n639), .B1(new_n645), .B2(new_n643), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n620), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(new_n645), .ZN(new_n649));
  INV_X1    g448(.A(new_n639), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n639), .A2(new_n643), .A3(new_n645), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(new_n619), .ZN(new_n653));
  XNOR2_X1  g452(.A(G134gat), .B(G162gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G99gat), .B(G106gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n432), .A2(new_n338), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT7), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT105), .B(G92gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(G99gat), .A2(G106gat), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n661), .A2(new_n432), .B1(KEYINPUT8), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n656), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n660), .A2(new_n656), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(G232gat), .A2(G233gat), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n232), .A2(new_n668), .B1(KEYINPUT41), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n217), .A2(new_n229), .A3(new_n667), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n655), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n669), .A2(KEYINPUT41), .ZN(new_n674));
  XNOR2_X1  g473(.A(G190gat), .B(G218gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n671), .A3(new_n655), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n676), .ZN(new_n679));
  INV_X1    g478(.A(new_n677), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n672), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n648), .A2(new_n653), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n640), .A2(new_n666), .A3(new_n665), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n635), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT10), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n668), .A2(KEYINPUT10), .A3(new_n640), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G230gat), .A2(G233gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n690), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n687), .B2(new_n688), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n690), .B1(new_n684), .B2(new_n685), .ZN(new_n697));
  XNOR2_X1  g496(.A(G120gat), .B(G148gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G176gat), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(G204gat), .Z(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n693), .A2(new_n696), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n695), .B2(new_n697), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n683), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n613), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n446), .A2(new_n453), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G1gat), .ZN(G1324gat));
  INV_X1    g510(.A(new_n583), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT16), .B(G8gat), .Z(new_n713));
  NAND4_X1  g512(.A1(new_n708), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n712), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n707), .B2(new_n583), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n715), .A2(new_n717), .A3(new_n713), .ZN(new_n719));
  OAI221_X1 g518(.A(new_n714), .B1(new_n718), .B2(new_n225), .C1(KEYINPUT42), .C2(new_n719), .ZN(G1325gat));
  OAI21_X1  g519(.A(G15gat), .B1(new_n707), .B2(new_n543), .ZN(new_n721));
  INV_X1    g520(.A(new_n605), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(G15gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n707), .B2(new_n723), .ZN(G1326gat));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n483), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT43), .B(G22gat), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  NAND2_X1  g526(.A1(new_n648), .A2(new_n653), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n703), .A2(new_n704), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n678), .A2(new_n681), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT109), .Z(new_n734));
  NAND4_X1  g533(.A1(new_n613), .A2(new_n202), .A3(new_n709), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT45), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n241), .A2(KEYINPUT95), .A3(new_n249), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n249), .B1(new_n241), .B2(KEYINPUT95), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n251), .A2(KEYINPUT110), .A3(new_n252), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n731), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n732), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n746), .B(new_n748), .C1(new_n598), .C2(new_n612), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n556), .A2(new_n563), .A3(new_n564), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n564), .B1(new_n556), .B2(new_n563), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n578), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n568), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n597), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n543), .A2(new_n485), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n612), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n750), .B1(new_n757), .B2(new_n732), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n745), .B1(new_n749), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT112), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n761), .B(new_n745), .C1(new_n749), .C2(new_n758), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n760), .A2(new_n709), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n736), .B1(new_n763), .B2(new_n202), .ZN(G1328gat));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n712), .A3(new_n762), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT113), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n760), .A2(new_n767), .A3(new_n712), .A4(new_n762), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(G36gat), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n613), .A2(new_n203), .A3(new_n712), .A4(new_n734), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT46), .Z(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1329gat));
  AND2_X1   g571(.A1(new_n613), .A2(new_n734), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(new_n209), .A3(new_n605), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n543), .ZN(new_n776));
  NAND2_X1  g575(.A1(KEYINPUT47), .A2(G43gat), .ZN(new_n777));
  OAI221_X1 g576(.A(new_n774), .B1(new_n775), .B2(KEYINPUT47), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n774), .A2(new_n775), .ZN(new_n779));
  INV_X1    g578(.A(new_n543), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n780), .A3(new_n762), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(G43gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n778), .B1(new_n782), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g582(.A1(new_n760), .A2(new_n484), .A3(new_n762), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n483), .A2(G50gat), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n784), .A2(G50gat), .B1(new_n773), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n759), .A2(new_n483), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n457), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT48), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n786), .A2(KEYINPUT48), .B1(new_n788), .B2(new_n790), .ZN(G1331gat));
  AND3_X1   g590(.A1(new_n742), .A2(new_n683), .A3(new_n730), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n757), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n709), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n430), .ZN(G1332gat));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n712), .B1(new_n797), .B2(new_n623), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT115), .ZN(new_n800));
  NOR2_X1   g599(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1333gat));
  NOR3_X1   g601(.A1(new_n793), .A2(G71gat), .A3(new_n722), .ZN(new_n803));
  INV_X1    g602(.A(new_n793), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n780), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(G71gat), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n484), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g608(.A1(new_n743), .A2(new_n729), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n705), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n749), .B2(new_n758), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT116), .B(new_n812), .C1(new_n749), .C2(new_n758), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n816), .A2(new_n818), .A3(new_n794), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n746), .B1(new_n598), .B2(new_n612), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n820), .B2(new_n810), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n730), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n709), .A2(new_n432), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n819), .A2(new_n432), .B1(new_n824), .B2(new_n825), .ZN(G1336gat));
  INV_X1    g625(.A(new_n661), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n813), .B2(new_n583), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n583), .A2(G92gat), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n828), .B(new_n829), .C1(new_n824), .C2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n712), .A3(new_n817), .ZN(new_n833));
  INV_X1    g632(.A(new_n823), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n705), .B1(new_n834), .B2(new_n821), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n833), .A2(new_n827), .B1(new_n835), .B2(new_n830), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n829), .ZN(G1337gat));
  AOI21_X1  g636(.A(G99gat), .B1(new_n835), .B2(new_n605), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n816), .A2(new_n818), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n543), .A2(new_n498), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(G1338gat));
  OAI21_X1  g640(.A(G106gat), .B1(new_n813), .B2(new_n483), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n483), .A2(G106gat), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n842), .B(new_n843), .C1(new_n824), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n815), .A2(new_n484), .A3(new_n817), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n847), .A2(G106gat), .B1(new_n835), .B2(new_n844), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n843), .ZN(G1339gat));
  NAND3_X1  g648(.A1(new_n742), .A2(new_n683), .A3(new_n705), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT117), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n742), .A2(new_n683), .A3(new_n852), .A4(new_n705), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n688), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n687), .A2(new_n694), .A3(new_n688), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n700), .B1(new_n695), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n855), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n703), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n693), .A2(new_n696), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT55), .B(new_n862), .C1(new_n866), .C2(new_n859), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n865), .A2(new_n741), .A3(new_n740), .A4(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n236), .A2(new_n237), .A3(new_n240), .A4(new_n249), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n231), .B1(new_n230), .B2(new_n233), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n238), .A2(new_n239), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n248), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n705), .A2(KEYINPUT118), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  INV_X1    g674(.A(new_n873), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n730), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n732), .B1(new_n868), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n867), .A3(new_n703), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(new_n746), .A3(new_n873), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n728), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n854), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n722), .A2(new_n484), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n794), .A2(new_n712), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n253), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n885), .A2(KEYINPUT119), .A3(new_n886), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G113gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n599), .B1(new_n540), .B2(new_n535), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n794), .B(new_n894), .C1(new_n854), .C2(new_n882), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n413), .A3(new_n743), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(G1340gat));
  AOI21_X1  g696(.A(G120gat), .B1(new_n895), .B2(new_n730), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n889), .A2(new_n891), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n705), .A2(new_n386), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(G1341gat));
  NOR2_X1   g700(.A1(new_n728), .A2(new_n391), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n895), .A2(KEYINPUT120), .A3(new_n729), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT120), .B1(new_n895), .B2(new_n729), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(G127gat), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n899), .A2(new_n902), .B1(new_n903), .B2(new_n905), .ZN(G1342gat));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n732), .A3(new_n891), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G134gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n895), .A2(new_n389), .A3(new_n732), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(KEYINPUT121), .B2(KEYINPUT56), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(G1343gat));
  NOR3_X1   g713(.A1(new_n780), .A2(new_n483), .A3(new_n712), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n253), .A2(G141gat), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n883), .A2(new_n709), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n794), .B1(new_n854), .B2(new_n882), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n915), .A4(new_n916), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n886), .A2(new_n543), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n483), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n851), .A2(new_n853), .ZN(new_n928));
  INV_X1    g727(.A(new_n881), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n705), .B2(new_n873), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n876), .A2(KEYINPUT122), .A3(new_n730), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n931), .B(new_n932), .C1(new_n880), .C2(new_n253), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n934), .B2(new_n732), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n728), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n881), .B1(new_n933), .B2(new_n746), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n937), .A3(new_n729), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n927), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n483), .B1(new_n854), .B2(new_n882), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(KEYINPUT57), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n743), .B(new_n924), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n922), .B1(new_n945), .B2(G141gat), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT58), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n883), .A2(new_n484), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n925), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n939), .A2(new_n729), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n854), .B1(new_n950), .B2(KEYINPUT123), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n926), .B1(new_n951), .B2(new_n940), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n923), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n359), .B1(new_n953), .B2(new_n890), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT58), .B1(new_n917), .B2(KEYINPUT125), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(KEYINPUT125), .B2(new_n917), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n946), .A2(new_n947), .B1(new_n954), .B2(new_n956), .ZN(G1344gat));
  AND2_X1   g756(.A1(new_n919), .A2(new_n915), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n360), .A3(new_n730), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G148gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n961), .B1(new_n953), .B2(new_n730), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n948), .A2(KEYINPUT57), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n483), .A2(KEYINPUT57), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n706), .A2(new_n253), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n950), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n963), .A2(new_n730), .A3(new_n924), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n960), .B1(new_n967), .B2(G148gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n959), .B1(new_n962), .B2(new_n968), .ZN(G1345gat));
  OR2_X1    g768(.A1(new_n354), .A2(new_n353), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n958), .A2(new_n971), .A3(new_n729), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n953), .A2(new_n729), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n971), .ZN(G1346gat));
  OR2_X1    g773(.A1(new_n355), .A2(new_n356), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n976), .A3(new_n732), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n953), .A2(new_n732), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n976), .ZN(G1347gat));
  NOR2_X1   g778(.A1(new_n709), .A2(new_n583), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n885), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n981), .A2(new_n260), .A3(new_n253), .ZN(new_n982));
  INV_X1    g781(.A(new_n980), .ZN(new_n983));
  AOI211_X1 g782(.A(new_n610), .B(new_n983), .C1(new_n854), .C2(new_n882), .ZN(new_n984));
  AOI21_X1  g783(.A(G169gat), .B1(new_n984), .B2(new_n743), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n982), .A2(new_n985), .ZN(G1348gat));
  OAI21_X1  g785(.A(G176gat), .B1(new_n981), .B2(new_n705), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n984), .A2(new_n261), .A3(new_n730), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1349gat));
  NAND4_X1  g788(.A1(new_n883), .A2(new_n729), .A3(new_n884), .A4(new_n980), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n729), .A2(new_n303), .A3(new_n304), .ZN(new_n991));
  AOI22_X1  g790(.A1(G183gat), .A2(new_n990), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n992), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n993));
  NOR2_X1   g792(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n994));
  AND2_X1   g793(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n993), .A2(new_n996), .ZN(G1350gat));
  NAND3_X1  g796(.A1(new_n984), .A2(new_n307), .A3(new_n732), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n885), .A2(new_n732), .A3(new_n980), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n999), .A2(new_n1000), .A3(G190gat), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n1000), .B1(new_n999), .B2(G190gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(G1351gat));
  NOR2_X1   g802(.A1(new_n780), .A2(new_n983), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n943), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1005), .A2(new_n742), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n966), .B(new_n1004), .C1(new_n943), .C2(new_n925), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n890), .A2(G197gat), .ZN(new_n1008));
  OAI22_X1  g807(.A1(new_n1006), .A2(G197gat), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(G1352gat));
  NOR3_X1   g809(.A1(new_n1005), .A2(G204gat), .A3(new_n705), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT62), .ZN(new_n1012));
  OAI211_X1 g811(.A(new_n730), .B(new_n966), .C1(new_n943), .C2(new_n925), .ZN(new_n1013));
  INV_X1    g812(.A(new_n1004), .ZN(new_n1014));
  OR3_X1    g813(.A1(new_n1013), .A2(KEYINPUT127), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g814(.A(KEYINPUT127), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1015), .A2(G204gat), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1012), .A2(new_n1017), .ZN(G1353gat));
  NAND4_X1  g817(.A1(new_n963), .A2(new_n729), .A3(new_n966), .A4(new_n1004), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1019), .B2(G211gat), .ZN(new_n1020));
  OAI211_X1 g819(.A(KEYINPUT63), .B(G211gat), .C1(new_n1007), .C2(new_n728), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n729), .A2(new_n314), .ZN(new_n1023));
  OAI22_X1  g822(.A1(new_n1020), .A2(new_n1022), .B1(new_n1005), .B2(new_n1023), .ZN(G1354gat));
  OAI21_X1  g823(.A(new_n315), .B1(new_n1005), .B2(new_n746), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n732), .A2(G218gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1025), .B1(new_n1007), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g826(.A(new_n1027), .ZN(G1355gat));
endmodule


