//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(new_n454), .B(KEYINPUT69), .Z(G261));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(G2106), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(KEYINPUT3), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n462), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n472), .A2(G2105), .A3(new_n464), .A4(new_n465), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n466), .A2(new_n467), .A3(new_n472), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(G136), .B2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n467), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI22_X1  g069(.A1(new_n487), .A2(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n467), .A3(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n479), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n467), .A2(G138), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n472), .A2(new_n464), .A3(new_n465), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n495), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  OAI211_X1 g080(.A(KEYINPUT73), .B(G62), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(KEYINPUT74), .A2(G75), .A3(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(G75), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n503), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n519), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT72), .A3(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(new_n522), .B1(KEYINPUT6), .B2(new_n503), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n515), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G88), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(new_n522), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(G543), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n518), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n524), .A3(new_n528), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n527), .A2(G543), .A3(new_n528), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT75), .B(G51), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AND2_X1   g115(.A1(G63), .A2(G651), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n524), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n534), .A2(new_n537), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n533), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n524), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n535), .A2(G52), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n545), .A2(new_n550), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n533), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n535), .A2(G43), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n554), .B(new_n555), .C1(new_n503), .C2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G860), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n557), .A2(new_n558), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n529), .B2(new_n565), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n547), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n533), .A2(G91), .B1(new_n571), .B2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n574), .B1(new_n518), .B2(new_n530), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n535), .A2(G50), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n578), .A2(KEYINPUT77), .A3(new_n579), .A4(new_n525), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n575), .A2(new_n580), .ZN(G303));
  NAND2_X1  g156(.A1(new_n535), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n523), .A2(G87), .A3(new_n524), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  OAI21_X1  g160(.A(G61), .B1(new_n504), .B2(new_n505), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n503), .B1(new_n529), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n532), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n523), .A2(KEYINPUT78), .A3(G86), .A4(new_n524), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n524), .A2(G60), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n503), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT79), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n533), .A2(G85), .B1(new_n535), .B2(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n523), .A2(G92), .A3(new_n524), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT10), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT80), .B(G66), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n524), .A2(new_n607), .B1(G79), .B2(G543), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n503), .B1(new_n608), .B2(new_n609), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n610), .A2(new_n611), .B1(G54), .B2(new_n535), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n606), .A2(KEYINPUT82), .A3(new_n612), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n604), .B1(new_n617), .B2(new_n603), .ZN(G284));
  AOI21_X1  g193(.A(new_n604), .B1(new_n617), .B2(new_n603), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(G860), .B2(new_n624), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  MUX2_X1   g201(.A(new_n557), .B(new_n626), .S(G868), .Z(G323));
  XNOR2_X1  g202(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g203(.A(G323), .B(new_n628), .ZN(G282));
  NOR3_X1   g204(.A1(new_n474), .A2(G2105), .A3(new_n479), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n637));
  INV_X1    g212(.A(G123), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n466), .A2(new_n467), .A3(new_n472), .ZN(new_n639));
  INV_X1    g214(.A(G135), .ZN(new_n640));
  OAI221_X1 g215(.A(new_n637), .B1(new_n638), .B2(new_n487), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n635), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT88), .B(G2438), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2430), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT87), .B(KEYINPUT14), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n653), .B(new_n657), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(G14), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n659), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n632), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G2096), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n678), .A2(KEYINPUT90), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(KEYINPUT90), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n676), .A2(new_n677), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(new_n687), .B(new_n686), .S(new_n682), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G21), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G168), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G1966), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT102), .Z(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G11), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G28), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n702), .B2(G28), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n701), .B1(new_n703), .B2(new_n705), .C1(new_n641), .C2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(G26), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  OAI21_X1  g283(.A(KEYINPUT98), .B1(G104), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g285(.A1(KEYINPUT98), .A2(G104), .A3(G2105), .ZN(new_n711));
  OAI221_X1 g286(.A(G2104), .B1(G116), .B2(new_n467), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G128), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n487), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n490), .B2(G140), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n708), .B1(new_n715), .B2(new_n704), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT99), .B(G2067), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G2084), .ZN(new_n719));
  INV_X1    g294(.A(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n720), .B2(KEYINPUT24), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT24), .B2(new_n720), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n483), .B2(new_n704), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n706), .B(new_n718), .C1(new_n719), .C2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G27), .A2(G29), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G164), .B2(G29), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n716), .A2(new_n717), .B1(new_n726), .B2(G2078), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n700), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n723), .A2(new_n719), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n704), .A2(G33), .ZN(new_n731));
  NAND2_X1  g306(.A1(G115), .A2(G2104), .ZN(new_n732));
  INV_X1    g307(.A(G127), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n479), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2105), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  INV_X1    g312(.A(G139), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n737), .C1(new_n639), .C2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT100), .Z(new_n740));
  OAI21_X1  g315(.A(new_n731), .B1(new_n740), .B2(new_n704), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2072), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n728), .A2(new_n730), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n696), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n696), .ZN(new_n745));
  INV_X1    g320(.A(G1961), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G162), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT29), .B(G2090), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n704), .A2(G32), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n490), .A2(G141), .ZN(new_n754));
  INV_X1    g329(.A(new_n487), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G129), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n475), .A2(G105), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n754), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n753), .B1(new_n763), .B2(new_n704), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n764), .B(new_n765), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n696), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n698), .A2(G1966), .B1(G2078), .B2(new_n726), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n752), .A2(new_n766), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  MUX2_X1   g348(.A(G19), .B(new_n557), .S(G16), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G1341), .Z(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n617), .B2(G16), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1348), .Z(new_n779));
  NAND4_X1  g354(.A1(new_n743), .A2(new_n773), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(G288), .A2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G23), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(G16), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n696), .A2(G22), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT94), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n696), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1971), .ZN(new_n790));
  INV_X1    g365(.A(G1971), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(new_n788), .C1(G166), .C2(new_n696), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n781), .B(new_n784), .C1(G16), .C2(new_n782), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n786), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n696), .A2(G6), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n595), .B2(new_n696), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n795), .B(new_n797), .C1(new_n595), .C2(new_n696), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n600), .A2(G16), .A3(new_n601), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n808));
  OR2_X1    g383(.A1(G16), .A2(G24), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(new_n812));
  OAI21_X1  g387(.A(G1986), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n812), .ZN(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(new_n815), .A3(new_n810), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n704), .A2(G25), .ZN(new_n818));
  OR2_X1    g393(.A1(G95), .A2(G2105), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n819), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n820));
  INV_X1    g395(.A(G119), .ZN(new_n821));
  INV_X1    g396(.A(G131), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n820), .B1(new_n821), .B2(new_n487), .C1(new_n639), .C2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT91), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n487), .B2(new_n821), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n490), .B2(G131), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT91), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n818), .B1(new_n829), .B2(G29), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT35), .B(G1991), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n704), .B1(new_n825), .B2(new_n828), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n831), .B1(new_n834), .B2(new_n818), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(KEYINPUT92), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n817), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(new_n835), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n839), .A2(new_n840), .B1(new_n802), .B2(new_n803), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n806), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT92), .B1(new_n833), .B2(new_n835), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n794), .A2(KEYINPUT34), .A3(new_n801), .ZN(new_n844));
  NOR4_X1   g419(.A1(new_n837), .A2(KEYINPUT95), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n805), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(new_n805), .C1(new_n842), .C2(new_n845), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n780), .B1(new_n847), .B2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n849), .ZN(new_n851));
  INV_X1    g426(.A(new_n780), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT103), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  AOI211_X1 g429(.A(new_n854), .B(new_n780), .C1(new_n847), .C2(new_n849), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(G150));
  NAND2_X1  g431(.A1(new_n617), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n533), .A2(G93), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n535), .A2(G55), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n859), .B(new_n860), .C1(new_n503), .C2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n557), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n557), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n858), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  AOI21_X1  g442(.A(G860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n762), .B(new_n715), .ZN(new_n873));
  INV_X1    g448(.A(new_n495), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n875));
  INV_X1    g450(.A(new_n498), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(KEYINPUT104), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n495), .B2(new_n501), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(new_n881), .ZN(new_n883));
  INV_X1    g458(.A(new_n740), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n884), .A2(new_n885), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n755), .A2(G130), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n467), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(G142), .B2(new_n490), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n631), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n823), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n889), .A2(new_n898), .A3(new_n890), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n641), .B(G160), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(G162), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n904), .A3(new_n901), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n862), .A2(new_n603), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n626), .B(new_n865), .Z(new_n912));
  NAND3_X1  g487(.A1(new_n621), .A2(new_n606), .A3(new_n612), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n613), .A2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n915), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(G305), .ZN(new_n923));
  XNOR2_X1  g498(.A(G166), .B(G288), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT42), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  OAI221_X1 g503(.A(new_n921), .B1(new_n922), .B2(new_n912), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n921), .B1(new_n922), .B2(new_n912), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(KEYINPUT106), .A3(new_n926), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n929), .A2(new_n931), .B1(new_n928), .B2(new_n927), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n911), .B1(new_n932), .B2(new_n603), .ZN(G295));
  OAI21_X1  g508(.A(new_n911), .B1(new_n932), .B2(new_n603), .ZN(G331));
  XOR2_X1   g509(.A(G301), .B(KEYINPUT107), .Z(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n864), .A3(new_n863), .ZN(new_n936));
  XNOR2_X1  g511(.A(G301), .B(KEYINPUT107), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n865), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G168), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n938), .A3(G168), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n915), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n918), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n943), .A2(new_n945), .A3(new_n939), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n919), .A2(KEYINPUT108), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n942), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n925), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT109), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n922), .B1(new_n943), .B2(new_n939), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n940), .A2(new_n919), .A3(new_n941), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n908), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n940), .B(new_n941), .C1(new_n944), .C2(new_n918), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n952), .B1(new_n957), .B2(new_n947), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n925), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n951), .A2(new_n956), .A3(new_n960), .A4(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT44), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n951), .A2(new_n956), .A3(new_n960), .A4(new_n962), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n955), .B2(new_n963), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(G397));
  NOR2_X1   g547(.A1(new_n881), .A2(G1384), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n473), .A2(new_n476), .A3(new_n482), .A4(G40), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(G1996), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT111), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n763), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n715), .B(G2067), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n979), .B2(new_n763), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n975), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n829), .A2(new_n832), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n715), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n976), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G290), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n975), .A2(new_n815), .A3(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n827), .B(new_n831), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n975), .A2(new_n993), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n981), .A2(new_n992), .A3(new_n984), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n976), .B1(new_n763), .B2(new_n982), .ZN(new_n996));
  INV_X1    g571(.A(new_n978), .ZN(new_n997));
  INV_X1    g572(.A(new_n980), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(KEYINPUT46), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n978), .B2(new_n980), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n989), .B(new_n995), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n575), .A2(G8), .A3(new_n580), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n575), .A2(KEYINPUT55), .A3(G8), .A4(new_n580), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n495), .B2(new_n501), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n974), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1014));
  INV_X1    g589(.A(G2090), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(new_n1012), .C1(new_n495), .C2(new_n501), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n878), .A2(new_n880), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n974), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1971), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1011), .B(G8), .C1(new_n1019), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n582), .A2(G1976), .A3(new_n583), .A4(new_n584), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1027), .C1(new_n1013), .C2(new_n974), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(G288), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT113), .B(G1976), .Z(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1028), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT112), .B1(new_n1028), .B2(KEYINPUT52), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n593), .A2(new_n594), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n503), .B1(new_n586), .B2(new_n587), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n535), .B2(G48), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n532), .A2(new_n592), .ZN(new_n1045));
  OAI21_X1  g620(.A(G1981), .B1(new_n590), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(KEYINPUT49), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1046), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT114), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1013), .A2(new_n974), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AND4_X1   g630(.A1(new_n1047), .A2(new_n1049), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1038), .A2(new_n1056), .A3(KEYINPUT115), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1033), .B1(new_n1061), .B2(new_n1035), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1049), .A2(new_n1052), .A3(new_n1055), .A4(new_n1047), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1058), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1026), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g640(.A1(G288), .A2(G1976), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1043), .B1(new_n1056), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1052), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n791), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1018), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1074), .A3(G8), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1011), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1025), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1078));
  INV_X1    g653(.A(G1966), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1021), .B1(new_n495), .B2(new_n501), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1023), .B2(KEYINPUT117), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1082), .B(new_n974), .C1(new_n1013), .C2(new_n1020), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1079), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1014), .A2(new_n719), .A3(new_n1017), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1051), .B(G286), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1077), .A2(new_n1078), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1025), .A2(KEYINPUT63), .ZN(new_n1090));
  OAI21_X1  g665(.A(G8), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1076), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT115), .B1(new_n1038), .B2(new_n1056), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1062), .A2(new_n1058), .A3(new_n1063), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(new_n1086), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1069), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1084), .A2(G168), .A3(new_n1085), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  AOI21_X1  g674(.A(G168), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT51), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(new_n1103), .A3(G8), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1051), .B1(new_n1106), .B2(new_n1073), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1011), .B1(new_n1107), .B2(new_n1070), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1025), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT124), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1077), .A2(new_n1078), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G2078), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1022), .A2(new_n1023), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1117));
  INV_X1    g692(.A(new_n974), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1017), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n746), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(G2078), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1081), .A2(new_n1083), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G171), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1105), .A2(new_n1110), .A3(new_n1112), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1102), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1097), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1114), .A2(new_n1115), .B1(new_n746), .B2(new_n1119), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n974), .A2(new_n1123), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1022), .B(new_n1131), .C1(new_n973), .C2(KEYINPUT45), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1132), .A3(KEYINPUT125), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(G171), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(G301), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1130), .A2(new_n1132), .A3(G301), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1125), .A2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1137), .A2(new_n1140), .B1(new_n1142), .B2(new_n1138), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1145), .A2(KEYINPUT126), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G299), .B(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1119), .A2(new_n770), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(G2072), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1022), .A2(new_n1023), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT119), .ZN(new_n1154));
  XNOR2_X1  g729(.A(G299), .B(KEYINPUT57), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1022), .A2(new_n1023), .A3(new_n1151), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1956), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1050), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(G2067), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1348), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n617), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1154), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1022), .A2(new_n1023), .A3(new_n979), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1165), .A2(KEYINPUT120), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT58), .B(G1341), .Z(new_n1167));
  AOI22_X1  g742(.A1(new_n1165), .A2(KEYINPUT120), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n557), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1158), .A2(KEYINPUT61), .A3(new_n1153), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1169), .B2(KEYINPUT59), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT60), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(new_n615), .A3(new_n616), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1162), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1175), .A2(new_n1162), .A3(new_n1177), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1184), .B(new_n1155), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1182), .B1(new_n1154), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1173), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1145), .A2(KEYINPUT126), .B1(new_n1164), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1129), .B1(new_n1146), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n991), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n990), .A2(new_n815), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1191), .B1(new_n975), .B2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT110), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(new_n981), .A3(new_n984), .A4(new_n994), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1006), .B1(new_n1190), .B2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g771(.A(G227), .ZN(new_n1198));
  AND3_X1   g772(.A1(new_n1198), .A2(KEYINPUT127), .A3(G319), .ZN(new_n1199));
  AOI21_X1  g773(.A(KEYINPUT127), .B1(new_n1198), .B2(G319), .ZN(new_n1200));
  NOR4_X1   g774(.A1(G229), .A2(G401), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND3_X1  g775(.A1(new_n969), .A2(new_n909), .A3(new_n1201), .ZN(G225));
  INV_X1    g776(.A(G225), .ZN(G308));
endmodule


