

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748;

  AND2_X1 U374 ( .A1(n537), .A2(KEYINPUT83), .ZN(n556) );
  AND2_X1 U375 ( .A1(n594), .A2(n660), .ZN(n595) );
  NAND2_X1 U376 ( .A1(n599), .A2(n598), .ZN(n604) );
  INV_X1 U377 ( .A(G953), .ZN(n735) );
  NAND2_X1 U378 ( .A1(n548), .A2(n549), .ZN(n649) );
  XOR2_X1 U379 ( .A(n503), .B(n502), .Z(n352) );
  NAND2_X2 U380 ( .A1(n617), .A2(n616), .ZN(n389) );
  XNOR2_X2 U381 ( .A(KEYINPUT112), .B(n595), .ZN(n742) );
  NOR2_X2 U382 ( .A1(n613), .A2(n492), .ZN(n392) );
  XNOR2_X2 U383 ( .A(n590), .B(KEYINPUT38), .ZN(n673) );
  NOR2_X2 U384 ( .A1(n556), .A2(n555), .ZN(n562) );
  NOR2_X2 U385 ( .A1(n424), .A2(n585), .ZN(n423) );
  NOR2_X2 U386 ( .A1(n573), .A2(n677), .ZN(n575) );
  XNOR2_X2 U387 ( .A(n578), .B(KEYINPUT1), .ZN(n660) );
  NOR2_X1 U388 ( .A1(n589), .A2(n588), .ZN(n606) );
  XOR2_X2 U389 ( .A(G122), .B(G104), .Z(n482) );
  OR2_X1 U390 ( .A1(n645), .A2(n355), .ZN(n402) );
  NOR2_X1 U391 ( .A1(n747), .A2(n748), .ZN(n381) );
  NAND2_X1 U392 ( .A1(n400), .A2(n367), .ZN(n555) );
  XNOR2_X1 U393 ( .A(KEYINPUT35), .B(n542), .ZN(n745) );
  XNOR2_X1 U394 ( .A(KEYINPUT42), .B(n580), .ZN(n748) );
  AND2_X1 U395 ( .A1(n570), .A2(n412), .ZN(n411) );
  NOR2_X1 U396 ( .A1(n577), .A2(n672), .ZN(n393) );
  NAND2_X1 U397 ( .A1(n584), .A2(n414), .ZN(n412) );
  XNOR2_X1 U398 ( .A(n416), .B(n417), .ZN(n656) );
  NAND2_X1 U399 ( .A1(n372), .A2(n369), .ZN(n578) );
  OR2_X1 U400 ( .A1(n715), .A2(G902), .ZN(n416) );
  XOR2_X1 U401 ( .A(n715), .B(KEYINPUT125), .Z(n718) );
  AND2_X2 U402 ( .A1(n389), .A2(n707), .ZN(n716) );
  XNOR2_X1 U403 ( .A(n377), .B(n440), .ZN(n703) );
  NOR2_X2 U404 ( .A1(n614), .A2(n697), .ZN(n465) );
  XNOR2_X2 U405 ( .A(n519), .B(n518), .ZN(n377) );
  XNOR2_X1 U406 ( .A(n455), .B(n435), .ZN(n524) );
  INV_X1 U407 ( .A(G119), .ZN(n435) );
  XOR2_X1 U408 ( .A(G146), .B(KEYINPUT4), .Z(n516) );
  INV_X1 U409 ( .A(KEYINPUT84), .ZN(n405) );
  NAND2_X1 U410 ( .A1(n746), .A2(n642), .ZN(n364) );
  AND2_X1 U411 ( .A1(n368), .A2(n633), .ZN(n367) );
  XNOR2_X1 U412 ( .A(n551), .B(KEYINPUT102), .ZN(n368) );
  INV_X1 U413 ( .A(KEYINPUT67), .ZN(n383) );
  NAND2_X1 U414 ( .A1(G237), .A2(G234), .ZN(n469) );
  XNOR2_X1 U415 ( .A(KEYINPUT5), .B(KEYINPUT93), .ZN(n520) );
  XOR2_X1 U416 ( .A(KEYINPUT73), .B(KEYINPUT94), .Z(n521) );
  NOR2_X1 U417 ( .A1(G953), .A2(G237), .ZN(n522) );
  XOR2_X1 U418 ( .A(G125), .B(KEYINPUT76), .Z(n462) );
  XNOR2_X1 U419 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n458) );
  XOR2_X1 U420 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n459) );
  XNOR2_X1 U421 ( .A(n568), .B(KEYINPUT108), .ZN(n569) );
  NOR2_X1 U422 ( .A1(n567), .A2(n566), .ZN(n584) );
  INV_X1 U423 ( .A(KEYINPUT75), .ZN(n414) );
  XNOR2_X1 U424 ( .A(n512), .B(n513), .ZN(n417) );
  INV_X1 U425 ( .A(KEYINPUT90), .ZN(n513) );
  AND2_X1 U426 ( .A1(n374), .A2(n373), .ZN(n372) );
  OR2_X1 U427 ( .A1(n703), .A2(n370), .ZN(n369) );
  NAND2_X1 U428 ( .A1(G469), .A2(G902), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n524), .B(n434), .ZN(n727) );
  XNOR2_X1 U430 ( .A(n457), .B(n534), .ZN(n434) );
  XOR2_X1 U431 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n456) );
  XNOR2_X1 U432 ( .A(G122), .B(G116), .ZN(n445) );
  XOR2_X1 U433 ( .A(KEYINPUT9), .B(G107), .Z(n446) );
  XOR2_X1 U434 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n450) );
  XNOR2_X1 U435 ( .A(n545), .B(KEYINPUT95), .ZN(n669) );
  OR2_X1 U436 ( .A1(n569), .A2(n410), .ZN(n409) );
  OR2_X1 U437 ( .A1(n584), .A2(n414), .ZN(n410) );
  BUF_X1 U438 ( .A(n610), .Z(n394) );
  XNOR2_X1 U439 ( .A(G478), .B(n491), .ZN(n549) );
  XNOR2_X1 U440 ( .A(n498), .B(KEYINPUT70), .ZN(n430) );
  INV_X1 U441 ( .A(KEYINPUT22), .ZN(n498) );
  BUF_X1 U442 ( .A(n656), .Z(n399) );
  XNOR2_X1 U443 ( .A(n533), .B(n441), .ZN(n440) );
  XNOR2_X1 U444 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U445 ( .A(n534), .B(n357), .ZN(n441) );
  NOR2_X1 U446 ( .A1(G952), .A2(n735), .ZN(n719) );
  NAND2_X1 U447 ( .A1(n429), .A2(n707), .ZN(n428) );
  NOR2_X1 U448 ( .A1(n605), .A2(n421), .ZN(n418) );
  NAND2_X1 U449 ( .A1(n422), .A2(KEYINPUT72), .ZN(n421) );
  INV_X1 U450 ( .A(KEYINPUT47), .ZN(n422) );
  XOR2_X1 U451 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n494) );
  OR2_X1 U452 ( .A1(G902), .A2(G237), .ZN(n466) );
  NAND2_X1 U453 ( .A1(n439), .A2(n371), .ZN(n370) );
  INV_X1 U454 ( .A(G902), .ZN(n371) );
  XNOR2_X1 U455 ( .A(G140), .B(KEYINPUT10), .ZN(n475) );
  INV_X1 U456 ( .A(KEYINPUT48), .ZN(n378) );
  INV_X1 U457 ( .A(n584), .ZN(n425) );
  NAND2_X1 U458 ( .A1(n656), .A2(n576), .ZN(n585) );
  INV_X1 U459 ( .A(n409), .ZN(n388) );
  NAND2_X1 U460 ( .A1(n660), .A2(n661), .ZN(n544) );
  NOR2_X1 U461 ( .A1(n656), .A2(n657), .ZN(n661) );
  XNOR2_X1 U462 ( .A(n363), .B(n362), .ZN(n471) );
  INV_X1 U463 ( .A(KEYINPUT88), .ZN(n362) );
  AND2_X1 U464 ( .A1(n674), .A2(n576), .ZN(n496) );
  XNOR2_X1 U465 ( .A(n526), .B(n525), .ZN(n627) );
  XNOR2_X1 U466 ( .A(n377), .B(n354), .ZN(n526) );
  XOR2_X1 U467 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n503) );
  XNOR2_X1 U468 ( .A(KEYINPUT100), .B(KEYINPUT98), .ZN(n478) );
  XNOR2_X1 U469 ( .A(G143), .B(G113), .ZN(n476) );
  XOR2_X1 U470 ( .A(G107), .B(G110), .Z(n534) );
  INV_X1 U471 ( .A(G101), .ZN(n531) );
  XNOR2_X1 U472 ( .A(n431), .B(n727), .ZN(n697) );
  XNOR2_X1 U473 ( .A(n464), .B(n358), .ZN(n432) );
  XNOR2_X1 U474 ( .A(n386), .B(n385), .ZN(n571) );
  INV_X1 U475 ( .A(KEYINPUT39), .ZN(n385) );
  NAND2_X1 U476 ( .A1(n387), .A2(n356), .ZN(n386) );
  NOR2_X1 U477 ( .A1(n407), .A2(n388), .ZN(n387) );
  NAND2_X1 U478 ( .A1(n661), .A2(n578), .ZN(n568) );
  XNOR2_X1 U479 ( .A(n529), .B(KEYINPUT6), .ZN(n530) );
  INV_X1 U480 ( .A(KEYINPUT103), .ZN(n529) );
  XNOR2_X1 U481 ( .A(n395), .B(n449), .ZN(n452) );
  XNOR2_X1 U482 ( .A(n451), .B(n450), .ZN(n395) );
  XNOR2_X1 U483 ( .A(n406), .B(KEYINPUT40), .ZN(n747) );
  NOR2_X1 U484 ( .A1(n571), .A2(n649), .ZN(n406) );
  XNOR2_X1 U485 ( .A(n592), .B(n591), .ZN(n594) );
  AND2_X1 U486 ( .A1(n438), .A2(n437), .ZN(n542) );
  INV_X1 U487 ( .A(n581), .ZN(n437) );
  NOR2_X1 U488 ( .A1(n536), .A2(n391), .ZN(n390) );
  XNOR2_X1 U489 ( .A(n375), .B(n547), .ZN(n652) );
  NOR2_X1 U490 ( .A1(n394), .A2(n583), .ZN(n645) );
  AND2_X1 U491 ( .A1(n409), .A2(n413), .ZN(n396) );
  NAND2_X1 U492 ( .A1(n353), .A2(n365), .ZN(n642) );
  NOR2_X1 U493 ( .A1(n404), .A2(n660), .ZN(n365) );
  OR2_X1 U494 ( .A1(n549), .A2(n548), .ZN(n651) );
  XNOR2_X1 U495 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U496 ( .A1(G953), .A2(n695), .ZN(n696) );
  XNOR2_X1 U497 ( .A(n427), .B(n426), .ZN(n695) );
  INV_X1 U498 ( .A(KEYINPUT123), .ZN(n426) );
  AND2_X1 U499 ( .A1(n554), .A2(n399), .ZN(n353) );
  XOR2_X1 U500 ( .A(n521), .B(n520), .Z(n354) );
  INV_X1 U501 ( .A(n660), .ZN(n593) );
  AND2_X1 U502 ( .A1(n361), .A2(KEYINPUT47), .ZN(n355) );
  AND2_X1 U503 ( .A1(n411), .A2(n408), .ZN(n356) );
  XOR2_X1 U504 ( .A(G140), .B(G104), .Z(n357) );
  INV_X1 U505 ( .A(G469), .ZN(n439) );
  NAND2_X1 U506 ( .A1(G224), .A2(n735), .ZN(n358) );
  AND2_X1 U507 ( .A1(n415), .A2(n655), .ZN(n359) );
  XOR2_X1 U508 ( .A(KEYINPUT34), .B(KEYINPUT79), .Z(n360) );
  NAND2_X1 U509 ( .A1(n716), .A2(G478), .ZN(n623) );
  INV_X1 U510 ( .A(n596), .ZN(n599) );
  NAND2_X1 U511 ( .A1(n579), .A2(n578), .ZN(n596) );
  NAND2_X1 U512 ( .A1(n603), .A2(KEYINPUT72), .ZN(n361) );
  NAND2_X1 U513 ( .A1(n470), .A2(G902), .ZN(n363) );
  XNOR2_X1 U514 ( .A(n384), .B(n383), .ZN(n382) );
  XNOR2_X1 U515 ( .A(n401), .B(n360), .ZN(n438) );
  XNOR2_X2 U516 ( .A(n364), .B(n405), .ZN(n557) );
  XNOR2_X2 U517 ( .A(n366), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U518 ( .A1(n554), .A2(n390), .ZN(n366) );
  NAND2_X1 U519 ( .A1(n703), .A2(G469), .ZN(n374) );
  NAND2_X1 U520 ( .A1(n652), .A2(n636), .ZN(n550) );
  NAND2_X1 U521 ( .A1(n669), .A2(n546), .ZN(n375) );
  XNOR2_X1 U522 ( .A(n377), .B(n376), .ZN(n737) );
  INV_X1 U523 ( .A(n732), .ZN(n376) );
  XNOR2_X2 U524 ( .A(n379), .B(n378), .ZN(n612) );
  NAND2_X1 U525 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U526 ( .A(n381), .B(KEYINPUT46), .ZN(n380) );
  AND2_X1 U527 ( .A1(n419), .A2(n420), .ZN(n384) );
  NAND2_X1 U528 ( .A1(n708), .A2(n389), .ZN(n712) );
  INV_X1 U529 ( .A(n399), .ZN(n391) );
  XNOR2_X1 U530 ( .A(n510), .B(n511), .ZN(n715) );
  XNOR2_X1 U531 ( .A(n618), .B(KEYINPUT45), .ZN(n722) );
  NAND2_X1 U532 ( .A1(n561), .A2(n562), .ZN(n618) );
  NAND2_X1 U533 ( .A1(n392), .A2(n403), .ZN(n617) );
  XNOR2_X1 U534 ( .A(n393), .B(KEYINPUT30), .ZN(n570) );
  XNOR2_X1 U535 ( .A(n618), .B(n563), .ZN(n613) );
  NAND2_X1 U536 ( .A1(n411), .A2(n396), .ZN(n582) );
  XNOR2_X1 U537 ( .A(n397), .B(n632), .ZN(G57) );
  NOR2_X2 U538 ( .A1(n631), .A2(n719), .ZN(n397) );
  XNOR2_X1 U539 ( .A(n398), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U540 ( .A1(n701), .A2(n719), .ZN(n398) );
  NAND2_X1 U541 ( .A1(n499), .A2(G217), .ZN(n500) );
  XNOR2_X1 U542 ( .A(n493), .B(n494), .ZN(n499) );
  XOR2_X2 U543 ( .A(G902), .B(KEYINPUT15), .Z(n614) );
  NOR2_X2 U544 ( .A1(G902), .A2(n627), .ZN(n528) );
  NAND2_X1 U545 ( .A1(n745), .A2(KEYINPUT83), .ZN(n400) );
  NOR2_X1 U546 ( .A1(n687), .A2(n540), .ZN(n401) );
  NOR2_X1 U547 ( .A1(n544), .A2(n589), .ZN(n541) );
  XNOR2_X1 U548 ( .A(n515), .B(n514), .ZN(n517) );
  NOR2_X1 U549 ( .A1(n742), .A2(n402), .ZN(n419) );
  XNOR2_X1 U550 ( .A(n461), .B(n463), .ZN(n433) );
  XNOR2_X1 U551 ( .A(n433), .B(n432), .ZN(n431) );
  XNOR2_X2 U552 ( .A(n460), .B(G134), .ZN(n519) );
  XNOR2_X1 U553 ( .A(n691), .B(KEYINPUT74), .ZN(n403) );
  BUF_X2 U554 ( .A(n667), .Z(n404) );
  NAND2_X1 U555 ( .A1(n557), .A2(n745), .ZN(n558) );
  NAND2_X1 U556 ( .A1(n569), .A2(n414), .ZN(n413) );
  INV_X1 U557 ( .A(n413), .ZN(n407) );
  INV_X1 U558 ( .A(n673), .ZN(n408) );
  NAND2_X1 U559 ( .A1(n612), .A2(n655), .ZN(n621) );
  AND2_X2 U560 ( .A1(n612), .A2(n359), .ZN(n691) );
  INV_X1 U561 ( .A(n654), .ZN(n415) );
  NOR2_X1 U562 ( .A1(n602), .A2(n418), .ZN(n420) );
  INV_X1 U563 ( .A(n667), .ZN(n577) );
  XNOR2_X1 U564 ( .A(n423), .B(KEYINPUT28), .ZN(n579) );
  NAND2_X1 U565 ( .A1(n667), .A2(n425), .ZN(n424) );
  NAND2_X1 U566 ( .A1(n428), .A2(n694), .ZN(n427) );
  NAND2_X1 U567 ( .A1(n722), .A2(n622), .ZN(n707) );
  NAND2_X1 U568 ( .A1(n693), .A2(n692), .ZN(n429) );
  XNOR2_X2 U569 ( .A(n497), .B(n430), .ZN(n554) );
  XNOR2_X2 U570 ( .A(n436), .B(G143), .ZN(n460) );
  XNOR2_X2 U571 ( .A(G128), .B(KEYINPUT64), .ZN(n436) );
  XNOR2_X1 U572 ( .A(n700), .B(n444), .ZN(n701) );
  BUF_X1 U573 ( .A(n691), .Z(n733) );
  XNOR2_X1 U574 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U575 ( .A(n703), .B(n702), .ZN(n704) );
  AND2_X1 U576 ( .A1(G210), .A2(n466), .ZN(n442) );
  XOR2_X1 U577 ( .A(n629), .B(n628), .Z(n443) );
  XOR2_X1 U578 ( .A(n699), .B(n698), .Z(n444) );
  INV_X1 U579 ( .A(KEYINPUT66), .ZN(n514) );
  INV_X1 U580 ( .A(KEYINPUT45), .ZN(n563) );
  XNOR2_X1 U581 ( .A(n462), .B(n516), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n482), .B(n456), .ZN(n457) );
  INV_X1 U584 ( .A(KEYINPUT59), .ZN(n709) );
  INV_X1 U585 ( .A(n597), .ZN(n598) );
  XNOR2_X1 U586 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U587 ( .A(n630), .B(n443), .ZN(n631) );
  XNOR2_X1 U588 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U589 ( .A(n446), .B(n445), .ZN(n451) );
  NAND2_X1 U590 ( .A1(n735), .A2(G234), .ZN(n448) );
  XNOR2_X1 U591 ( .A(KEYINPUT65), .B(KEYINPUT8), .ZN(n447) );
  XNOR2_X1 U592 ( .A(n448), .B(n447), .ZN(n507) );
  NAND2_X1 U593 ( .A1(G217), .A2(n507), .ZN(n449) );
  XOR2_X1 U594 ( .A(n519), .B(n452), .Z(n624) );
  XOR2_X1 U595 ( .A(G101), .B(KEYINPUT3), .Z(n454) );
  XNOR2_X1 U596 ( .A(G116), .B(G113), .ZN(n453) );
  XNOR2_X1 U597 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U598 ( .A(n459), .B(n458), .ZN(n464) );
  XNOR2_X1 U599 ( .A(n460), .B(KEYINPUT86), .ZN(n461) );
  XNOR2_X2 U600 ( .A(n465), .B(n442), .ZN(n610) );
  NAND2_X1 U601 ( .A1(G214), .A2(n466), .ZN(n467) );
  XNOR2_X1 U602 ( .A(KEYINPUT87), .B(n467), .ZN(n672) );
  NOR2_X1 U603 ( .A1(n610), .A2(n672), .ZN(n468) );
  XNOR2_X1 U604 ( .A(n468), .B(KEYINPUT19), .ZN(n597) );
  XNOR2_X1 U605 ( .A(n469), .B(KEYINPUT14), .ZN(n470) );
  NAND2_X1 U606 ( .A1(G952), .A2(n470), .ZN(n686) );
  NOR2_X1 U607 ( .A1(G953), .A2(n686), .ZN(n567) );
  NAND2_X1 U608 ( .A1(G953), .A2(n471), .ZN(n564) );
  NOR2_X1 U609 ( .A1(G898), .A2(n564), .ZN(n472) );
  NOR2_X1 U610 ( .A1(n567), .A2(n472), .ZN(n473) );
  NOR2_X2 U611 ( .A1(n597), .A2(n473), .ZN(n474) );
  XNOR2_X2 U612 ( .A(n474), .B(KEYINPUT0), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n475), .B(G125), .ZN(n732) );
  XNOR2_X1 U614 ( .A(G146), .B(n732), .ZN(n511) );
  INV_X1 U615 ( .A(n511), .ZN(n488) );
  XOR2_X1 U616 ( .A(KEYINPUT99), .B(G131), .Z(n477) );
  XNOR2_X1 U617 ( .A(n477), .B(n476), .ZN(n481) );
  XOR2_X1 U618 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n479) );
  XNOR2_X1 U619 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U620 ( .A(n481), .B(n480), .ZN(n486) );
  XOR2_X1 U621 ( .A(n482), .B(KEYINPUT97), .Z(n484) );
  NAND2_X1 U622 ( .A1(n522), .A2(G214), .ZN(n483) );
  XNOR2_X1 U623 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U624 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U625 ( .A(n488), .B(n487), .ZN(n710) );
  NOR2_X1 U626 ( .A1(G902), .A2(n710), .ZN(n490) );
  XNOR2_X1 U627 ( .A(KEYINPUT13), .B(G475), .ZN(n489) );
  XNOR2_X1 U628 ( .A(n490), .B(n489), .ZN(n548) );
  NOR2_X1 U629 ( .A1(n624), .A2(G902), .ZN(n491) );
  INV_X1 U630 ( .A(n549), .ZN(n538) );
  NOR2_X1 U631 ( .A1(n548), .A2(n538), .ZN(n674) );
  INV_X1 U632 ( .A(n614), .ZN(n492) );
  NAND2_X1 U633 ( .A1(G234), .A2(n492), .ZN(n493) );
  NAND2_X1 U634 ( .A1(n499), .A2(G221), .ZN(n495) );
  XOR2_X1 U635 ( .A(KEYINPUT21), .B(n495), .Z(n576) );
  INV_X1 U636 ( .A(n576), .ZN(n657) );
  NAND2_X1 U637 ( .A1(n546), .A2(n496), .ZN(n497) );
  XOR2_X1 U638 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n501) );
  XNOR2_X1 U639 ( .A(n501), .B(n500), .ZN(n512) );
  XNOR2_X1 U640 ( .A(KEYINPUT68), .B(KEYINPUT89), .ZN(n502) );
  XNOR2_X1 U641 ( .A(G128), .B(G137), .ZN(n505) );
  XOR2_X1 U642 ( .A(G110), .B(G119), .Z(n504) );
  XNOR2_X1 U643 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U644 ( .A(n352), .B(n506), .ZN(n509) );
  NAND2_X1 U645 ( .A1(G221), .A2(n507), .ZN(n508) );
  XNOR2_X1 U646 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U647 ( .A(G137), .B(G131), .ZN(n515) );
  NAND2_X1 U648 ( .A1(G210), .A2(n522), .ZN(n523) );
  XNOR2_X1 U649 ( .A(KEYINPUT69), .B(G472), .ZN(n527) );
  XNOR2_X2 U650 ( .A(n528), .B(n527), .ZN(n667) );
  XNOR2_X2 U651 ( .A(n404), .B(n530), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT80), .B(n589), .ZN(n535) );
  NAND2_X1 U653 ( .A1(G227), .A2(n735), .ZN(n532) );
  NAND2_X1 U654 ( .A1(n535), .A2(n660), .ZN(n536) );
  NAND2_X1 U655 ( .A1(KEYINPUT44), .A2(n557), .ZN(n537) );
  NAND2_X1 U656 ( .A1(n548), .A2(n538), .ZN(n539) );
  XNOR2_X1 U657 ( .A(KEYINPUT104), .B(n539), .ZN(n581) );
  INV_X1 U658 ( .A(n546), .ZN(n540) );
  XNOR2_X1 U659 ( .A(n541), .B(KEYINPUT33), .ZN(n687) );
  NOR2_X1 U660 ( .A1(n404), .A2(n568), .ZN(n543) );
  NAND2_X1 U661 ( .A1(n543), .A2(n546), .ZN(n636) );
  XOR2_X1 U662 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n547) );
  OR2_X1 U663 ( .A1(n544), .A2(n577), .ZN(n545) );
  NAND2_X1 U664 ( .A1(n649), .A2(n651), .ZN(n676) );
  NAND2_X1 U665 ( .A1(n550), .A2(n676), .ZN(n551) );
  NAND2_X1 U666 ( .A1(n593), .A2(n589), .ZN(n552) );
  NOR2_X1 U667 ( .A1(n399), .A2(n552), .ZN(n553) );
  NAND2_X1 U668 ( .A1(n554), .A2(n553), .ZN(n633) );
  XNOR2_X1 U669 ( .A(n558), .B(KEYINPUT44), .ZN(n560) );
  INV_X1 U670 ( .A(KEYINPUT83), .ZN(n559) );
  NAND2_X1 U671 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U672 ( .A(KEYINPUT105), .B(n564), .Z(n565) );
  NOR2_X1 U673 ( .A1(G900), .A2(n565), .ZN(n566) );
  INV_X1 U674 ( .A(n610), .ZN(n590) );
  NOR2_X1 U675 ( .A1(n651), .A2(n571), .ZN(n654) );
  INV_X1 U676 ( .A(n674), .ZN(n573) );
  NOR2_X1 U677 ( .A1(n673), .A2(n672), .ZN(n572) );
  XNOR2_X1 U678 ( .A(n572), .B(KEYINPUT109), .ZN(n677) );
  XNOR2_X1 U679 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n574) );
  XNOR2_X1 U680 ( .A(n575), .B(n574), .ZN(n688) );
  NOR2_X1 U681 ( .A1(n688), .A2(n596), .ZN(n580) );
  OR2_X1 U682 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U683 ( .A1(n672), .A2(n584), .ZN(n587) );
  NOR2_X1 U684 ( .A1(n649), .A2(n585), .ZN(n586) );
  NAND2_X1 U685 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U686 ( .A1(n606), .A2(n590), .ZN(n592) );
  XNOR2_X1 U687 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n591) );
  NOR2_X1 U688 ( .A1(KEYINPUT72), .A2(n604), .ZN(n600) );
  NOR2_X1 U689 ( .A1(KEYINPUT47), .A2(n600), .ZN(n601) );
  NOR2_X1 U690 ( .A1(n676), .A2(n601), .ZN(n602) );
  INV_X1 U691 ( .A(n604), .ZN(n603) );
  NOR2_X1 U692 ( .A1(n649), .A2(n604), .ZN(n647) );
  NOR2_X1 U693 ( .A1(n651), .A2(n604), .ZN(n643) );
  NOR2_X1 U694 ( .A1(n647), .A2(n643), .ZN(n605) );
  XOR2_X1 U695 ( .A(n606), .B(KEYINPUT106), .Z(n607) );
  NOR2_X1 U696 ( .A1(n660), .A2(n607), .ZN(n608) );
  XNOR2_X1 U697 ( .A(KEYINPUT43), .B(n608), .ZN(n609) );
  XNOR2_X1 U698 ( .A(n609), .B(KEYINPUT107), .ZN(n611) );
  NAND2_X1 U699 ( .A1(n611), .A2(n394), .ZN(n655) );
  XNOR2_X1 U700 ( .A(n614), .B(KEYINPUT82), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n615), .A2(KEYINPUT2), .ZN(n616) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n692) );
  OR2_X1 U703 ( .A1(n692), .A2(n654), .ZN(n619) );
  XOR2_X1 U704 ( .A(KEYINPUT81), .B(n619), .Z(n620) );
  NOR2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U706 ( .A(n623), .B(n624), .ZN(n625) );
  NOR2_X2 U707 ( .A1(n625), .A2(n719), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT124), .ZN(G63) );
  INV_X1 U709 ( .A(KEYINPUT63), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n716), .A2(G472), .ZN(n630) );
  XNOR2_X1 U711 ( .A(KEYINPUT62), .B(KEYINPUT114), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n627), .B(KEYINPUT113), .ZN(n628) );
  XNOR2_X1 U713 ( .A(G101), .B(n633), .ZN(G3) );
  NOR2_X1 U714 ( .A1(n649), .A2(n636), .ZN(n635) );
  XNOR2_X1 U715 ( .A(G104), .B(KEYINPUT115), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n635), .B(n634), .ZN(G6) );
  NOR2_X1 U717 ( .A1(n651), .A2(n636), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n638) );
  XNOR2_X1 U719 ( .A(G107), .B(KEYINPUT26), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U721 ( .A(KEYINPUT116), .B(n639), .ZN(n640) );
  XNOR2_X1 U722 ( .A(n641), .B(n640), .ZN(G9) );
  XNOR2_X1 U723 ( .A(G110), .B(n642), .ZN(G12) );
  XNOR2_X1 U724 ( .A(G128), .B(n643), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n644), .B(KEYINPUT29), .ZN(G30) );
  XOR2_X1 U726 ( .A(n645), .B(G143), .Z(n646) );
  XNOR2_X1 U727 ( .A(KEYINPUT118), .B(n646), .ZN(G45) );
  XNOR2_X1 U728 ( .A(G146), .B(n647), .ZN(n648) );
  XNOR2_X1 U729 ( .A(n648), .B(KEYINPUT119), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n652), .A2(n649), .ZN(n650) );
  XOR2_X1 U731 ( .A(G113), .B(n650), .Z(G15) );
  NOR2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U733 ( .A(G116), .B(n653), .Z(G18) );
  XOR2_X1 U734 ( .A(G134), .B(n654), .Z(G36) );
  XNOR2_X1 U735 ( .A(G140), .B(n655), .ZN(G42) );
  NAND2_X1 U736 ( .A1(n657), .A2(n399), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n658), .B(KEYINPUT121), .ZN(n659) );
  XNOR2_X1 U738 ( .A(KEYINPUT49), .B(n659), .ZN(n665) );
  OR2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(KEYINPUT122), .ZN(n663) );
  XNOR2_X1 U741 ( .A(KEYINPUT50), .B(n663), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U743 ( .A1(n404), .A2(n666), .ZN(n668) );
  NOR2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U745 ( .A(KEYINPUT51), .B(n670), .Z(n671) );
  NOR2_X1 U746 ( .A1(n688), .A2(n671), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n673), .A2(n672), .ZN(n675) );
  AND2_X1 U748 ( .A1(n675), .A2(n674), .ZN(n680) );
  INV_X1 U749 ( .A(n676), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U752 ( .A1(n681), .A2(n687), .ZN(n682) );
  NOR2_X1 U753 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U754 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  NOR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U758 ( .A1(n733), .A2(n722), .ZN(n693) );
  XNOR2_X1 U759 ( .A(KEYINPUT53), .B(n696), .ZN(G75) );
  NAND2_X1 U760 ( .A1(n716), .A2(G210), .ZN(n700) );
  XOR2_X1 U761 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n699) );
  XNOR2_X1 U762 ( .A(n697), .B(KEYINPUT85), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n716), .A2(G469), .ZN(n705) );
  XOR2_X1 U764 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  NOR2_X1 U765 ( .A1(n719), .A2(n706), .ZN(G54) );
  AND2_X1 U766 ( .A1(G475), .A2(n707), .ZN(n708) );
  NOR2_X1 U767 ( .A1(n719), .A2(n713), .ZN(n714) );
  XNOR2_X1 U768 ( .A(KEYINPUT60), .B(n714), .ZN(G60) );
  NAND2_X1 U769 ( .A1(n716), .A2(G217), .ZN(n717) );
  XNOR2_X1 U770 ( .A(n717), .B(n718), .ZN(n720) );
  NOR2_X2 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n721), .B(KEYINPUT126), .ZN(G66) );
  NAND2_X1 U773 ( .A1(n735), .A2(n722), .ZN(n726) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n723) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n731) );
  XOR2_X1 U778 ( .A(KEYINPUT127), .B(n727), .Z(n729) );
  NOR2_X1 U779 ( .A1(G898), .A2(n735), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(G69) );
  INV_X1 U782 ( .A(n737), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n734), .B(n733), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n741) );
  XNOR2_X1 U785 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U789 ( .A(KEYINPUT120), .B(KEYINPUT37), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U791 ( .A(G125), .B(n744), .ZN(G27) );
  XNOR2_X1 U792 ( .A(n745), .B(G122), .ZN(G24) );
  XNOR2_X1 U793 ( .A(n746), .B(G119), .ZN(G21) );
  XOR2_X1 U794 ( .A(n747), .B(G131), .Z(G33) );
  XOR2_X1 U795 ( .A(G137), .B(n748), .Z(G39) );
endmodule

