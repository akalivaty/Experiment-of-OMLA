//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G50), .A2(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n212), .B(new_n214), .C1(G77), .C2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n208), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT64), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n231), .A2(G1), .A3(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n206), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g0036(.A(G50), .B1(G58), .B2(G68), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n225), .B(new_n228), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G226), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n244), .B(KEYINPUT68), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G264), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n219), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n252), .B(KEYINPUT69), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT70), .ZN(new_n254));
  XOR2_X1   g0054(.A(G107), .B(G116), .Z(new_n255));
  XNOR2_X1  g0055(.A(G87), .B(G97), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(KEYINPUT10), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(KEYINPUT75), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n233), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G222), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G223), .A2(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n264), .B(new_n272), .C1(G77), .C2(new_n268), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT71), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G41), .A2(G45), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(G1), .ZN(new_n279));
  INV_X1    g0079(.A(new_n278), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(KEYINPUT71), .A3(new_n205), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n276), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n205), .A2(KEYINPUT72), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n274), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G226), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n273), .A2(new_n282), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI211_X1 g0091(.A(new_n260), .B(new_n291), .C1(G200), .C2(new_n289), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n230), .A2(new_n232), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n206), .A2(G33), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT73), .ZN(new_n297));
  XOR2_X1   g0097(.A(KEYINPUT8), .B(G58), .Z(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G58), .A2(G68), .ZN(new_n300));
  INV_X1    g0100(.A(G50), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n206), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(G150), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n295), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n294), .B1(G20), .B2(new_n286), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(G50), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n286), .A2(G13), .A3(G20), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n301), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT9), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n292), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT75), .A3(new_n259), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n259), .A2(KEYINPUT75), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n292), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n289), .A2(G179), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT74), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n289), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(KEYINPUT74), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n318), .A2(new_n311), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n298), .ZN(new_n323));
  INV_X1    g0123(.A(new_n303), .ZN(new_n324));
  INV_X1    g0124(.A(G77), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n323), .A2(new_n324), .B1(new_n206), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n296), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n294), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n306), .A2(G77), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(G77), .C2(new_n308), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n269), .A2(G232), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n268), .B(new_n333), .C1(new_n211), .C2(new_n269), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n264), .B(new_n334), .C1(G107), .C2(new_n268), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n287), .A2(G244), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n282), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n338), .B2(G190), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n338), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n314), .A2(new_n316), .A3(new_n322), .A4(new_n341), .ZN(new_n342));
  OR3_X1    g0142(.A1(new_n308), .A2(KEYINPUT12), .A3(G68), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT12), .B1(new_n308), .B2(G68), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(new_n306), .B2(G68), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n297), .A2(G77), .B1(G20), .B2(new_n210), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n301), .B2(new_n324), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT11), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n347), .A2(new_n348), .A3(new_n294), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(new_n347), .B2(new_n294), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n287), .A2(G238), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n282), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n269), .A2(G232), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n268), .B(new_n355), .C1(G226), .C2(G1698), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n263), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT13), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n354), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n264), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n352), .A4(new_n282), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n290), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n340), .B1(new_n358), .B2(new_n362), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n351), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(G169), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n358), .A2(new_n362), .A3(G179), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n370), .A3(G169), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n366), .B1(new_n372), .B2(new_n351), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n265), .ZN(new_n375));
  NAND2_X1  g0175(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(G33), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G226), .A2(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n269), .A2(G223), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n377), .A2(new_n266), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT77), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  NOR2_X1   g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  AND2_X1   g0185(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n388), .B2(G33), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n379), .A2(new_n378), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n384), .B(new_n381), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n383), .A2(new_n391), .A3(new_n264), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n287), .A2(G232), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n393), .A2(new_n282), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(G179), .A3(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n392), .A2(new_n394), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n319), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n389), .A2(new_n398), .A3(new_n206), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n377), .A2(new_n206), .A3(new_n266), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT7), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(G68), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G58), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n210), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n404), .B2(new_n300), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n303), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  AOI21_X1  g0210(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT7), .B(new_n411), .C1(new_n388), .C2(G33), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n266), .A2(new_n206), .A3(new_n267), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n398), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n210), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n410), .B1(new_n415), .B2(new_n407), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n409), .A2(new_n294), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n308), .A2(new_n323), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n306), .B2(new_n323), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n397), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n397), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n392), .A2(G190), .A3(new_n394), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n417), .A2(new_n427), .A3(new_n419), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n392), .A2(new_n394), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G200), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n426), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n419), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n375), .A2(new_n376), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n398), .B1(new_n434), .B2(new_n261), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n411), .B1(new_n398), .B2(new_n413), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n408), .B1(new_n436), .B2(new_n210), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n295), .B1(new_n437), .B2(new_n410), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n433), .B1(new_n438), .B2(new_n409), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(KEYINPUT17), .A3(new_n430), .A4(new_n427), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n337), .A2(new_n319), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(new_n332), .C1(G179), .C2(new_n337), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n373), .A2(new_n425), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n342), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT78), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n342), .B2(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n268), .A2(new_n206), .A3(G87), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT22), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n206), .A2(G107), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT23), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n261), .A2(new_n218), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n377), .B2(new_n266), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(G87), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n452), .B(new_n454), .C1(new_n457), .C2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT24), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n451), .B(new_n216), .C1(new_n377), .C2(new_n266), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n206), .B1(new_n461), .B2(new_n455), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(KEYINPUT24), .A3(new_n452), .A4(new_n454), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n294), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  OR2_X1    g0265(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n466));
  NAND2_X1  g0266(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n309), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT85), .B(KEYINPUT25), .C1(new_n308), .C2(G107), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n286), .A2(G33), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n294), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n286), .A2(KEYINPUT79), .A3(G33), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n308), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G107), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n464), .A2(new_n468), .A3(new_n469), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n377), .A2(new_n266), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(G257), .A3(G1698), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G294), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n482), .A2(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(KEYINPUT87), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n483), .A2(G33), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(G1698), .B1(new_n377), .B2(new_n266), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(G250), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n478), .A2(KEYINPUT86), .A3(G257), .A4(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n481), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n264), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT5), .B(G41), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n286), .A2(new_n491), .A3(G45), .ZN(new_n492));
  INV_X1    g0292(.A(new_n274), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G264), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT88), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n276), .A2(G45), .A3(new_n286), .A4(new_n491), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT88), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n490), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n340), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n490), .A2(new_n290), .A3(new_n500), .A4(new_n497), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n477), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n477), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n492), .A2(new_n275), .A3(new_n274), .ZN(new_n508));
  OAI21_X1  g0308(.A(G169), .B1(new_n498), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n499), .A2(G179), .A3(new_n500), .A4(new_n502), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n500), .B1(new_n494), .B2(new_n219), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT82), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n377), .A2(new_n266), .B1(new_n495), .B2(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n222), .A2(new_n269), .ZN(new_n517));
  INV_X1    g0317(.A(new_n268), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n516), .A2(new_n517), .B1(G303), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n515), .B1(new_n519), .B2(new_n263), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n495), .A2(G1698), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n386), .A2(new_n387), .A3(new_n261), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n517), .B(new_n521), .C1(new_n522), .C2(new_n385), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(G303), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(KEYINPUT82), .A3(new_n264), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n514), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n472), .A2(G116), .A3(new_n308), .A4(new_n473), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(new_n206), .C1(G33), .C2(new_n221), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n218), .A2(G20), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n294), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n294), .A2(KEYINPUT20), .A3(new_n530), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n308), .A2(G116), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n528), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G169), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n513), .B1(new_n527), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT84), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n514), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT82), .B1(new_n525), .B2(new_n264), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n515), .B(new_n263), .C1(new_n523), .C2(new_n524), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n537), .B1(new_n534), .B2(new_n535), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n319), .B1(new_n548), .B2(new_n528), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(KEYINPUT84), .A3(new_n513), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(G200), .ZN(new_n553));
  INV_X1    g0353(.A(new_n539), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n554), .C1(new_n290), .C2(new_n547), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT83), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n547), .A2(KEYINPUT21), .A3(new_n549), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n520), .A2(new_n526), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n558), .A2(G179), .A3(new_n539), .A4(new_n544), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n556), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n557), .A2(new_n556), .A3(new_n559), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n552), .B(new_n555), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT80), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n286), .A2(G45), .A3(new_n275), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n493), .ZN(new_n565));
  AOI21_X1  g0365(.A(G250), .B1(new_n286), .B2(G45), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n283), .A2(new_n285), .ZN(new_n568));
  INV_X1    g0368(.A(G45), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n217), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n570), .A2(KEYINPUT80), .A3(new_n493), .A4(new_n564), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G238), .A2(G1698), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n269), .A2(G244), .ZN(new_n574));
  AOI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n377), .C2(new_n266), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n264), .B1(new_n575), .B2(new_n455), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT81), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n572), .A2(new_n576), .A3(KEYINPUT81), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n319), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G179), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n572), .A2(KEYINPUT81), .A3(new_n576), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(new_n577), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n478), .A2(new_n206), .A3(G68), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n206), .B1(new_n354), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G87), .B2(new_n203), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n354), .B2(G20), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(new_n294), .B1(new_n309), .B2(new_n328), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n328), .B2(new_n474), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n580), .A2(new_n583), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n578), .A2(G200), .A3(new_n579), .ZN(new_n593));
  OAI21_X1  g0393(.A(G190), .B1(new_n582), .B2(new_n577), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n475), .A2(G87), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n595), .A2(new_n590), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n475), .A2(G97), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n309), .A2(new_n221), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n324), .A2(new_n325), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n221), .A2(new_n465), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n202), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n206), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n412), .A2(new_n414), .ZN(new_n606));
  AOI211_X1 g0406(.A(new_n600), .B(new_n605), .C1(new_n606), .C2(G107), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n598), .B(new_n599), .C1(new_n607), .C2(new_n295), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT4), .B1(new_n486), .B2(G244), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n269), .ZN(new_n611));
  INV_X1    g0411(.A(G244), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n529), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n264), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n494), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G257), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n500), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n319), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n614), .A2(new_n581), .A3(new_n500), .A4(new_n616), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n608), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n607), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(new_n294), .B1(G97), .B2(new_n475), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(G200), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n614), .A2(G190), .A3(new_n500), .A4(new_n616), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n599), .A4(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n592), .A2(new_n597), .A3(new_n620), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n562), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n449), .A2(new_n512), .A3(new_n627), .ZN(G372));
  AND2_X1   g0428(.A1(new_n557), .A2(new_n559), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT84), .B1(new_n550), .B2(new_n513), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n542), .B(KEYINPUT21), .C1(new_n547), .C2(new_n549), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT89), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n510), .A2(new_n509), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n477), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n552), .A2(KEYINPUT89), .A3(new_n629), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n572), .A2(new_n576), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G200), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n594), .A2(new_n596), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n625), .A3(new_n620), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n501), .B1(new_n490), .B2(new_n497), .ZN(new_n643));
  AOI211_X1 g0443(.A(KEYINPUT88), .B(new_n496), .C1(new_n489), .C2(new_n264), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n643), .A2(new_n644), .A3(new_n508), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n505), .B1(new_n645), .B2(G200), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n642), .B1(new_n507), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n638), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n639), .A2(new_n319), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n583), .A2(new_n591), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n620), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n641), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g0455(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n656));
  NAND4_X1  g0456(.A1(new_n592), .A2(new_n597), .A3(new_n652), .A4(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n449), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n372), .A2(new_n351), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n366), .A2(new_n443), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n441), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n397), .A2(new_n420), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n397), .B2(new_n420), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n423), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n319), .B1(new_n392), .B2(new_n394), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(G179), .B2(new_n396), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT91), .B1(new_n671), .B2(new_n439), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(KEYINPUT18), .A3(new_n666), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n314), .A2(new_n316), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n322), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n660), .A2(new_n679), .ZN(G369));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n634), .A2(new_n637), .ZN(new_n682));
  INV_X1    g0482(.A(G13), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G20), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n286), .A2(new_n684), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n685), .A2(KEYINPUT92), .A3(KEYINPUT27), .ZN(new_n686));
  INV_X1    g0486(.A(G213), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n685), .B2(KEYINPUT27), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT92), .B1(new_n685), .B2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n554), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n682), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n562), .A2(new_n694), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n681), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT93), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n507), .B2(new_n693), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n477), .A2(KEYINPUT93), .A3(new_n692), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n512), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n511), .A2(new_n692), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n511), .A2(new_n693), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n557), .A2(new_n559), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT83), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n557), .A2(new_n559), .A3(new_n556), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n543), .B2(new_n551), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n692), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n512), .A2(new_n710), .A3(new_n699), .A4(new_n700), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n704), .A2(new_n705), .A3(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n226), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G1), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n202), .A2(new_n216), .A3(new_n218), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(new_n237), .B2(new_n715), .ZN(new_n718));
  XOR2_X1   g0518(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n719));
  XNOR2_X1  g0519(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n659), .A2(new_n721), .A3(new_n693), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n709), .A2(new_n636), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n651), .B1(new_n723), .B2(new_n647), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n641), .A2(new_n650), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT26), .A4(new_n652), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT95), .B1(new_n653), .B2(new_n654), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n592), .A2(new_n597), .A3(new_n652), .ZN(new_n729));
  INV_X1    g0529(.A(new_n656), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n692), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n722), .B1(new_n721), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  INV_X1    g0535(.A(new_n617), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n499), .A2(new_n502), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(G179), .B(new_n527), .C1(new_n582), .C2(new_n577), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n643), .A2(new_n644), .A3(new_n617), .ZN(new_n740));
  OAI211_X1 g0540(.A(G179), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n578), .B2(new_n579), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n736), .A2(new_n527), .A3(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n503), .A2(new_n639), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n746), .B2(new_n692), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n627), .A2(new_n512), .A3(new_n693), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n681), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n734), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n720), .B1(new_n752), .B2(G1), .ZN(G364));
  OR2_X1    g0553(.A1(new_n237), .A2(G45), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n713), .A2(new_n478), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(new_n254), .C2(new_n569), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n226), .A2(G355), .A3(new_n268), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n757), .C1(G116), .C2(new_n226), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT96), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n234), .B1(G20), .B2(new_n319), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT97), .Z(new_n765));
  NAND2_X1  g0565(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n716), .B1(G45), .B2(new_n684), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n695), .A2(new_n696), .A3(new_n763), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(G20), .B1(new_n770), .B2(new_n290), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT99), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n483), .A2(new_n484), .ZN(new_n776));
  INV_X1    g0576(.A(G326), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n206), .A2(new_n581), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT100), .Z(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n268), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n778), .A2(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G200), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n770), .A2(new_n206), .A3(G190), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n784), .A2(G322), .B1(new_n785), .B2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(new_n778), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(new_n340), .A3(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI211_X1 g0590(.A(new_n782), .B(new_n786), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n581), .A2(G200), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT98), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n290), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n794), .A2(G190), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n791), .A2(new_n798), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n785), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT32), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n268), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n796), .A2(new_n216), .B1(new_n301), .B2(new_n779), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G107), .C2(new_n799), .ZN(new_n814));
  INV_X1    g0614(.A(new_n784), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n775), .A2(new_n221), .B1(new_n403), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n811), .B2(new_n810), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n814), .B(new_n817), .C1(new_n325), .C2(new_n804), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G68), .B2(new_n788), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n760), .B1(new_n807), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n697), .ZN(new_n822));
  INV_X1    g0622(.A(new_n767), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n695), .A2(new_n696), .A3(new_n681), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(new_n825), .ZN(G396));
  AOI21_X1  g0626(.A(new_n692), .B1(new_n648), .B2(new_n658), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n443), .A2(new_n692), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n332), .A2(new_n692), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n341), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n829), .B1(new_n443), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n827), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(new_n751), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n823), .ZN(new_n835));
  INV_X1    g0635(.A(new_n832), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n761), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G150), .A2(new_n788), .B1(new_n784), .B2(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n779), .C1(new_n809), .C2(new_n804), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  AOI22_X1  g0641(.A1(G50), .A2(new_n795), .B1(new_n799), .B2(G68), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT101), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n478), .B1(new_n844), .B2(new_n808), .C1(new_n775), .C2(new_n403), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n841), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G87), .A2(new_n799), .B1(new_n795), .B2(G107), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n218), .B2(new_n804), .C1(new_n801), .C2(new_n789), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n808), .A2(new_n805), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n815), .A2(new_n482), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n518), .B1(new_n797), .B2(new_n779), .C1(new_n775), .C2(new_n221), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n760), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n760), .A2(new_n761), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n325), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n837), .A2(new_n853), .A3(new_n767), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n835), .A2(new_n856), .ZN(G384));
  AND2_X1   g0657(.A1(new_n603), .A2(new_n604), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT35), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n236), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n860), .B(G116), .C1(new_n859), .C2(new_n858), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT36), .ZN(new_n862));
  OAI21_X1  g0662(.A(G77), .B1(new_n403), .B2(new_n210), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n863), .A2(new_n237), .B1(G50), .B2(new_n210), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n683), .A3(new_n568), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n422), .A2(new_n432), .A3(new_n440), .A4(new_n424), .ZN(new_n866));
  INV_X1    g0666(.A(new_n690), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n409), .A2(new_n294), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT16), .B1(new_n402), .B2(new_n408), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n419), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n439), .A2(new_n430), .A3(new_n427), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n420), .A2(new_n867), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n872), .A2(new_n421), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n428), .A2(new_n431), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n671), .A2(new_n690), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n875), .B1(new_n878), .B2(new_n874), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n871), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n661), .A2(new_n692), .ZN(new_n888));
  INV_X1    g0688(.A(new_n883), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n876), .B1(new_n672), .B2(new_n666), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n873), .B1(new_n890), .B2(KEYINPUT102), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT102), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n892), .B(new_n876), .C1(new_n672), .C2(new_n666), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n875), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n873), .B1(new_n674), .B2(new_n441), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n889), .B1(new_n898), .B2(new_n881), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n887), .B(new_n888), .C1(new_n899), .C2(KEYINPUT39), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n674), .A2(new_n867), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n661), .A2(new_n693), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n351), .A2(new_n692), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n373), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n659), .A2(new_n693), .A3(new_n832), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(new_n828), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n901), .B1(new_n909), .B2(new_n884), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n678), .B1(new_n734), .B2(new_n449), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n911), .B(new_n912), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n906), .A2(new_n832), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n749), .B2(new_n750), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n895), .B2(new_n897), .ZN(new_n916));
  OAI211_X1 g0716(.A(KEYINPUT40), .B(new_n915), .C1(new_n916), .C2(new_n889), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n746), .A2(new_n692), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT31), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n750), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n914), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n884), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n917), .A2(G330), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n449), .A2(G330), .A3(new_n922), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n917), .A2(new_n449), .A3(new_n926), .A4(new_n922), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n913), .A2(new_n931), .B1(new_n286), .B2(new_n684), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT103), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n913), .A2(new_n931), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n862), .B(new_n865), .C1(new_n933), .C2(new_n934), .ZN(G367));
  OAI22_X1  g0735(.A1(new_n403), .A2(new_n796), .B1(new_n800), .B2(new_n325), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G150), .B2(new_n784), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n785), .A2(G137), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n775), .A2(new_n210), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT109), .ZN(new_n940));
  AOI22_X1  g0740(.A1(G50), .A2(new_n803), .B1(new_n788), .B2(G159), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n518), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n937), .A2(new_n938), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(G143), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n943), .B1(new_n940), .B2(new_n941), .C1(new_n944), .C2(new_n779), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n775), .A2(new_n465), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n795), .A2(G116), .ZN(new_n947));
  OR2_X1    g0747(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n948));
  NAND2_X1  g0748(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n789), .A2(new_n776), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n804), .A2(new_n801), .ZN(new_n952));
  NOR4_X1   g0752(.A1(new_n950), .A2(new_n478), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n785), .A2(G317), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n800), .A2(new_n221), .B1(new_n805), .B2(new_n779), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n947), .B2(new_n949), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n784), .A2(G303), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n953), .A2(new_n954), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n945), .B1(new_n946), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT47), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n760), .ZN(new_n961));
  INV_X1    g0761(.A(new_n755), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n764), .B1(new_n226), .B2(new_n328), .C1(new_n248), .C2(new_n962), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n961), .A2(new_n767), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n596), .A2(new_n693), .ZN(new_n965));
  MUX2_X1   g0765(.A(new_n725), .B(new_n651), .S(new_n965), .Z(new_n966));
  OR3_X1    g0766(.A1(new_n966), .A2(G20), .A3(new_n762), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n205), .B1(new_n684), .B2(G45), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n711), .A2(new_n705), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n608), .A2(new_n692), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n625), .A2(new_n620), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n652), .A2(new_n692), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT45), .B1(new_n971), .B2(new_n976), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n711), .A2(new_n982), .A3(new_n705), .A4(new_n975), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n971), .A2(new_n976), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n697), .B(new_n703), .C1(new_n984), .C2(new_n988), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n981), .A2(new_n983), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n990), .A2(new_n704), .A3(new_n980), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT106), .B1(new_n703), .B2(new_n710), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT106), .ZN(new_n994));
  INV_X1    g0794(.A(new_n710), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n701), .A2(new_n994), .A3(new_n702), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n711), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n697), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n993), .A2(new_n822), .A3(new_n711), .A4(new_n996), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n752), .ZN(new_n1001));
  OAI21_X1  g0801(.A(KEYINPUT107), .B1(new_n992), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n752), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n998), .B2(new_n999), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT107), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1004), .A2(new_n989), .A3(new_n991), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n752), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n714), .B(KEYINPUT41), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n970), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n711), .A2(new_n976), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT42), .Z(new_n1012));
  OR2_X1    g0812(.A1(new_n636), .A2(new_n973), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n692), .B1(new_n1013), .B2(new_n620), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n966), .B(KEYINPUT43), .Z(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT104), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT104), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n1016), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n704), .A2(new_n976), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n968), .B1(new_n1010), .B2(new_n1026), .ZN(G387));
  NAND3_X1  g0827(.A1(new_n1003), .A2(new_n999), .A3(new_n998), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1001), .A2(new_n1028), .A3(new_n714), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1000), .A2(new_n970), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n389), .B1(new_n808), .B2(new_n777), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G311), .A2(new_n788), .B1(new_n784), .B2(G317), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n779), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(G322), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(new_n797), .C2(new_n804), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT48), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n801), .B2(new_n775), .C1(new_n776), .C2(new_n796), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT49), .Z(new_n1038));
  AOI211_X1 g0838(.A(new_n1031), .B(new_n1038), .C1(G116), .C2(new_n799), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n804), .A2(new_n210), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n775), .A2(new_n328), .B1(new_n323), .B2(new_n789), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n799), .A2(G97), .B1(G150), .B2(new_n785), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1042), .B(new_n478), .C1(new_n325), .C2(new_n796), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT110), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .C1(new_n809), .C2(new_n779), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1040), .B(new_n1046), .C1(G50), .C2(new_n784), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n760), .B1(new_n1039), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n298), .A2(new_n301), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n210), .A2(new_n325), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1050), .A2(G45), .A3(new_n1051), .A4(new_n717), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n755), .B1(new_n244), .B2(new_n569), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n226), .A2(new_n268), .A3(new_n717), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n226), .A2(G107), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n765), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n701), .A2(new_n702), .A3(new_n763), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1048), .A2(new_n767), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1029), .A2(new_n1030), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT111), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(G393));
  NAND3_X1  g0862(.A1(new_n989), .A2(new_n970), .A3(new_n991), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n764), .B1(new_n221), .B2(new_n226), .C1(new_n962), .C2(new_n257), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n823), .B1(new_n976), .B2(new_n763), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G311), .A2(new_n784), .B1(new_n1033), .B2(G317), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n268), .B1(new_n785), .B2(G322), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n218), .B2(new_n775), .C1(new_n800), .C2(new_n465), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(G283), .C2(new_n795), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n482), .B2(new_n804), .C1(new_n797), .C2(new_n789), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT114), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n775), .A2(new_n325), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G87), .B2(new_n799), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT113), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n796), .A2(new_n210), .B1(new_n944), .B2(new_n808), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1074), .B(new_n478), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n803), .A2(new_n298), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n788), .A2(G50), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G159), .A2(new_n784), .B1(new_n1033), .B2(G150), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1072), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n760), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1064), .B(new_n1065), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1063), .A2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1002), .A2(new_n1006), .B1(new_n992), .B2(new_n1001), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n714), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G390));
  AOI21_X1  g0891(.A(KEYINPUT115), .B1(new_n912), .B2(new_n928), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n723), .A2(new_n647), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n732), .A2(new_n650), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n721), .B1(new_n1094), .B2(new_n693), .ZN(new_n1095));
  AOI211_X1 g0895(.A(KEYINPUT29), .B(new_n692), .C1(new_n648), .C2(new_n658), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n449), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1097), .A2(new_n928), .A3(KEYINPUT115), .A4(new_n679), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n908), .A2(new_n828), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n906), .B1(new_n751), .B2(new_n832), .ZN(new_n1102));
  AND4_X1   g0902(.A1(G330), .A2(new_n922), .A3(new_n832), .A4(new_n906), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n922), .A2(G330), .A3(new_n832), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n907), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n751), .A2(new_n832), .A3(new_n906), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n831), .A2(new_n443), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n829), .B1(new_n733), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n888), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n896), .B1(new_n894), .B2(new_n875), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n883), .B1(new_n1113), .B2(KEYINPUT38), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(new_n1109), .C2(new_n907), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n888), .B1(new_n1101), .B2(new_n906), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n886), .B1(new_n1114), .B2(new_n885), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1103), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1115), .B(new_n1107), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1100), .A2(new_n1111), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1097), .A2(new_n679), .A3(new_n928), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT115), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1111), .A2(new_n1124), .A3(new_n1098), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n887), .B1(new_n899), .B2(KEYINPUT39), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n829), .B1(new_n827), .B2(new_n832), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1112), .B1(new_n1127), .B2(new_n907), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1107), .B1(new_n1129), .B2(new_n1115), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1120), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1121), .A2(new_n1132), .A3(new_n714), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1119), .A2(new_n970), .A3(new_n1120), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1126), .A2(new_n761), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n854), .A2(new_n323), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n795), .A2(G150), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT53), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n518), .B(new_n1138), .C1(G125), .C2(new_n785), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1033), .A2(G128), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n775), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(G159), .B1(G50), .B2(new_n799), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G137), .A2(new_n788), .B1(new_n784), .B2(G132), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT54), .B(G143), .Z(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n803), .B2(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n800), .A2(new_n210), .B1(new_n465), .B2(new_n789), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1073), .B(new_n1147), .C1(G97), .C2(new_n803), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n784), .A2(G116), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n795), .A2(G87), .B1(G283), .B2(new_n1033), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1148), .A2(new_n518), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G294), .B2(new_n785), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n760), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1135), .A2(new_n767), .A3(new_n1136), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT116), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1134), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1134), .B2(new_n1154), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1133), .B1(new_n1156), .B2(new_n1157), .ZN(G378));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n676), .A2(new_n322), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT119), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n311), .A2(new_n867), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT119), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1161), .B(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(new_n1163), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1160), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1163), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n1159), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n927), .A2(new_n910), .A3(new_n900), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n927), .B1(new_n900), .B2(new_n910), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n927), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n911), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n927), .A2(new_n910), .A3(new_n900), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1178), .A2(new_n1172), .A3(new_n1169), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1100), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n1184), .A3(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n714), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1169), .A2(new_n761), .A3(new_n1172), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1141), .A2(G150), .B1(G125), .B2(new_n1033), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT118), .Z(new_n1191));
  INV_X1    g0991(.A(G128), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n815), .C1(new_n839), .C2(new_n804), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G132), .B2(new_n788), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1145), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n796), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n1196), .B2(KEYINPUT59), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G33), .B1(new_n785), .B2(G124), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n809), .C2(new_n800), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT58), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n796), .A2(new_n325), .B1(new_n465), .B2(new_n815), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n939), .B(new_n1202), .C1(G116), .C2(new_n1033), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n800), .A2(new_n403), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n377), .A2(new_n262), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n804), .A2(new_n328), .B1(new_n801), .B2(new_n808), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1204), .A2(new_n385), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1203), .B(new_n1207), .C1(new_n221), .C2(new_n789), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1199), .A2(new_n1200), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1208), .A2(new_n1201), .B1(new_n301), .B2(new_n1205), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT117), .Z(new_n1211));
  OAI21_X1  g1011(.A(new_n760), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n854), .A2(new_n301), .ZN(new_n1213));
  AND4_X1   g1013(.A1(new_n767), .A2(new_n1189), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1181), .B2(new_n970), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1188), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(G375));
  AOI22_X1  g1017(.A1(new_n1141), .A2(new_n327), .B1(G97), .B2(new_n795), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n218), .B2(new_n789), .C1(new_n482), .C2(new_n779), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n518), .B1(new_n465), .B2(new_n804), .C1(new_n800), .C2(new_n325), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n801), .B2(new_n815), .C1(new_n797), .C2(new_n808), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1141), .A2(G50), .B1(G150), .B2(new_n803), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT122), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n478), .B1(new_n796), .B2(new_n809), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n815), .A2(new_n839), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n789), .A2(new_n1195), .B1(new_n844), .B2(new_n779), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1225), .A2(new_n1204), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1224), .B(new_n1228), .C1(new_n1192), .C2(new_n808), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1086), .B1(new_n1222), .B2(new_n1229), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n823), .B(new_n1230), .C1(new_n210), .C2(new_n854), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n907), .A2(new_n761), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT121), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1111), .A2(new_n970), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1100), .A2(new_n1111), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1009), .B(KEYINPUT120), .Z(new_n1236));
  NAND2_X1  g1036(.A1(new_n1125), .A2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1235), .B2(new_n1237), .ZN(G381));
  OAI211_X1 g1038(.A(new_n968), .B(new_n1090), .C1(new_n1010), .C2(new_n1026), .ZN(new_n1239));
  OR2_X1    g1039(.A1(G381), .A2(G384), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1239), .A2(G396), .A3(G393), .A4(new_n1240), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1134), .A2(new_n1154), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1133), .A2(KEYINPUT123), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT123), .B1(new_n1133), .B2(new_n1242), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1241), .A2(new_n1216), .A3(new_n1246), .ZN(G407));
  NOR2_X1   g1047(.A1(new_n1241), .A2(new_n691), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1216), .A2(new_n1246), .ZN(new_n1249));
  OAI21_X1  g1049(.A(G213), .B1(new_n1248), .B2(new_n1249), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n687), .A2(G343), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G378), .B(new_n1215), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1181), .A2(new_n1184), .A3(new_n1236), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1215), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1252), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1124), .A2(new_n1098), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(KEYINPUT60), .A3(new_n1183), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n714), .A3(new_n1125), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT60), .B1(new_n1258), .B2(new_n1183), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1234), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G384), .B(new_n1234), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1252), .A2(G2897), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1251), .B1(new_n1257), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1266), .B(new_n1252), .C1(new_n1253), .C2(new_n1256), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(KEYINPUT125), .B(new_n1251), .C1(new_n1257), .C2(new_n1271), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1266), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1252), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1274), .A2(new_n1278), .A3(new_n1279), .A4(new_n1284), .ZN(new_n1285));
  XOR2_X1   g1085(.A(G393), .B(G396), .Z(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1239), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1003), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1009), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n969), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1025), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1090), .B1(new_n1292), .B2(new_n968), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1288), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(G390), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(G393), .B(G396), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1287), .A4(new_n1239), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1285), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(KEYINPUT63), .B2(new_n1276), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT63), .B1(new_n1257), .B2(new_n1271), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1301), .B2(new_n1283), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(G405));
  OAI21_X1  g1104(.A(new_n1253), .B1(new_n1216), .B2(new_n1245), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(KEYINPUT127), .B2(new_n1281), .ZN(new_n1306));
  XOR2_X1   g1106(.A(new_n1266), .B(KEYINPUT127), .Z(new_n1307));
  OAI211_X1 g1107(.A(new_n1307), .B(new_n1253), .C1(new_n1216), .C2(new_n1245), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1298), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1298), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


