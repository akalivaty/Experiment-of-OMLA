//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n203), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n215), .A2(new_n217), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n223), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n222), .A2(new_n224), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT25), .B1(new_n220), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT23), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n237), .B1(new_n219), .B2(new_n213), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n221), .B(new_n230), .C1(new_n227), .C2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n225), .B2(new_n226), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n236), .B(new_n238), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT68), .B1(new_n232), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n219), .A2(new_n213), .ZN(new_n245));
  INV_X1    g044(.A(new_n217), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT65), .B1(new_n216), .B2(KEYINPUT23), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n231), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n237), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n242), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n213), .A2(KEYINPUT26), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n235), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n218), .B(new_n254), .C1(new_n255), .C2(KEYINPUT26), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n225), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G183gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(new_n229), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n229), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n258), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n262), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n267), .A2(KEYINPUT71), .B1(KEYINPUT28), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n258), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n265), .B1(new_n264), .B2(new_n229), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n257), .B1(new_n269), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n209), .B1(new_n253), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n257), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n268), .A2(KEYINPUT28), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n273), .B2(new_n274), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n209), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n244), .A4(new_n252), .ZN(new_n284));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n277), .A2(new_n284), .A3(new_n285), .A4(new_n287), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n292));
  XOR2_X1   g091(.A(G15gat), .B(G43gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G71gat), .B(G99gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n285), .B1(new_n277), .B2(new_n284), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(KEYINPUT33), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n277), .A2(new_n284), .ZN(new_n301));
  INV_X1    g100(.A(new_n285), .ZN(new_n302));
  AOI221_X4 g101(.A(new_n298), .B1(KEYINPUT33), .B2(new_n295), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n292), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT33), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n308), .A3(new_n295), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n297), .A2(new_n299), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n289), .B2(new_n290), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n202), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n291), .B1(new_n300), .B2(new_n303), .ZN(new_n316));
  INV_X1    g115(.A(new_n291), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(new_n310), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n314), .A2(new_n315), .B1(new_n319), .B2(new_n202), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n313), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT74), .ZN(new_n323));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT0), .ZN(new_n325));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  INV_X1    g128(.A(G141gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G148gat), .ZN(new_n331));
  INV_X1    g130(.A(G148gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G141gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n331), .A2(new_n333), .B1(KEYINPUT2), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT77), .A3(new_n334), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT77), .B1(new_n336), .B2(new_n334), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n329), .B(new_n335), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n333), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n334), .A2(KEYINPUT2), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n339), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n337), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(new_n334), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT78), .B1(new_n335), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n283), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT84), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n283), .A2(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n348), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n209), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n207), .A2(KEYINPUT80), .A3(new_n208), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n367));
  INV_X1    g166(.A(new_n346), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n329), .B1(new_n343), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n370), .A2(KEYINPUT79), .A3(KEYINPUT3), .A4(new_n340), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n362), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n348), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n348), .A2(new_n374), .A3(new_n375), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT83), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n375), .ZN(new_n381));
  AOI211_X1 g180(.A(KEYINPUT82), .B(new_n381), .C1(new_n370), .C2(new_n340), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n376), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n383), .A2(new_n372), .A3(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n356), .B(new_n359), .C1(new_n380), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n358), .B1(new_n353), .B2(new_n350), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n373), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n384), .B1(new_n383), .B2(new_n372), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n366), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n352), .B1(new_n393), .B2(new_n348), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n358), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT6), .B(new_n328), .C1(new_n387), .C2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n386), .B(new_n327), .C1(new_n392), .C2(new_n396), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n390), .A2(new_n391), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n388), .ZN(new_n403));
  INV_X1    g202(.A(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n327), .B1(new_n405), .B2(new_n386), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n398), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  NAND2_X1  g209(.A1(new_n250), .A2(new_n242), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n282), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT22), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n417), .A2(KEYINPUT75), .B1(G211gat), .B2(G218gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(KEYINPUT75), .B2(new_n417), .ZN(new_n419));
  XNOR2_X1  g218(.A(G197gat), .B(G204gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G211gat), .B(G218gat), .Z(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT76), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n282), .A2(new_n414), .A3(new_n244), .A4(new_n252), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n282), .A2(new_n244), .A3(new_n252), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n415), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n282), .A2(new_n414), .A3(new_n411), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n424), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n410), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n410), .ZN(new_n433));
  INV_X1    g232(.A(new_n412), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n434), .A2(new_n414), .B1(new_n428), .B2(new_n415), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n426), .B(new_n433), .C1(new_n435), .C2(new_n424), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(KEYINPUT30), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(new_n410), .C1(new_n427), .C2(new_n431), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n407), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT88), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n423), .B(KEYINPUT76), .Z(new_n445));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n382), .B2(new_n376), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n423), .A2(new_n446), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n370), .B(new_n340), .C1(new_n449), .C2(new_n381), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n444), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT3), .B1(new_n423), .B2(new_n446), .ZN(new_n452));
  OAI211_X1 g251(.A(G228gat), .B(G233gat), .C1(new_n452), .C2(new_n348), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n445), .B2(new_n447), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G22gat), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT89), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(G50gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT86), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n455), .B2(new_n456), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(G22gat), .C1(new_n451), .C2(new_n454), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n462), .B(KEYINPUT87), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n455), .A2(new_n456), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n451), .A2(G22gat), .A3(new_n454), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n320), .A2(new_n323), .B1(new_n441), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n394), .A2(new_n358), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n390), .A2(new_n391), .B1(new_n354), .B2(new_n355), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT39), .B(new_n474), .C1(new_n475), .C2(new_n357), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n402), .A2(new_n356), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n358), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n327), .B(KEYINPUT90), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n440), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT40), .A4(new_n481), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n480), .B1(new_n387), .B2(new_n397), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n400), .A3(new_n399), .ZN(new_n489));
  INV_X1    g288(.A(new_n432), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n433), .A2(KEYINPUT37), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n436), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n435), .B2(new_n424), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n416), .A2(new_n425), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n445), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT38), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n490), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n436), .A2(new_n491), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n427), .A2(new_n431), .A3(new_n493), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT38), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n489), .A2(new_n498), .A3(new_n398), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n488), .A2(new_n502), .A3(new_n471), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n471), .A2(new_n321), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT35), .B1(new_n441), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT35), .B1(new_n489), .B2(new_n398), .ZN(new_n506));
  INV_X1    g305(.A(new_n319), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n506), .A2(new_n440), .A3(new_n471), .A4(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n473), .A2(new_n503), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT13), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G8gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT16), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G1gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n516), .B2(KEYINPUT96), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(G1gat), .B2(new_n514), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI221_X1 g318(.A(new_n516), .B1(KEYINPUT96), .B2(new_n513), .C1(G1gat), .C2(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(G43gat), .A2(G50gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(G43gat), .A2(G50gat), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT15), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(KEYINPUT92), .A2(G29gat), .A3(G36gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n528), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(KEYINPUT93), .A2(G50gat), .ZN(new_n538));
  INV_X1    g337(.A(G43gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT93), .A2(G50gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n541), .A2(KEYINPUT94), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT94), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n537), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n536), .ZN(new_n546));
  INV_X1    g345(.A(new_n531), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n537), .B(new_n549), .C1(new_n543), .C2(new_n544), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n522), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n528), .A2(new_n531), .A3(new_n536), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  INV_X1    g354(.A(new_n540), .ZN(new_n556));
  NOR2_X1   g355(.A1(KEYINPUT93), .A2(G50gat), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n556), .A2(new_n557), .A3(G43gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n541), .A2(KEYINPUT94), .A3(new_n542), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT95), .B1(new_n546), .B2(new_n547), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n552), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n521), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n512), .B1(new_n553), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n552), .B(new_n567), .C1(new_n562), .C2(new_n563), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n551), .B2(new_n552), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n522), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n510), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n572), .B1(new_n564), .B2(new_n521), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n564), .A2(KEYINPUT17), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n521), .B1(new_n577), .B2(new_n568), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n510), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT97), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581));
  AOI211_X1 g380(.A(new_n575), .B(new_n572), .C1(new_n564), .C2(new_n521), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n571), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G169gat), .B(G197gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT12), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n576), .A2(new_n584), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n576), .B2(new_n584), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT97), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n581), .B1(new_n571), .B2(new_n582), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n573), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n575), .B1(new_n578), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n566), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n595), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n576), .A2(new_n584), .A3(new_n590), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT98), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n594), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n509), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(G71gat), .A2(G78gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G57gat), .B(G64gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT9), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT99), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n617), .A3(new_n614), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n612), .A2(KEYINPUT100), .A3(new_n616), .A4(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(G57gat), .A2(G64gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(G57gat), .A2(G64gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G71gat), .B(G78gat), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n616), .A2(new_n622), .A3(new_n623), .A4(new_n618), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n614), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(KEYINPUT21), .ZN(new_n630));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n624), .A2(new_n625), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n624), .A2(new_n625), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n522), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n632), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT101), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n638), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT102), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT103), .ZN(new_n650));
  XOR2_X1   g449(.A(G134gat), .B(G162gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654));
  INV_X1    g453(.A(G99gat), .ZN(new_n655));
  INV_X1    g454(.A(G106gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G99gat), .A2(G106gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G85gat), .A2(G92gat), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT7), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(KEYINPUT8), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(G85gat), .B2(G92gat), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n654), .B(new_n659), .C1(new_n662), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n654), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n660), .B(KEYINPUT7), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n657), .A2(KEYINPUT104), .A3(new_n658), .ZN(new_n668));
  INV_X1    g467(.A(G85gat), .ZN(new_n669));
  INV_X1    g468(.A(G92gat), .ZN(new_n670));
  AOI22_X1  g469(.A1(KEYINPUT8), .A2(new_n658), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n666), .A2(new_n667), .A3(new_n668), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n577), .B2(new_n568), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n646), .A2(new_n647), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n564), .B2(new_n673), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(G190gat), .B(G218gat), .Z(new_n678));
  NOR3_X1   g477(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  INV_X1    g479(.A(new_n673), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n569), .B2(new_n570), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n682), .B2(new_n676), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n653), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n680), .A3(new_n676), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(new_n652), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(G230gat), .A2(G233gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT106), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n627), .A2(new_n628), .A3(new_n673), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n673), .B1(new_n627), .B2(new_n628), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT105), .B(KEYINPUT10), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n627), .A2(new_n628), .A3(new_n673), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT10), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n691), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n636), .A2(new_n681), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n691), .B1(new_n701), .B2(new_n697), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(G120gat), .B(G148gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(G176gat), .B(G204gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(new_n706));
  NAND3_X1  g505(.A1(new_n700), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n706), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n701), .A2(new_n697), .A3(new_n694), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n692), .A2(KEYINPUT10), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n690), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n711), .B2(new_n702), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n712), .A3(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n714), .B(new_n708), .C1(new_n711), .C2(new_n702), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n645), .A2(new_n688), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n607), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n407), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g521(.A1(new_n718), .A2(new_n440), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT108), .B(KEYINPUT16), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(new_n513), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n725), .ZN(new_n729));
  INV_X1    g528(.A(new_n723), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n730), .A2(KEYINPUT109), .A3(G8gat), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT109), .B1(new_n730), .B2(G8gat), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n728), .B(new_n729), .C1(new_n731), .C2(new_n732), .ZN(G1325gat));
  NAND2_X1  g532(.A1(new_n320), .A2(new_n323), .ZN(new_n734));
  OAI21_X1  g533(.A(G15gat), .B1(new_n718), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n319), .A2(G15gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n718), .B2(new_n736), .ZN(G1326gat));
  NOR2_X1   g536(.A1(new_n718), .A2(new_n471), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT43), .B(G22gat), .Z(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1327gat));
  INV_X1    g539(.A(new_n645), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n716), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n688), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n607), .A2(new_n524), .A3(new_n720), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT45), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n509), .B2(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n441), .A2(new_n472), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n503), .A2(new_n734), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n505), .A2(new_n508), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n688), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n591), .A2(new_n592), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n743), .A2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n755), .A2(new_n720), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n747), .B1(new_n524), .B2(new_n758), .ZN(G1328gat));
  NOR2_X1   g558(.A1(new_n440), .A2(G36gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n607), .A2(new_n745), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT46), .Z(new_n762));
  NAND4_X1  g561(.A1(new_n749), .A2(new_n754), .A3(new_n485), .A4(new_n757), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G36gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(KEYINPUT110), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n761), .B(KEYINPUT46), .ZN(new_n767));
  INV_X1    g566(.A(new_n764), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n765), .A2(new_n769), .ZN(G1329gat));
  INV_X1    g569(.A(new_n734), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n755), .A2(G43gat), .A3(new_n771), .A4(new_n757), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n607), .A2(new_n745), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n539), .B1(new_n773), .B2(new_n319), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(new_n777), .A3(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1330gat));
  AOI21_X1  g578(.A(new_n471), .B1(new_n538), .B2(new_n540), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n755), .A2(new_n757), .A3(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n538), .B(new_n540), .C1(new_n773), .C2(new_n471), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g583(.A(new_n716), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n603), .A2(new_n604), .ZN(new_n786));
  NOR4_X1   g585(.A1(new_n645), .A2(new_n785), .A3(new_n786), .A4(new_n688), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n753), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n407), .ZN(new_n789));
  XNOR2_X1  g588(.A(KEYINPUT111), .B(G57gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1332gat));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n440), .ZN(new_n792));
  NOR2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n792), .B2(new_n793), .ZN(G1333gat));
  NOR3_X1   g595(.A1(new_n788), .A2(G71gat), .A3(new_n319), .ZN(new_n797));
  INV_X1    g596(.A(new_n788), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n771), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(G71gat), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n472), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g602(.A1(new_n741), .A2(new_n786), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n716), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT112), .Z(new_n806));
  NAND2_X1  g605(.A1(new_n755), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G85gat), .B1(new_n807), .B2(new_n407), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n753), .A2(new_n688), .A3(new_n804), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n744), .B1(new_n751), .B2(new_n752), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n804), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n720), .A2(new_n669), .A3(new_n716), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n808), .B1(new_n815), .B2(new_n816), .ZN(G1336gat));
  NOR3_X1   g616(.A1(new_n440), .A2(new_n785), .A3(G92gat), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n749), .A2(new_n754), .A3(new_n485), .A4(new_n806), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n814), .A2(new_n818), .B1(new_n819), .B2(G92gat), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n819), .B2(G92gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n820), .A2(KEYINPUT52), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n809), .A2(new_n810), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT51), .B1(new_n812), .B2(new_n804), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n818), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n819), .A2(G92gat), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n826), .B(new_n827), .C1(KEYINPUT113), .C2(KEYINPUT52), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n823), .A2(new_n829), .ZN(G1337gat));
  OAI21_X1  g629(.A(G99gat), .B1(new_n807), .B2(new_n734), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n507), .A2(new_n655), .A3(new_n716), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n815), .B2(new_n832), .ZN(G1338gat));
  NAND4_X1  g632(.A1(new_n749), .A2(new_n754), .A3(new_n472), .A4(new_n806), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n656), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n471), .A2(G106gat), .A3(new_n785), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n814), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n834), .A2(G106gat), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n838), .B(KEYINPUT114), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n815), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(G1339gat));
  NOR4_X1   g644(.A1(new_n645), .A2(new_n786), .A3(new_n688), .A4(new_n716), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n709), .A2(new_n690), .A3(new_n710), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n700), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n706), .B1(new_n711), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n850), .A3(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n707), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n848), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n510), .B1(new_n571), .B2(new_n565), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n553), .A2(new_n565), .A3(new_n512), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n589), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n604), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n688), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n854), .A2(new_n786), .B1(new_n858), .B2(new_n716), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(new_n688), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n846), .B1(new_n861), .B2(new_n645), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n407), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n504), .A2(new_n485), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n786), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n863), .A2(new_n440), .A3(new_n471), .A4(new_n507), .ZN(new_n868));
  INV_X1    g667(.A(G113gat), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n868), .A2(new_n869), .A3(new_n606), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n867), .A2(new_n870), .ZN(G1340gat));
  AOI21_X1  g670(.A(G120gat), .B1(new_n866), .B2(new_n716), .ZN(new_n872));
  INV_X1    g671(.A(G120gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n868), .A2(new_n873), .A3(new_n785), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n868), .B2(new_n645), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n645), .A2(G127gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n865), .B2(new_n877), .ZN(G1342gat));
  OAI21_X1  g677(.A(G134gat), .B1(new_n868), .B2(new_n744), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT116), .Z(new_n880));
  NOR3_X1   g679(.A1(new_n865), .A2(G134gat), .A3(new_n744), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT56), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1343gat));
  NAND2_X1  g682(.A1(new_n734), .A2(new_n472), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n485), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n863), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n606), .A2(G141gat), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n471), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n848), .A2(new_n850), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT55), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n707), .A3(new_n851), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n756), .A2(KEYINPUT98), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n786), .A2(new_n593), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n604), .A2(new_n713), .A3(new_n715), .A4(new_n857), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n744), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n741), .B1(new_n902), .B2(new_n859), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n892), .B1(new_n903), .B2(new_n846), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n891), .B1(new_n862), .B2(new_n471), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n734), .A2(new_n720), .A3(new_n440), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G141gat), .B1(new_n909), .B2(new_n606), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT58), .B1(new_n890), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n906), .A2(KEYINPUT117), .A3(new_n908), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT58), .B(G141gat), .C1(new_n915), .C2(new_n756), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n888), .B1(new_n889), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n911), .B1(new_n916), .B2(new_n918), .ZN(G1344gat));
  NAND3_X1  g718(.A1(new_n886), .A2(new_n332), .A3(new_n716), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G148gat), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n913), .A2(new_n914), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n716), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n741), .A2(new_n756), .A3(new_n744), .A4(new_n785), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n688), .A2(new_n604), .A3(new_n857), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n896), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n900), .B1(new_n896), .B2(new_n756), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n744), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n929), .B2(new_n741), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n892), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n854), .B1(new_n594), .B2(new_n605), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n688), .B1(new_n932), .B2(new_n900), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n645), .B1(new_n933), .B2(new_n927), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n717), .A2(new_n606), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n471), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n931), .B1(new_n936), .B2(KEYINPUT57), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n716), .A3(new_n908), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n921), .B1(new_n938), .B2(G148gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n920), .B1(new_n924), .B2(new_n939), .ZN(G1345gat));
  OAI21_X1  g739(.A(G155gat), .B1(new_n915), .B2(new_n645), .ZN(new_n941));
  INV_X1    g740(.A(new_n886), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n645), .A2(G155gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1346gat));
  OAI21_X1  g743(.A(G162gat), .B1(new_n915), .B2(new_n744), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n744), .A2(G162gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n942), .B2(new_n946), .ZN(G1347gat));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n862), .B2(new_n720), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n930), .A2(KEYINPUT119), .A3(new_n407), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n504), .A2(new_n440), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G169gat), .B1(new_n954), .B2(new_n786), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n472), .A2(new_n440), .A3(new_n319), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n930), .A2(new_n407), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT120), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n958), .A2(new_n211), .A3(new_n606), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n955), .A2(new_n959), .ZN(G1348gat));
  OAI21_X1  g759(.A(G176gat), .B1(new_n958), .B2(new_n785), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n785), .A2(G176gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n961), .B1(new_n953), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT121), .Z(G1349gat));
  OAI21_X1  g764(.A(G183gat), .B1(new_n958), .B2(new_n645), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n741), .A2(new_n264), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n953), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n229), .A3(new_n688), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n958), .A2(new_n744), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n972), .A2(new_n973), .A3(G190gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n972), .B2(G190gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1351gat));
  NOR2_X1   g775(.A1(new_n884), .A2(new_n440), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n951), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n786), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n771), .A2(new_n720), .A3(new_n440), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n937), .A2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(G197gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n606), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(G1352gat));
  NAND3_X1  g784(.A1(new_n937), .A2(new_n716), .A3(new_n981), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT124), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n937), .A2(new_n988), .A3(new_n716), .A4(new_n981), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n987), .A2(G204gat), .A3(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n991), .A2(KEYINPUT123), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n785), .A2(G204gat), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n734), .A2(new_n485), .A3(new_n472), .A4(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT122), .B1(new_n951), .B2(new_n995), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT122), .ZN(new_n997));
  AOI211_X1 g796(.A(new_n997), .B(new_n994), .C1(new_n949), .C2(new_n950), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n992), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n862), .A2(new_n948), .A3(new_n720), .ZN(new_n1000));
  AOI21_X1  g799(.A(KEYINPUT119), .B1(new_n930), .B2(new_n407), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n995), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(new_n997), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n951), .A2(KEYINPUT122), .A3(new_n995), .ZN(new_n1004));
  XNOR2_X1  g803(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT125), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n990), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1353gat));
  OR3_X1    g811(.A1(new_n978), .A2(G211gat), .A3(new_n645), .ZN(new_n1013));
  OAI21_X1  g812(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1014), .B1(new_n982), .B2(new_n741), .ZN(new_n1015));
  AND2_X1   g814(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(G1354gat));
  INV_X1    g818(.A(G218gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1020), .B1(new_n978), .B2(new_n744), .ZN(new_n1021));
  OR2_X1    g820(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n744), .A2(new_n1020), .ZN(new_n1024));
  AOI22_X1  g823(.A1(new_n1022), .A2(new_n1023), .B1(new_n982), .B2(new_n1024), .ZN(G1355gat));
endmodule


