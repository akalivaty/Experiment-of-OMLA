//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n548, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  OR4_X1    g030(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n462), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G113), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT68), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G113), .A3(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n471), .B(new_n473), .C1(new_n466), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n467), .A2(G136), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n463), .A2(new_n465), .A3(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n483), .B2(G112), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT69), .Z(G162));
  NAND4_X1  g061(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n483), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G138), .A4(new_n483), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT70), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n480), .A2(G126), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n492), .A2(new_n500), .A3(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n514), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  AND2_X1   g097(.A1(new_n511), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  INV_X1    g099(.A(new_n518), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n524), .A2(new_n526), .A3(new_n527), .A4(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(G90), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n523), .A2(new_n532), .B1(new_n525), .B2(G52), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT75), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AOI22_X1  g114(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n513), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n542), .A2(new_n543), .B1(G43), .B2(new_n525), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n523), .A2(G81), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT77), .Z(G188));
  NAND2_X1  g128(.A1(new_n525), .A2(G53), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n523), .A2(G91), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n511), .A2(G65), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT78), .Z(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n556), .A3(new_n560), .ZN(G299));
  NAND2_X1  g136(.A1(new_n523), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n525), .A2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n513), .ZN(new_n567));
  INV_X1    g142(.A(G86), .ZN(new_n568));
  INV_X1    g143(.A(G48), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n516), .A2(new_n568), .B1(new_n518), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n513), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  INV_X1    g151(.A(G47), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n516), .A2(new_n576), .B1(new_n518), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n575), .A2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n523), .A2(G92), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT10), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n513), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n525), .A2(G54), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n580), .B1(new_n587), .B2(G868), .ZN(G284));
  XOR2_X1   g163(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g164(.A1(G286), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G299), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(G868), .ZN(G297));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(G868), .ZN(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G860), .ZN(G148));
  NOR2_X1   g170(.A1(new_n546), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n585), .A2(new_n586), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(G559), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n596), .B1(new_n599), .B2(G868), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n489), .A2(new_n468), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT13), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(G2100), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n467), .A2(G135), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n480), .A2(G123), .ZN(new_n608));
  OR2_X1    g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G2104), .C1(G111), .C2(new_n483), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n606), .A2(new_n612), .ZN(G156));
  XNOR2_X1  g188(.A(KEYINPUT15), .B(G2435), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT81), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2427), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT14), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2451), .B(G2454), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n619), .B(new_n625), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n626), .A2(G14), .ZN(G401));
  XOR2_X1   g202(.A(G2084), .B(G2090), .Z(new_n628));
  XNOR2_X1  g203(.A(G2067), .B(G2678), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n630), .A2(KEYINPUT17), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT18), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n630), .B2(KEYINPUT18), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2096), .B(G2100), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(G227));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n639));
  XOR2_X1   g214(.A(G1961), .B(G1966), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(new_n641));
  XOR2_X1   g216(.A(G1956), .B(G2474), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1971), .B(G1976), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT19), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n641), .A2(new_n642), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n648), .A2(new_n645), .A3(new_n643), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n643), .A2(new_n639), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n650), .A2(new_n647), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n646), .B(new_n649), .C1(new_n651), .C2(new_n645), .ZN(new_n652));
  XOR2_X1   g227(.A(G1991), .B(G1996), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1981), .B(G1986), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G229));
  NOR2_X1   g233(.A1(G29), .A2(G33), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n467), .A2(G139), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n468), .A2(G103), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT25), .Z(new_n662));
  AOI22_X1  g237(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT87), .Z(new_n664));
  OAI211_X1 g239(.A(new_n660), .B(new_n662), .C1(new_n664), .C2(new_n483), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT88), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n659), .B1(new_n667), .B2(G29), .ZN(new_n668));
  NAND2_X1  g243(.A1(KEYINPUT91), .A2(G2072), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(KEYINPUT24), .A2(G34), .ZN(new_n671));
  INV_X1    g246(.A(G29), .ZN(new_n672));
  NAND2_X1  g247(.A1(KEYINPUT24), .A2(G34), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G160), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT89), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G2084), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT90), .ZN(new_n678));
  NOR2_X1   g253(.A1(KEYINPUT91), .A2(G2072), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n467), .A2(G141), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT92), .ZN(new_n682));
  NAND3_X1  g257(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT26), .Z(new_n684));
  AOI22_X1  g259(.A1(new_n480), .A2(G129), .B1(G105), .B2(new_n468), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT93), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G29), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n692), .B(KEYINPUT94), .C1(G29), .C2(G32), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(KEYINPUT94), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT27), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT95), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n670), .B(new_n680), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT96), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n672), .A2(G26), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n467), .A2(G140), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n480), .A2(G128), .ZN(new_n701));
  OR2_X1    g276(.A1(G104), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G116), .C2(new_n483), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n672), .ZN(new_n706));
  MUX2_X1   g281(.A(new_n699), .B(new_n706), .S(KEYINPUT28), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT86), .B(G2067), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G290), .A2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G24), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT83), .B1(new_n711), .B2(G16), .ZN(new_n712));
  OR3_X1    g287(.A1(new_n711), .A2(KEYINPUT83), .A3(G16), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1986), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(G6), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n571), .B2(new_n716), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT32), .B(G1981), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT84), .B1(G16), .B2(G23), .ZN(new_n725));
  OR3_X1    g300(.A1(KEYINPUT84), .A2(G16), .A3(G23), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(G288), .C2(new_n716), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT33), .B(G1976), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n720), .A2(new_n724), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n715), .B1(new_n730), .B2(KEYINPUT34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n467), .A2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n480), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(new_n483), .B2(G107), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G25), .B(new_n736), .S(G29), .Z(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT35), .B(G1991), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n737), .B(new_n738), .Z(new_n739));
  OAI211_X1 g314(.A(new_n731), .B(new_n739), .C1(KEYINPUT34), .C2(new_n730), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(KEYINPUT85), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n676), .A2(G2084), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT97), .ZN(new_n745));
  NAND2_X1  g320(.A1(G171), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G5), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n716), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n716), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1966), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT30), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n611), .B2(new_n672), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n745), .A2(new_n749), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n694), .A2(new_n696), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT31), .B(G11), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n716), .A2(G19), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n546), .B2(new_n716), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n747), .A2(new_n748), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n716), .A2(G20), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT99), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G299), .B2(G16), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G1956), .Z(new_n768));
  NOR3_X1   g343(.A1(new_n762), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n672), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n672), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT29), .Z(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT98), .ZN(new_n776));
  NOR2_X1   g351(.A1(G27), .A2(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G164), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2078), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n716), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n587), .B2(new_n716), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n773), .B2(new_n774), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n770), .A2(new_n776), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n698), .A2(new_n709), .A3(new_n743), .A4(new_n785), .ZN(G150));
  INV_X1    g361(.A(G150), .ZN(G311));
  AOI22_X1  g362(.A1(new_n523), .A2(G93), .B1(new_n525), .B2(G55), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n513), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT100), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G860), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT37), .Z(new_n794));
  NOR2_X1   g369(.A1(new_n597), .A2(new_n594), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n546), .A2(new_n790), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n544), .A2(new_n545), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n797), .B(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n794), .B1(new_n802), .B2(G860), .ZN(G145));
  XNOR2_X1  g378(.A(G162), .B(new_n477), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n688), .A2(new_n501), .A3(new_n689), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n501), .B1(new_n688), .B2(new_n689), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n807), .A2(new_n704), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n497), .A2(new_n499), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n488), .B2(new_n491), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n690), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n705), .B1(new_n814), .B2(new_n806), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n667), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n704), .B1(new_n807), .B2(new_n808), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n705), .A3(new_n806), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n817), .A2(new_n665), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n611), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n611), .B1(new_n816), .B2(new_n819), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n736), .B(new_n604), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n467), .A2(G142), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n480), .A2(G130), .ZN(new_n825));
  NOR2_X1   g400(.A1(G106), .A2(G2105), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(new_n483), .B2(G118), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n823), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n821), .A2(new_n822), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n611), .ZN(new_n832));
  INV_X1    g407(.A(new_n819), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n666), .B1(new_n817), .B2(new_n818), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n829), .B1(new_n835), .B2(new_n820), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n805), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G37), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n830), .B1(new_n821), .B2(new_n822), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n829), .A3(new_n820), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n804), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n837), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT101), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n837), .A2(new_n844), .A3(new_n838), .A4(new_n841), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n843), .A2(KEYINPUT40), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT40), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(G395));
  XNOR2_X1  g423(.A(G290), .B(G288), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT105), .ZN(new_n850));
  XNOR2_X1  g425(.A(G303), .B(KEYINPUT104), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G305), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(KEYINPUT105), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT42), .ZN(new_n857));
  OR2_X1    g432(.A1(G299), .A2(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g433(.A1(G299), .A2(KEYINPUT102), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n587), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n597), .A2(KEYINPUT102), .A3(G299), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT103), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n860), .A2(KEYINPUT41), .A3(new_n861), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT41), .B1(new_n860), .B2(new_n861), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n798), .A2(new_n800), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n599), .ZN(new_n868));
  MUX2_X1   g443(.A(new_n863), .B(new_n866), .S(new_n868), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n857), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(G868), .B2(new_n791), .ZN(G295));
  OAI21_X1  g447(.A(new_n871), .B1(G868), .B2(new_n791), .ZN(G331));
  XNOR2_X1  g448(.A(G301), .B(G168), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n801), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n867), .A2(new_n874), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(KEYINPUT107), .A3(new_n877), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n867), .A2(new_n874), .A3(KEYINPUT107), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n861), .A3(new_n860), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n866), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n866), .A3(KEYINPUT106), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n856), .ZN(new_n888));
  INV_X1    g463(.A(new_n856), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n881), .A2(new_n885), .A3(new_n889), .A4(new_n886), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n838), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT43), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n878), .A2(new_n866), .A3(new_n879), .ZN(new_n893));
  INV_X1    g468(.A(new_n863), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n882), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n856), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n890), .A2(new_n896), .A3(new_n838), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n888), .A2(new_n903), .A3(new_n838), .A4(new_n890), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n904), .A3(KEYINPUT44), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(G397));
  XOR2_X1   g483(.A(KEYINPUT113), .B(G8), .Z(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(G168), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n469), .A2(new_n476), .A3(G40), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n813), .B2(G1384), .ZN(new_n916));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n501), .A2(KEYINPUT110), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT50), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G2084), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n492), .A2(new_n500), .A3(KEYINPUT71), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT71), .B1(new_n492), .B2(new_n500), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n923), .A2(new_n924), .A3(G1384), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT111), .B1(new_n925), .B2(new_n920), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n503), .A2(new_n917), .A3(new_n504), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT50), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n921), .A2(new_n922), .A3(new_n926), .A4(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n916), .A2(new_n931), .A3(new_n918), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n917), .A4(new_n504), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n913), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1966), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n912), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n909), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT120), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(KEYINPUT120), .A3(new_n909), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n912), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G8), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n930), .B2(new_n936), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT51), .B1(new_n946), .B2(new_n911), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n937), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT126), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n942), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n910), .B1(new_n930), .B2(new_n936), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n912), .B1(new_n952), .B2(KEYINPUT120), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n947), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n937), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT126), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n914), .B1(new_n916), .B2(new_n918), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n910), .ZN(new_n961));
  INV_X1    g536(.A(G288), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G1976), .ZN(new_n963));
  INV_X1    g538(.A(G1976), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT52), .B1(G288), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G305), .A2(G1981), .ZN(new_n967));
  INV_X1    g542(.A(G1981), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n571), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT49), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(KEYINPUT49), .A3(new_n969), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n961), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT110), .B1(new_n501), .B2(new_n917), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n915), .B(G1384), .C1(new_n492), .C2(new_n500), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n913), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n909), .A3(new_n963), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT52), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n978), .B2(KEYINPUT52), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n966), .B(new_n974), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n925), .B2(KEYINPUT45), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n501), .A2(new_n917), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n913), .B1(new_n990), .B2(new_n931), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n927), .A2(KEYINPUT109), .A3(new_n931), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n916), .A2(KEYINPUT50), .A3(new_n918), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n503), .A2(new_n920), .A3(new_n917), .A4(new_n504), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n995), .A2(new_n913), .A3(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n994), .A2(new_n719), .B1(new_n997), .B2(new_n774), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n987), .B1(new_n998), .B2(new_n910), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n921), .A2(new_n774), .A3(new_n926), .A4(new_n929), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n927), .A2(KEYINPUT109), .A3(new_n931), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT109), .B1(new_n927), .B2(new_n931), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n991), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1003), .B2(G1971), .ZN(new_n1004));
  OR3_X1    g579(.A1(new_n985), .A2(KEYINPUT112), .A3(new_n986), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT112), .B1(new_n985), .B2(new_n986), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n983), .A2(new_n999), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT123), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT123), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n983), .A2(new_n999), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n954), .A2(new_n949), .A3(new_n955), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n921), .A2(new_n926), .A3(new_n929), .ZN(new_n1015));
  INV_X1    g590(.A(G2078), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n989), .A2(new_n1016), .A3(new_n992), .A4(new_n993), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n748), .A2(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n932), .A2(new_n1016), .A3(new_n913), .A4(new_n933), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1018), .B1(new_n1020), .B2(KEYINPUT121), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(KEYINPUT121), .B2(new_n1020), .ZN(new_n1022));
  AOI21_X1  g597(.A(G301), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  AND4_X1   g598(.A1(KEYINPUT125), .A2(new_n1013), .A3(new_n1014), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G171), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT125), .B1(new_n1027), .B2(new_n1014), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n959), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT127), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n974), .A2(new_n964), .A3(new_n962), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n969), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n961), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1008), .B2(new_n982), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT63), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n952), .A2(G168), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1009), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1004), .A2(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1041), .B2(new_n987), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n1008), .A3(new_n983), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1040), .B1(new_n1043), .B2(new_n1039), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1037), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT56), .B(G2072), .Z(new_n1046));
  OAI22_X1  g621(.A1(new_n994), .A2(new_n1046), .B1(new_n997), .B2(G1956), .ZN(new_n1047));
  XNOR2_X1  g622(.A(G299), .B(KEYINPUT57), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G2067), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1015), .A2(new_n782), .B1(new_n1050), .B2(new_n960), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT116), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(new_n587), .C1(new_n1048), .C2(new_n1047), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n587), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1051), .B(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1055), .A2(new_n1058), .B1(new_n1054), .B2(new_n1052), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(G1996), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1003), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1003), .A2(KEYINPUT118), .A3(new_n1060), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT58), .B(G1341), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1063), .B(new_n1064), .C1(new_n960), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n546), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n1070), .A2(KEYINPUT119), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(KEYINPUT59), .A3(new_n546), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1070), .B1(KEYINPUT119), .B2(new_n1071), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1049), .B(new_n1053), .C1(new_n1059), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n990), .A2(new_n931), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n992), .A2(KEYINPUT53), .A3(new_n1016), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1019), .A2(G301), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1081), .B2(new_n1023), .ZN(new_n1082));
  AOI22_X1  g657(.A1(KEYINPUT122), .A2(new_n1082), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1015), .A2(new_n748), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1079), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1019), .A2(new_n1022), .A3(G301), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(KEYINPUT54), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n1026), .B2(new_n1080), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1092), .A2(new_n1093), .B1(new_n954), .B2(new_n955), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1083), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1045), .B1(new_n1076), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n959), .B(KEYINPUT127), .C1(new_n1024), .C2(new_n1028), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1031), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1078), .A2(new_n914), .ZN(new_n1099));
  INV_X1    g674(.A(G1996), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n691), .A2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n736), .A2(new_n738), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n704), .B(new_n1050), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n690), .A2(G1996), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n738), .B2(new_n736), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G290), .A2(G1986), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G290), .A2(G1986), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1099), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1098), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT46), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1099), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(G1996), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1099), .A2(KEYINPUT46), .A3(new_n1100), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n691), .A2(new_n1103), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1114), .B(new_n1115), .C1(new_n1116), .C2(new_n1113), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT47), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1109), .A2(new_n1099), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT48), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1122), .A2(new_n1102), .B1(G2067), .B2(new_n704), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1099), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1118), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1111), .A2(new_n1125), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g701(.A1(new_n843), .A2(new_n845), .ZN(new_n1128));
  INV_X1    g702(.A(G319), .ZN(new_n1129));
  OR2_X1    g703(.A1(G229), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g704(.A(new_n1130), .B1(new_n892), .B2(new_n898), .ZN(new_n1131));
  NOR2_X1   g705(.A1(G401), .A2(G227), .ZN(new_n1132));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .ZN(G225));
  INV_X1    g707(.A(G225), .ZN(G308));
endmodule


