//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT10), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT65), .B1(new_n191), .B2(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(new_n191), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT65), .A3(G143), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n190), .B1(new_n194), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n200), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n188), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n201), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(G107), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n218));
  XNOR2_X1  g032(.A(G104), .B(G107), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT78), .A3(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n187), .B1(new_n207), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n233), .A3(new_n236), .A4(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n209), .A2(new_n212), .A3(new_n214), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n215), .A2(new_n216), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n215), .A2(new_n216), .ZN(new_n243));
  OAI211_X1 g057(.A(KEYINPUT4), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  OR2_X1    g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n196), .A2(new_n198), .A3(new_n191), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(new_n204), .ZN(new_n249));
  INV_X1    g063(.A(new_n246), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n202), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n243), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n215), .A2(new_n216), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n224), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n195), .B2(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n258), .B(new_n191), .C1(new_n196), .C2(new_n198), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n189), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  OAI21_X1  g077(.A(G128), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n248), .A2(new_n204), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n256), .A2(new_n267), .A3(KEYINPUT10), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n227), .A2(new_n239), .A3(new_n253), .A4(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G110), .B(G140), .ZN(new_n270));
  INV_X1    g084(.A(G227), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n270), .B(new_n272), .Z(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT79), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n227), .A2(new_n253), .A3(new_n268), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n238), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT79), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n269), .A2(new_n278), .A3(new_n273), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n262), .B1(new_n202), .B2(new_n205), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n256), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n202), .A2(new_n189), .B1(new_n264), .B2(new_n265), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n226), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT12), .B1(new_n285), .B2(new_n238), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n287), .B(new_n239), .C1(new_n282), .C2(new_n284), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n269), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n273), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n280), .A2(new_n291), .A3(G469), .ZN(new_n292));
  INV_X1    g106(.A(G469), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT70), .B(G902), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n286), .ZN(new_n296));
  INV_X1    g110(.A(new_n288), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n274), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n273), .B1(new_n277), .B2(new_n269), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n293), .B(new_n295), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n292), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G221), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT76), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n307), .B2(new_n301), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(KEYINPUT80), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(G125), .A2(G140), .ZN(new_n315));
  NOR2_X1   g129(.A1(G125), .A2(G140), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT16), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G125), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(G146), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n320), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n195), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n317), .A2(new_n325), .A3(G146), .A4(new_n320), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G237), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G214), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n191), .ZN(new_n332));
  NOR2_X1   g146(.A1(G237), .A2(G953), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(G143), .A3(G214), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT87), .B1(new_n335), .B2(G131), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(G131), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT87), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n332), .A2(new_n339), .A3(new_n236), .A4(new_n334), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n336), .A2(new_n337), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(KEYINPUT17), .A3(G131), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n328), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n208), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n345), .B(KEYINPUT89), .Z(new_n346));
  XNOR2_X1  g160(.A(G125), .B(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n199), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n195), .B2(new_n347), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT18), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(new_n236), .ZN(new_n351));
  OAI221_X1 g165(.A(new_n349), .B1(new_n335), .B2(new_n351), .C1(new_n338), .C2(new_n350), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n343), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n345), .B1(new_n343), .B2(new_n352), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n301), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT91), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT91), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(new_n301), .C1(new_n353), .C2(new_n354), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(G475), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(G475), .A2(G902), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT88), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n347), .A2(new_n361), .A3(KEYINPUT19), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT19), .B1(new_n347), .B2(new_n361), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n321), .B1(new_n365), .B2(new_n193), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n336), .A2(new_n338), .A3(new_n340), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n352), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n345), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n343), .A2(new_n346), .A3(new_n352), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n370), .A2(KEYINPUT90), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT90), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  OAI211_X1 g187(.A(KEYINPUT20), .B(new_n360), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n360), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n359), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT92), .ZN(new_n380));
  INV_X1    g194(.A(G478), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(KEYINPUT15), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n191), .A2(G128), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n188), .A2(G143), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n229), .ZN(new_n386));
  INV_X1    g200(.A(G116), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT14), .A3(G122), .ZN(new_n388));
  XNOR2_X1  g202(.A(G116), .B(G122), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(G107), .B(new_n388), .C1(new_n390), .C2(KEYINPUT14), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n386), .B(new_n391), .C1(G107), .C2(new_n390), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n229), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n389), .B(new_n211), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT13), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT93), .B1(new_n383), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(new_n395), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT93), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n398), .A2(new_n191), .A3(KEYINPUT13), .A4(G128), .ZN(new_n399));
  AND4_X1   g213(.A1(new_n384), .A2(new_n396), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n393), .B(new_n394), .C1(new_n400), .C2(new_n229), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n307), .A2(G217), .A3(new_n330), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n405));
  INV_X1    g219(.A(new_n403), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n392), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n406), .A2(KEYINPUT94), .A3(new_n401), .A4(new_n392), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n295), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n382), .B1(new_n410), .B2(KEYINPUT95), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(KEYINPUT95), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(new_n382), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n359), .A2(new_n374), .A3(new_n414), .A4(new_n378), .ZN(new_n415));
  OR2_X1    g229(.A1(KEYINPUT96), .A2(G952), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT96), .A2(G952), .ZN(new_n417));
  AOI21_X1  g231(.A(G953), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G234), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n329), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n294), .B(G953), .C1(new_n419), .C2(new_n329), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT21), .B(G898), .Z(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n380), .A2(new_n413), .A3(new_n415), .A4(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G214), .B1(G237), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G125), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT82), .B1(new_n251), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n283), .A2(new_n428), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n246), .B1(new_n194), .B2(new_n200), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n431), .B(G125), .C1(new_n432), .C2(new_n249), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n330), .A2(G224), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT83), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n429), .A2(new_n436), .A3(new_n430), .A4(new_n433), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  INV_X1    g255(.A(G119), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G116), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n387), .A2(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G116), .B(G119), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT68), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT2), .B(G113), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n445), .A2(new_n451), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n244), .A2(new_n454), .A3(new_n252), .ZN(new_n455));
  OAI21_X1  g269(.A(G113), .B1(new_n443), .B2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT5), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n450), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n217), .A2(new_n459), .A3(new_n453), .A4(new_n225), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT81), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n441), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n455), .B2(new_n460), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT6), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n440), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n436), .A2(KEYINPUT7), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n429), .A2(new_n430), .A3(new_n433), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n466), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n262), .A2(new_n428), .A3(new_n266), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n202), .A2(new_n250), .ZN(new_n477));
  INV_X1    g291(.A(new_n249), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n428), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n472), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n445), .A2(new_n458), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n453), .B1(new_n481), .B2(new_n456), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n217), .A2(new_n225), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n462), .B(KEYINPUT8), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n459), .A2(new_n453), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n256), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n301), .B1(new_n475), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(new_n301), .C1(new_n475), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n466), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT6), .B1(new_n493), .B2(new_n468), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n465), .A2(new_n441), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n440), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n471), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT86), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n471), .A2(new_n492), .A3(new_n498), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n427), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n314), .A2(new_n425), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n507));
  NOR2_X1   g321(.A1(G472), .A2(G902), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n509));
  INV_X1    g323(.A(new_n231), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n229), .A2(G137), .ZN(new_n511));
  OAI21_X1  g325(.A(G131), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n237), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT67), .B1(new_n267), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n516), .B(new_n513), .C1(new_n262), .C2(new_n266), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n477), .A2(new_n238), .A3(new_n478), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT66), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n251), .A2(new_n521), .A3(new_n238), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n509), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n267), .A2(new_n514), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n525), .A2(new_n519), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT30), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n454), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n454), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n333), .A2(G210), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(new_n213), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n528), .A2(new_n537), .A3(new_n530), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR4_X1   g353(.A1(new_n239), .A2(new_n432), .A3(KEYINPUT66), .A4(new_n249), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n521), .B1(new_n251), .B2(new_n238), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n516), .B1(new_n283), .B2(new_n513), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n267), .A2(KEYINPUT67), .A3(new_n514), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n529), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n530), .B1(new_n546), .B2(KEYINPUT69), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n548), .B(new_n529), .C1(new_n542), .C2(new_n545), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT28), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n530), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT28), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n534), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n508), .B1(new_n539), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT32), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT32), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n557), .B(new_n508), .C1(new_n539), .C2(new_n554), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n550), .A2(new_n553), .A3(new_n534), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n528), .A2(new_n530), .ZN(new_n560));
  INV_X1    g374(.A(new_n534), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT29), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n525), .A2(new_n519), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n454), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n530), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(KEYINPUT28), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n552), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(KEYINPUT29), .A3(new_n534), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(new_n295), .A3(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n556), .A2(new_n558), .B1(G472), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n188), .A2(KEYINPUT71), .A3(G119), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n188), .A2(G119), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT71), .B1(new_n188), .B2(G119), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(KEYINPUT24), .A2(G110), .ZN(new_n576));
  NOR2_X1   g390(.A1(KEYINPUT24), .A2(G110), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n442), .B2(G128), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n442), .A2(G128), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G110), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n327), .A2(new_n579), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n574), .A2(new_n573), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n188), .A2(KEYINPUT71), .A3(G119), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n578), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G110), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n581), .A2(new_n583), .A3(new_n590), .A4(new_n582), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT73), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT73), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n594), .B(new_n591), .C1(new_n575), .C2(new_n578), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n593), .A2(new_n595), .A3(new_n321), .A4(new_n348), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT74), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n586), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT22), .B(G137), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n305), .A2(new_n419), .A3(G953), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n597), .B1(new_n586), .B2(new_n596), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n597), .B(new_n601), .C1(new_n586), .C2(new_n596), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n295), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT25), .ZN(new_n607));
  INV_X1    g421(.A(G217), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n295), .B2(G234), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT25), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n610), .B(new_n295), .C1(new_n604), .C2(new_n605), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(G902), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n604), .A2(new_n605), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n507), .B1(new_n571), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n570), .A2(G472), .ZN(new_n618));
  INV_X1    g432(.A(new_n558), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n454), .B1(new_n518), .B2(new_n523), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n548), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n546), .A2(KEYINPUT69), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n530), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n552), .B1(new_n623), .B2(KEYINPUT28), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n538), .B(new_n536), .C1(new_n624), .C2(new_n534), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n557), .B1(new_n625), .B2(new_n508), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n618), .B1(new_n619), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n616), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT75), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n506), .B1(new_n617), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n213), .ZN(G3));
  OAI21_X1  g445(.A(new_n295), .B1(new_n539), .B2(new_n554), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n632), .A2(new_n633), .A3(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n632), .B2(G472), .ZN(new_n635));
  INV_X1    g449(.A(new_n555), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n304), .A2(KEYINPUT80), .A3(new_n309), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT80), .B1(new_n304), .B2(new_n309), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n638), .A2(new_n616), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT98), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n502), .A2(KEYINPUT99), .A3(new_n504), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n503), .A2(new_n471), .A3(new_n492), .A4(new_n498), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n427), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n380), .A2(new_n415), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n404), .A2(new_n651), .A3(new_n407), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n402), .A2(KEYINPUT100), .A3(new_n403), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n408), .A2(new_n409), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n655), .B2(new_n650), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n294), .A2(new_n381), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n656), .A2(new_n657), .B1(new_n381), .B2(new_n410), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n423), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n648), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  OAI21_X1  g479(.A(new_n360), .B1(new_n372), .B2(new_n373), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n377), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n374), .A3(new_n359), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n413), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n648), .A2(new_n423), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT35), .B(G107), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n670), .B(new_n673), .ZN(G9));
  OAI21_X1  g488(.A(new_n505), .B1(new_n639), .B2(new_n640), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n424), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n586), .A2(new_n596), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n601), .A2(KEYINPUT36), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n613), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n612), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n677), .B1(new_n612), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n676), .A2(new_n637), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G12));
  NAND3_X1  g501(.A1(new_n684), .A2(new_n647), .A3(new_n644), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n571), .A2(new_n641), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n420), .B1(new_n421), .B2(G900), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n413), .A2(new_n668), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT104), .B(G128), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G30));
  NOR2_X1   g509(.A1(new_n684), .A2(new_n427), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n556), .A2(new_n558), .ZN(new_n697));
  INV_X1    g511(.A(new_n535), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n561), .B2(new_n566), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n699), .B2(G902), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n502), .A2(new_n504), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n413), .B1(new_n380), .B2(new_n415), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n690), .B(KEYINPUT39), .Z(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n314), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT106), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n696), .B(new_n706), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  AND3_X1   g528(.A1(new_n684), .A2(new_n647), .A3(new_n644), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n691), .B(new_n658), .C1(new_n380), .C2(new_n415), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n627), .A2(new_n715), .A3(new_n314), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n697), .A2(new_n618), .B1(new_n312), .B2(new_n313), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(KEYINPUT107), .A3(new_n715), .A4(new_n716), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  INV_X1    g537(.A(new_n299), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n269), .B(new_n273), .C1(new_n286), .C2(new_n288), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n293), .B1(new_n726), .B2(new_n295), .ZN(new_n727));
  INV_X1    g541(.A(new_n300), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n308), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n647), .A2(new_n644), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n628), .A2(new_n731), .A3(new_n627), .A4(new_n662), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT41), .B(G113), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND2_X1  g548(.A1(new_n669), .A2(new_n423), .ZN(new_n735));
  NOR4_X1   g549(.A1(new_n571), .A2(new_n730), .A3(new_n616), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n387), .ZN(G18));
  AOI21_X1  g551(.A(new_n424), .B1(new_n697), .B2(new_n618), .ZN(new_n738));
  INV_X1    g552(.A(new_n729), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n688), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  INV_X1    g556(.A(G472), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n625), .B2(new_n295), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n561), .B1(new_n567), .B2(new_n552), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n536), .A2(new_n745), .A3(new_n538), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n508), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n744), .A2(new_n747), .A3(new_n616), .A4(new_n661), .ZN(new_n748));
  AND4_X1   g562(.A1(new_n644), .A2(new_n647), .A3(new_n705), .A4(new_n729), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NAND2_X1  g565(.A1(new_n632), .A2(G472), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n746), .A2(new_n508), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n683), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n612), .A2(new_n677), .A3(new_n681), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n716), .A4(new_n731), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n716), .A2(new_n752), .A3(new_n684), .A4(new_n753), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n761), .B2(new_n730), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n571), .B2(new_n616), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n304), .A2(KEYINPUT109), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n292), .A2(new_n300), .A3(new_n768), .A4(new_n303), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n309), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n649), .A2(new_n659), .A3(new_n690), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n502), .A2(new_n426), .A3(new_n504), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n627), .A2(KEYINPUT110), .A3(new_n628), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n770), .A2(new_n773), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n627), .A2(new_n777), .A3(new_n628), .A4(new_n716), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n772), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  AND4_X1   g595(.A1(new_n628), .A2(new_n627), .A3(new_n777), .A4(new_n692), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n229), .ZN(G36));
  AND3_X1   g597(.A1(new_n280), .A2(new_n291), .A3(KEYINPUT45), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT45), .B1(new_n280), .B2(new_n291), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT46), .B(new_n303), .C1(new_n786), .C2(new_n293), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n300), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n784), .A2(new_n785), .A3(new_n293), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(new_n792), .B2(new_n302), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT112), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n787), .A2(KEYINPUT111), .A3(new_n300), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(KEYINPUT112), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n790), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n309), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n707), .ZN(new_n799));
  INV_X1    g613(.A(new_n773), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n380), .A2(new_n659), .A3(new_n415), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n638), .A2(KEYINPUT44), .A3(new_n684), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT44), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n684), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n637), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n799), .A2(new_n800), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n798), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n771), .A2(new_n773), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n627), .A2(new_n628), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NOR2_X1   g631(.A1(new_n727), .A2(new_n728), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n427), .B1(new_n819), .B2(KEYINPUT49), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n309), .C1(KEYINPUT49), .C2(new_n819), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n697), .A2(new_n628), .A3(new_n700), .ZN(new_n822));
  OR4_X1    g636(.A1(new_n704), .A2(new_n821), .A3(new_n822), .A4(new_n801), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n630), .A2(new_n732), .A3(new_n736), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n782), .B1(new_n776), .B2(new_n779), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n738), .A2(new_n740), .B1(new_n748), .B2(new_n749), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n702), .A2(new_n423), .A3(new_n426), .ZN(new_n829));
  INV_X1    g643(.A(new_n413), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n415), .A3(new_n380), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n660), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n637), .A2(new_n832), .A3(new_n628), .A4(new_n314), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n828), .A2(new_n833), .A3(new_n685), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n761), .A2(new_n773), .A3(new_n770), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n757), .A2(new_n668), .A3(new_n691), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n773), .A2(new_n830), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n627), .A2(new_n836), .A3(new_n314), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT113), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n720), .A2(new_n840), .A3(new_n837), .A4(new_n836), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n835), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n826), .A2(new_n827), .A3(new_n834), .A4(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n760), .A2(new_n762), .B1(new_n689), .B2(new_n692), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n612), .A2(new_n681), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n697), .B2(new_n700), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n647), .A2(new_n705), .A3(new_n644), .ZN(new_n847));
  INV_X1    g661(.A(new_n770), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n846), .A2(new_n690), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n722), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n844), .A2(new_n722), .A3(new_n849), .A4(KEYINPUT52), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n843), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n825), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n853), .ZN(new_n857));
  INV_X1    g671(.A(new_n843), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n855), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(KEYINPUT118), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n851), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n850), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n858), .A3(KEYINPUT53), .A4(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n824), .A2(new_n856), .A3(new_n861), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n857), .A2(new_n858), .A3(new_n855), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n854), .A2(KEYINPUT117), .A3(new_n855), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n863), .A2(new_n858), .A3(new_n864), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n866), .B1(KEYINPUT54), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n420), .B1(new_n803), .B2(new_n804), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n754), .A2(new_n616), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n819), .A2(new_n309), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n800), .B(new_n881), .C1(new_n813), .C2(new_n882), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n739), .A2(new_n420), .A3(new_n773), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n884), .A2(new_n822), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n885), .A2(new_n649), .A3(new_n659), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n427), .A3(new_n729), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(new_n887), .B2(new_n704), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT50), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT50), .ZN(new_n890));
  OAI211_X1 g704(.A(KEYINPUT119), .B(new_n890), .C1(new_n887), .C2(new_n704), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n884), .B1(new_n804), .B2(new_n803), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n758), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n883), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT51), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n883), .A2(new_n892), .A3(new_n897), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n766), .A2(new_n775), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n893), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT48), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n885), .A2(new_n660), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n418), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n731), .B2(new_n881), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n899), .A2(KEYINPUT120), .A3(new_n905), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n878), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n823), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NAND3_X1  g726(.A1(new_n856), .A2(new_n861), .A3(new_n865), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n913), .A2(new_n294), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n501), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n496), .B(new_n440), .Z(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n915), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n330), .A2(G952), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G51));
  XOR2_X1   g736(.A(new_n726), .B(KEYINPUT121), .Z(new_n923));
  NAND2_X1  g737(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n856), .A2(new_n861), .A3(new_n824), .A4(new_n865), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n302), .B(KEYINPUT57), .Z(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n914), .A2(new_n792), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(G54));
  NAND3_X1  g745(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n372), .A2(new_n373), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n921), .ZN(G60));
  INV_X1    g750(.A(new_n656), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n926), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n921), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(KEYINPUT122), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n937), .B1(new_n878), .B2(new_n939), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  INV_X1    g759(.A(new_n940), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n924), .B2(new_n925), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n945), .B1(new_n947), .B2(new_n921), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n943), .A2(new_n944), .A3(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT60), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n913), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n615), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n913), .A2(new_n680), .A3(new_n951), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n942), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT61), .B1(new_n954), .B2(KEYINPUT123), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G66));
  AOI21_X1  g771(.A(new_n330), .B1(new_n422), .B2(G224), .ZN(new_n958));
  INV_X1    g772(.A(new_n826), .ZN(new_n959));
  INV_X1    g773(.A(new_n834), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n958), .B1(new_n962), .B2(new_n330), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n494), .B(new_n495), .C1(G898), .C2(new_n330), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(G69));
  NAND2_X1  g779(.A1(new_n844), .A2(new_n722), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n810), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n799), .A2(new_n847), .A3(new_n900), .ZN(new_n971));
  INV_X1    g785(.A(new_n827), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(G953), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n970), .A2(new_n816), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n271), .B2(new_n330), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n524), .A2(new_n527), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(new_n365), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n977), .A2(G227), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n330), .B1(new_n979), .B2(G900), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n617), .A2(new_n629), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n773), .B1(new_n660), .B2(new_n831), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n710), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT124), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n983), .A2(KEYINPUT124), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n810), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  INV_X1    g801(.A(new_n816), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n713), .A2(new_n967), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n713), .A2(KEYINPUT62), .A3(new_n967), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n977), .A2(G953), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n980), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n978), .A2(new_n996), .ZN(G72));
  NAND3_X1  g811(.A1(new_n987), .A2(new_n993), .A3(new_n961), .ZN(new_n998));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n560), .B(KEYINPUT127), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1001), .A2(new_n534), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n962), .A2(new_n972), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n970), .A2(new_n816), .A3(new_n1005), .A4(new_n971), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n1000), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n561), .A3(new_n1002), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1004), .A2(new_n1008), .A3(new_n942), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n560), .A2(new_n561), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n535), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n877), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1009), .B1(new_n1000), .B2(new_n1012), .ZN(G57));
endmodule


