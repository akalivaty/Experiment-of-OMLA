//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT66), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n211), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  OR2_X1    g0024(.A1(KEYINPUT65), .A2(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(KEYINPUT65), .A2(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n203), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n209), .B(new_n224), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n221), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  INV_X1    g0042(.A(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n246), .B(KEYINPUT68), .Z(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n220), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT10), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT70), .B(G1698), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(G222), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G223), .A3(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(new_n255), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(G274), .C1(G41), .C2(G45), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT69), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G226), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n263), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G200), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT75), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT74), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n270), .A2(KEYINPUT75), .A3(G200), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n273), .A2(new_n275), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  INV_X1    g0079(.A(G20), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n279), .A2(new_n280), .A3(G1), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT72), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR3_X1   g0087(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G150), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n291), .B(G20), .C1(new_n201), .C2(new_n203), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(G33), .A3(new_n227), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n285), .A2(new_n290), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n228), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n283), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n264), .B2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G50), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n273), .A2(new_n277), .A3(new_n275), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n253), .B(new_n278), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n273), .A2(new_n277), .A3(new_n275), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(new_n305), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n309), .B(new_n310), .C1(new_n276), .C2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n270), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n302), .B(new_n313), .C1(G179), .C2(new_n270), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n308), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  INV_X1    g0116(.A(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G33), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n318), .A2(new_n320), .A3(G232), .A4(G1698), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n318), .B(new_n320), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n316), .B(new_n321), .C1(new_n324), .C2(new_n221), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n262), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n268), .A2(G238), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n266), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(KEYINPUT76), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n330), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n326), .A2(new_n327), .A3(new_n266), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(G179), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n328), .A2(new_n329), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n326), .A2(KEYINPUT13), .A3(new_n327), .A4(new_n266), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G169), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n337), .A2(new_n341), .A3(G169), .A4(new_n338), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n331), .A2(KEYINPUT77), .A3(G179), .A4(new_n333), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n336), .A2(new_n340), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G68), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G20), .ZN(new_n346));
  AND2_X1   g0146(.A1(KEYINPUT65), .A2(G20), .ZN(new_n347));
  NOR2_X1   g0147(.A1(KEYINPUT65), .A2(G20), .ZN(new_n348));
  OAI211_X1 g0148(.A(G33), .B(G77), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n287), .A2(new_n288), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n346), .B(new_n349), .C1(new_n350), .C2(new_n220), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n298), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT11), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n281), .A2(new_n345), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n298), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n300), .A2(G68), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n354), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n344), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n337), .A2(G200), .A3(new_n338), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n331), .A2(G190), .A3(new_n333), .ZN(new_n362));
  INV_X1    g0162(.A(new_n359), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n315), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n282), .A2(new_n293), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n300), .B2(new_n293), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n298), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n250), .A2(new_n345), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n202), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n350), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT78), .B1(new_n317), .B2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT78), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(new_n319), .A3(G33), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n377), .A3(new_n318), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n280), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT7), .B1(new_n225), .B2(new_n226), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n379), .A2(KEYINPUT7), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n374), .B1(new_n381), .B2(G68), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n370), .B1(new_n382), .B2(KEYINPUT16), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n319), .B2(G33), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n317), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n320), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n255), .B2(G20), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n345), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n384), .B1(new_n392), .B2(new_n374), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n369), .B1(new_n383), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n268), .A2(G232), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n317), .A2(new_n212), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G226), .A2(G1698), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n322), .A2(new_n323), .ZN(new_n398));
  INV_X1    g0198(.A(G223), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n375), .A2(new_n377), .A3(new_n318), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n266), .B(new_n395), .C1(new_n402), .C2(new_n261), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G169), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n254), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n405), .A2(new_n378), .B1(new_n317), .B2(new_n212), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n262), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(G179), .A3(new_n266), .A4(new_n395), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT80), .B(KEYINPUT18), .C1(new_n394), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n379), .A2(KEYINPUT7), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n378), .A2(new_n380), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(G68), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n374), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(new_n298), .A3(new_n393), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n368), .ZN(new_n418));
  NOR2_X1   g0218(.A1(KEYINPUT80), .A2(KEYINPUT18), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(KEYINPUT80), .A2(KEYINPUT18), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n418), .A2(new_n409), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT81), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n403), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n407), .A2(new_n274), .A3(new_n266), .A4(new_n395), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n417), .A3(new_n368), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n424), .A2(new_n425), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n426), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n394), .B2(new_n430), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n411), .B(new_n423), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT82), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n282), .A2(G77), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(G33), .A3(new_n227), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n347), .A2(new_n348), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G77), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n444), .C1(new_n350), .C2(new_n293), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(new_n445), .B2(new_n298), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n300), .A2(G77), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n266), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n254), .A2(new_n255), .A3(G232), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n243), .C2(new_n255), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n452), .B2(new_n262), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n268), .A2(G244), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n448), .B(KEYINPUT73), .C1(new_n455), .C2(G169), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT73), .ZN(new_n457));
  AOI21_X1  g0257(.A(G169), .B1(new_n453), .B2(new_n454), .ZN(new_n458));
  INV_X1    g0258(.A(new_n447), .ZN(new_n459));
  AOI211_X1 g0259(.A(new_n439), .B(new_n459), .C1(new_n445), .C2(new_n298), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G179), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n456), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n455), .A2(G190), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n460), .C1(new_n427), .C2(new_n455), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n436), .B2(new_n437), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n366), .A2(new_n438), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G274), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n261), .B(G250), .C1(G1), .C2(new_n471), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G116), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G244), .A2(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(G238), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n398), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(new_n401), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n473), .B(new_n474), .C1(new_n480), .C2(new_n261), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n312), .ZN(new_n482));
  OAI211_X1 g0282(.A(G33), .B(G97), .C1(new_n347), .C2(new_n348), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n212), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n316), .A2(new_n484), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n443), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n227), .A2(new_n318), .A3(new_n375), .A4(new_n377), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n485), .B(new_n489), .C1(new_n490), .C2(new_n345), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n298), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n440), .A2(new_n281), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n264), .A2(G33), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n282), .A2(new_n370), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n441), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n254), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n475), .B1(new_n499), .B2(new_n378), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n262), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(new_n462), .A3(new_n473), .A4(new_n474), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n482), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(G87), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n492), .A2(new_n493), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n481), .A2(new_n427), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n501), .A2(new_n274), .A3(new_n473), .A4(new_n474), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n389), .A2(new_n391), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n243), .A2(KEYINPUT6), .A3(G97), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n214), .A2(new_n243), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(new_n486), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n443), .B1(new_n289), .B2(G77), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n298), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n282), .A2(G97), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n496), .B2(G97), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(G244), .B1(new_n322), .B2(new_n323), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT4), .B1(new_n401), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G283), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n318), .A2(new_n320), .A3(G250), .A4(G1698), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT4), .B(G244), .C1(new_n322), .C2(new_n323), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n318), .A2(new_n320), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n262), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(KEYINPUT5), .A2(G41), .ZN(new_n531));
  AND2_X1   g0331(.A1(KEYINPUT5), .A2(G41), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n472), .B(G274), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n472), .B1(new_n532), .B2(new_n531), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n261), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n535), .B2(new_n215), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n312), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n378), .B2(new_n522), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n526), .A2(new_n525), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n528), .C2(new_n527), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n536), .B1(new_n544), .B2(new_n262), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n540), .B1(new_n545), .B2(new_n462), .ZN(new_n546));
  AND4_X1   g0346(.A1(new_n540), .A2(new_n530), .A3(new_n462), .A4(new_n537), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n521), .B(new_n539), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT83), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n545), .B2(new_n427), .ZN(new_n550));
  INV_X1    g0350(.A(new_n520), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n517), .B2(new_n298), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(G190), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n538), .A2(KEYINPUT83), .A3(G200), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n509), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n534), .A2(G264), .A3(new_n261), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT89), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(G294), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n317), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G257), .A2(G1698), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n254), .B2(G250), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n565), .B2(new_n378), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n262), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(new_n533), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n563), .B1(new_n398), .B2(new_n213), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n561), .B1(new_n569), .B2(new_n401), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n533), .B(new_n557), .C1(new_n570), .C2(new_n261), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n427), .A2(new_n568), .B1(new_n572), .B2(new_n274), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT22), .B1(new_n255), .B2(G87), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n225), .A2(new_n575), .A3(new_n226), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n475), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n280), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n401), .A2(KEYINPUT22), .A3(G87), .A4(new_n227), .ZN(new_n582));
  NAND2_X1  g0382(.A1(KEYINPUT23), .A2(G107), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT24), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n581), .A2(new_n582), .A3(new_n586), .A4(new_n583), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n370), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n281), .A2(KEYINPUT25), .A3(new_n243), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT25), .B1(new_n281), .B2(new_n243), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n495), .B2(new_n243), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n573), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n559), .A2(G179), .A3(new_n533), .A4(new_n567), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n571), .A2(G169), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n588), .B2(new_n592), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT86), .ZN(new_n601));
  INV_X1    g0401(.A(G303), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n255), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(G257), .B1(new_n322), .B2(new_n323), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G264), .A2(G1698), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n606), .B2(new_n401), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n607), .B2(new_n261), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n528), .A2(G303), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n254), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n378), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(KEYINPUT86), .A3(new_n262), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n534), .A2(G270), .A3(new_n261), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n533), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT85), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n617), .A3(new_n533), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n317), .A2(G97), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n620), .B(new_n525), .C1(new_n347), .C2(new_n348), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n297), .A2(new_n228), .B1(G20), .B2(new_n245), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT88), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT88), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n282), .A2(G116), .A3(new_n370), .A4(new_n494), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n621), .A2(KEYINPUT88), .A3(new_n622), .A4(new_n624), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n264), .A2(new_n245), .A3(G13), .A4(G20), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT87), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n613), .A2(G179), .A3(new_n619), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n619), .A2(new_n608), .A3(new_n612), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  INV_X1    g0435(.A(new_n632), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n619), .A2(G190), .A3(new_n608), .A4(new_n612), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n632), .A2(G169), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n634), .A2(new_n639), .A3(KEYINPUT21), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n633), .A2(new_n638), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n470), .A2(new_n556), .A3(new_n600), .A4(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n314), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT18), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT90), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n418), .A2(new_n649), .A3(new_n409), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n418), .B2(new_n409), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n418), .A2(new_n409), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT90), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n418), .A2(new_n649), .A3(new_n409), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(KEYINPUT18), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n364), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n464), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n359), .B2(new_n344), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n433), .A2(new_n435), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n308), .A2(new_n311), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n647), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n482), .A2(new_n498), .A3(new_n502), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n597), .A2(new_n642), .A3(new_n633), .A4(new_n643), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n568), .A2(new_n427), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(G190), .B2(new_n571), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n588), .A2(new_n592), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n665), .B1(new_n671), .B2(new_n556), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n506), .A2(new_n507), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n665), .B1(new_n674), .B2(new_n505), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n675), .B2(new_n548), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT84), .B1(new_n538), .B2(G179), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n545), .A2(new_n540), .A3(new_n462), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n552), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n509), .A2(KEYINPUT26), .A3(new_n679), .A4(new_n539), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n672), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n664), .B1(new_n470), .B2(new_n682), .ZN(G369));
  NAND2_X1  g0483(.A1(new_n227), .A2(G13), .ZN(new_n684));
  OR3_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .A3(G1), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT27), .B1(new_n684), .B2(G1), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n644), .B1(new_n636), .B2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n634), .A2(new_n639), .A3(KEYINPUT21), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT21), .B1(new_n634), .B2(new_n639), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n619), .A2(G179), .A3(new_n608), .A4(new_n612), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n636), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n690), .A2(new_n636), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n599), .B1(new_n669), .B2(new_n690), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n597), .B2(new_n690), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n671), .A2(new_n689), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n207), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n487), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n230), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n593), .B1(new_n696), .B2(new_n597), .ZN(new_n718));
  INV_X1    g0518(.A(new_n556), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n503), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n676), .A2(new_n680), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n689), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n717), .B1(new_n722), .B2(KEYINPUT29), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n690), .B1(new_n672), .B2(new_n681), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(KEYINPUT91), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n718), .A2(new_n719), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT92), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n676), .A2(new_n680), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n548), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n509), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n728), .A2(new_n730), .A3(new_n665), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .A3(new_n690), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n719), .A2(new_n644), .A3(new_n599), .A4(new_n690), .ZN(new_n735));
  INV_X1    g0535(.A(new_n694), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n559), .A2(new_n567), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n538), .A2(new_n481), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n481), .A2(new_n462), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n538), .A3(new_n634), .A4(new_n568), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n736), .A2(KEYINPUT30), .A3(new_n737), .A4(new_n738), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n689), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n746), .A2(KEYINPUT31), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n727), .A2(new_n734), .B1(G330), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n716), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(new_n703), .ZN(new_n752));
  INV_X1    g0552(.A(new_n684), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n264), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n711), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n701), .A2(new_n702), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n752), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT93), .Z(new_n760));
  NOR4_X1   g0560(.A1(new_n227), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT102), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n427), .A2(G179), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n443), .A2(new_n274), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT100), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n763), .A2(G329), .B1(new_n770), .B2(G283), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT103), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n227), .A2(new_n462), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G317), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(KEYINPUT33), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(KEYINPUT33), .B2(new_n777), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(G190), .A3(new_n427), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G322), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n443), .A2(G179), .A3(new_n274), .A4(new_n427), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n255), .B1(new_n784), .B2(G311), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n779), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n774), .A2(new_n274), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n274), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n227), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n787), .A2(G326), .B1(G294), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT101), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n786), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n764), .A2(G20), .A3(G190), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n772), .B(new_n795), .C1(new_n602), .C2(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n776), .A2(new_n345), .B1(new_n769), .B2(new_n243), .ZN(new_n798));
  INV_X1    g0598(.A(new_n761), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT99), .B(G159), .Z(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(KEYINPUT32), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n214), .B2(new_n789), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n799), .A2(KEYINPUT32), .A3(new_n801), .ZN(new_n804));
  OR3_X1    g0604(.A1(new_n798), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G77), .B1(G58), .B2(new_n781), .ZN(new_n810));
  INV_X1    g0610(.A(new_n787), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n220), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n805), .B1(KEYINPUT98), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n813), .B1(KEYINPUT98), .B2(new_n812), .C1(new_n212), .C2(new_n796), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n797), .B1(new_n814), .B2(new_n528), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n312), .A2(KEYINPUT95), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n312), .A2(KEYINPUT95), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n816), .A2(new_n817), .A3(G20), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n818), .A2(G1), .A3(G13), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT96), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G13), .A2(G33), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n251), .A2(G45), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n401), .A2(new_n710), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G45), .C2(new_n230), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n710), .A2(new_n528), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT94), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G355), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n828), .B(new_n831), .C1(G116), .C2(new_n207), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n815), .A2(new_n821), .B1(new_n825), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n824), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n700), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n760), .B1(new_n757), .B2(new_n835), .ZN(G396));
  NOR2_X1   g0636(.A1(new_n690), .A2(new_n460), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n464), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n464), .B2(new_n466), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n724), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n749), .A2(G330), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n757), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G137), .A2(new_n787), .B1(new_n775), .B2(G150), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT104), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n780), .C1(new_n808), .C2(new_n801), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT34), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n770), .A2(G68), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n250), .B2(new_n789), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n401), .B1(new_n220), .B2(new_n796), .C1(new_n762), .C2(new_n854), .ZN(new_n855));
  OR4_X1    g0655(.A1(new_n850), .A2(new_n851), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G311), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n762), .A2(new_n857), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n780), .A2(new_n560), .B1(new_n214), .B2(new_n789), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n809), .B2(G116), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n770), .A2(G87), .B1(new_n787), .B2(G303), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n528), .B1(new_n796), .B2(new_n243), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n775), .B2(G283), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n856), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n821), .A2(new_n822), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n865), .A2(new_n821), .B1(new_n258), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n867), .B(new_n756), .C1(new_n823), .C2(new_n840), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n844), .A2(new_n868), .ZN(G384));
  NAND2_X1  g0669(.A1(new_n414), .A2(new_n415), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n384), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n369), .B1(new_n383), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n431), .B1(new_n872), .B2(new_n687), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n410), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n687), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n418), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n653), .A2(new_n877), .A3(new_n878), .A4(new_n431), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n872), .A2(new_n687), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n411), .A2(new_n423), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n661), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n875), .A2(KEYINPUT106), .A3(new_n879), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n877), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n431), .A2(new_n426), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n394), .A2(new_n430), .B1(new_n424), .B2(new_n425), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n426), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n652), .A3(new_n656), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n654), .A2(new_n655), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n877), .A2(new_n431), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n888), .A2(new_n892), .B1(new_n895), .B2(new_n879), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n887), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n359), .A2(new_n689), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT105), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n359), .A2(new_n900), .A3(new_n689), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n658), .B(new_n902), .C1(new_n344), .C2(new_n359), .ZN(new_n903));
  INV_X1    g0703(.A(new_n902), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n360), .B2(new_n364), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AND4_X1   g0706(.A1(new_n747), .A2(new_n906), .A3(new_n748), .A4(new_n840), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n897), .A2(new_n907), .A3(KEYINPUT40), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n747), .A2(new_n906), .A3(new_n748), .A4(new_n840), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n885), .A2(new_n886), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT106), .B1(new_n875), .B2(new_n879), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n911), .B1(new_n887), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n910), .B1(new_n916), .B2(KEYINPUT40), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n887), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n907), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(KEYINPUT107), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n909), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n469), .A2(new_n749), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G330), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n360), .A2(new_n689), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n918), .A2(KEYINPUT39), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n887), .B(new_n929), .C1(new_n896), .C2(KEYINPUT38), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n903), .A2(new_n905), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n690), .B(new_n840), .C1(new_n672), .C2(new_n681), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n464), .A2(new_n689), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n918), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n657), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n687), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n723), .A2(new_n469), .A3(new_n734), .A4(new_n726), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n664), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n925), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n264), .B2(new_n753), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n245), .B1(new_n515), .B2(KEYINPUT35), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n946), .B(new_n229), .C1(KEYINPUT35), .C2(new_n515), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT36), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n230), .A2(new_n258), .A3(new_n371), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n201), .A2(new_n345), .ZN(new_n950));
  OAI211_X1 g0750(.A(G1), .B(new_n279), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n945), .A2(new_n948), .A3(new_n951), .ZN(G367));
  INV_X1    g0752(.A(KEYINPUT112), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n521), .A2(new_n689), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n539), .A2(new_n679), .B1(new_n555), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n548), .A2(new_n689), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n955), .A2(KEYINPUT109), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT109), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT45), .B1(new_n959), .B2(new_n708), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(KEYINPUT45), .A3(new_n708), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT44), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n959), .B2(new_n708), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n957), .A2(KEYINPUT44), .A3(new_n707), .A4(new_n958), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n961), .A2(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT110), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n706), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n965), .ZN(new_n969));
  INV_X1    g0769(.A(new_n962), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n970), .B2(new_n960), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n971), .A2(KEYINPUT110), .A3(new_n703), .A4(new_n705), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n696), .A2(new_n689), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n705), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT111), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n973), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n600), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT111), .B1(new_n705), .B2(new_n973), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n703), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n752), .A2(new_n976), .A3(new_n979), .A4(new_n980), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n968), .A2(new_n972), .A3(new_n750), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n750), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n711), .B(KEYINPUT41), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n755), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n505), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n509), .B1(new_n989), .B2(new_n690), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n503), .A2(new_n505), .A3(new_n689), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT108), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n959), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT42), .B1(new_n996), .B2(new_n979), .ZN(new_n997));
  INV_X1    g0797(.A(new_n956), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n959), .A2(new_n598), .A3(new_n690), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT42), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n959), .A2(new_n1000), .A3(new_n978), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n703), .A2(new_n705), .A3(new_n959), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1003), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n995), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1007), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(new_n994), .A3(new_n1005), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n953), .B1(new_n988), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1011), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n987), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n985), .B2(new_n750), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1013), .B(KEYINPUT112), .C1(new_n755), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n770), .A2(G77), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n255), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT113), .Z(new_n1020));
  AOI22_X1  g0820(.A1(G143), .A2(new_n787), .B1(new_n775), .B2(new_n800), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n796), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n790), .A2(G68), .B1(G58), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(G150), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1023), .C1(new_n1024), .C2(new_n780), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n201), .B2(new_n809), .ZN(new_n1026));
  INV_X1    g0826(.A(G137), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1020), .B(new_n1026), .C1(new_n1027), .C2(new_n799), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n789), .A2(new_n243), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n776), .A2(new_n560), .B1(new_n769), .B2(new_n214), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G311), .B2(new_n787), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT46), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n796), .B2(new_n245), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1022), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n799), .C2(new_n777), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n401), .B(new_n1035), .C1(G303), .C2(new_n781), .ZN(new_n1036));
  INV_X1    g0836(.A(G283), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1031), .B(new_n1036), .C1(new_n1037), .C2(new_n808), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1028), .B1(new_n1029), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT47), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n821), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n827), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n825), .B1(new_n207), .B2(new_n440), .C1(new_n239), .C2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n990), .A2(new_n824), .A3(new_n991), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n756), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1017), .A2(new_n1045), .ZN(G387));
  OR2_X1    g0846(.A1(new_n750), .A2(new_n984), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n750), .A2(new_n984), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n711), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G311), .A2(new_n775), .B1(new_n787), .B2(G322), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n777), .B2(new_n780), .C1(new_n602), .C2(new_n808), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT48), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n1037), .B2(new_n789), .C1(new_n560), .C2(new_n796), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT49), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n761), .A2(G326), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n401), .B1(new_n770), .B2(G116), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n780), .A2(new_n220), .B1(new_n345), .B2(new_n783), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n789), .A2(new_n440), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n796), .A2(new_n258), .ZN(new_n1060));
  OR3_X1    g0860(.A1(new_n1059), .A2(new_n378), .A3(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1058), .B(new_n1061), .C1(G150), .C2(new_n761), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n770), .A2(G97), .B1(new_n787), .B2(G159), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n293), .C2(new_n776), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n820), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n293), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1066));
  OAI21_X1  g0866(.A(KEYINPUT50), .B1(new_n293), .B2(G50), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n471), .A4(new_n713), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G68), .B2(G77), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n827), .B1(new_n236), .B2(new_n471), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n830), .B1(G116), .B2(new_n487), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n207), .A2(G107), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n825), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n705), .B2(new_n834), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1065), .A2(new_n757), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n755), .B2(new_n984), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1049), .A2(new_n1077), .ZN(G393));
  XNOR2_X1  g0878(.A(new_n966), .B(new_n706), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1079), .A2(new_n754), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n775), .A2(G303), .B1(G116), .B2(new_n790), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n560), .B2(new_n783), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT114), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n255), .B1(new_n1022), .B2(G283), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n811), .A2(new_n777), .B1(new_n857), .B2(new_n780), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n770), .A2(G107), .B1(G322), .B2(new_n761), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT115), .Z(new_n1089));
  OAI22_X1  g0889(.A1(new_n811), .A2(new_n1024), .B1(new_n373), .B2(new_n780), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n770), .A2(G87), .B1(new_n775), .B2(new_n201), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n789), .A2(new_n258), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n401), .B1(new_n345), .B2(new_n796), .C1(new_n799), .C2(new_n847), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n809), .C2(new_n294), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1091), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n820), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n959), .A2(new_n834), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n246), .A2(new_n1042), .B1(new_n214), .B2(new_n207), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1099), .A2(new_n824), .A3(new_n821), .ZN(new_n1100));
  NOR4_X1   g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n757), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1080), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1079), .A2(new_n1048), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n711), .A3(new_n985), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  NAND4_X1  g0906(.A1(new_n747), .A2(new_n748), .A3(G330), .A4(new_n840), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n932), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n930), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n933), .A2(new_n934), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n926), .B1(new_n1110), .B2(new_n906), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n929), .B1(new_n915), .B2(new_n887), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n897), .A2(new_n927), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n733), .A2(new_n690), .A3(new_n840), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n932), .B1(new_n1115), .B2(new_n934), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1108), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n928), .B(new_n930), .C1(new_n926), .C2(new_n935), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1107), .A2(new_n932), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1115), .A2(new_n934), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n927), .B(new_n897), .C1(new_n1121), .C2(new_n932), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1118), .A2(new_n755), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1118), .A2(new_n1123), .A3(KEYINPUT116), .A4(new_n755), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1107), .A2(new_n932), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1110), .B1(new_n1129), .B2(new_n1108), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1107), .A2(new_n932), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1120), .A2(new_n1121), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n469), .A2(new_n749), .A3(G330), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n941), .A2(new_n664), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1113), .A2(new_n1108), .A3(new_n1117), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1120), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1135), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1142), .A3(new_n711), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT54), .B(G143), .Z(new_n1144));
  AOI22_X1  g0944(.A1(new_n809), .A2(new_n1144), .B1(G137), .B2(new_n775), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT117), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n373), .B2(new_n789), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT118), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n787), .A2(G128), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n201), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n762), .A2(new_n1150), .B1(new_n1151), .B2(new_n769), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n255), .B1(new_n780), .B2(new_n854), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1022), .A2(G150), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1148), .A2(new_n1149), .A3(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n763), .A2(G294), .B1(G107), .B2(new_n775), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1158), .B(new_n852), .C1(new_n1037), .C2(new_n811), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n796), .A2(new_n212), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n808), .A2(new_n214), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n528), .B1(new_n258), .B2(new_n789), .C1(new_n780), .C2(new_n245), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT119), .Z(new_n1164));
  NAND2_X1  g0964(.A1(new_n1157), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n757), .B1(new_n1165), .B2(new_n821), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n928), .A2(new_n822), .A3(new_n930), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n866), .A2(new_n293), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1128), .A2(new_n1143), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT120), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1169), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n1143), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(G378));
  AOI21_X1  g0976(.A(KEYINPUT107), .B1(new_n919), .B2(new_n920), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n910), .B(KEYINPUT40), .C1(new_n918), .C2(new_n907), .ZN(new_n1178));
  OAI211_X1 g0978(.A(G330), .B(new_n908), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT56), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n302), .A2(new_n876), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n315), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT55), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n308), .A2(new_n311), .A3(new_n314), .A4(new_n1181), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT55), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(KEYINPUT56), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n931), .A2(new_n1193), .A3(new_n939), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n926), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n918), .A2(new_n935), .B1(new_n937), .B2(new_n687), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1179), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1193), .B1(new_n931), .B2(new_n939), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1197), .A3(new_n1195), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n922), .A2(new_n1200), .A3(G330), .A4(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n754), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1193), .A2(new_n822), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1150), .A2(new_n811), .B1(new_n776), .B2(new_n854), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n781), .A2(G128), .B1(G150), .B2(new_n790), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1027), .B2(new_n783), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(new_n1022), .C2(new_n1144), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT59), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G41), .B1(new_n770), .B2(new_n800), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G33), .B1(new_n761), .B2(G124), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n375), .A2(new_n377), .A3(G33), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n220), .B1(new_n1213), .B2(G41), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n781), .A2(G107), .B1(new_n441), .B2(new_n784), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n345), .B2(new_n789), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1216), .A2(G41), .A3(new_n401), .A4(new_n1060), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n770), .A2(G58), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n763), .A2(G283), .B1(G116), .B2(new_n787), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n775), .A2(G97), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT58), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1212), .A2(new_n1214), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n757), .B1(new_n1223), .B2(new_n821), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1204), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1151), .B2(new_n866), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1203), .A2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1202), .A2(new_n1199), .B1(new_n1142), .B2(new_n1136), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n711), .B1(new_n1228), .B2(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1142), .A2(new_n1136), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1230), .A2(KEYINPUT57), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1227), .B1(new_n1229), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n932), .A2(new_n822), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n762), .A2(new_n602), .B1(new_n245), .B2(new_n776), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1059), .B(new_n1235), .C1(G294), .C2(new_n787), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n809), .A2(G107), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n528), .B1(new_n796), .B2(new_n214), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n781), .B2(G283), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1018), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n811), .A2(new_n854), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n763), .A2(G128), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n401), .B1(new_n789), .B2(new_n220), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n780), .A2(new_n1027), .B1(new_n1024), .B2(new_n783), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(G159), .C2(new_n1022), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n775), .A2(new_n1144), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1242), .A2(new_n1245), .A3(new_n1218), .A4(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1240), .B1(new_n1241), .B2(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1248), .A2(new_n821), .B1(new_n345), .B2(new_n866), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1234), .A2(new_n756), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1133), .B2(new_n755), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1135), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n987), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1253), .B2(new_n1141), .ZN(G381));
  OR2_X1    g1054(.A1(new_n1203), .A2(new_n1226), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT57), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n712), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1228), .A2(KEYINPUT57), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1255), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1170), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1262), .A2(G384), .A3(G381), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(G390), .A2(G393), .A3(G396), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n1017), .A3(new_n1045), .A4(new_n1264), .ZN(G407));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G343), .C2(new_n1262), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  INV_X1    g1067(.A(G213), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(G343), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n1259), .A3(new_n711), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1174), .B1(new_n1173), .B2(new_n1143), .ZN(new_n1272));
  AND4_X1   g1072(.A1(new_n1174), .A2(new_n1128), .A3(new_n1143), .A4(new_n1169), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1271), .B(new_n1227), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1228), .A2(new_n987), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1227), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1261), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1269), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n712), .B1(new_n1252), .B2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1280), .B(new_n1137), .C1(new_n1279), .C2(new_n1252), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(G384), .A3(new_n1251), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1281), .B2(new_n1251), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT121), .B1(new_n1278), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1170), .B1(new_n1227), .B2(new_n1275), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1260), .B2(G378), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT121), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1285), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1269), .A4(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1267), .B1(new_n1286), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT122), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G390), .B1(new_n1017), .B2(new_n1045), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  XOR2_X1   g1096(.A(G393), .B(G396), .Z(new_n1297));
  NAND3_X1  g1097(.A1(new_n1017), .A2(new_n1045), .A3(G390), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1297), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1045), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1301), .B(new_n1105), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1295), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1284), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(G2897), .A3(new_n1269), .A4(new_n1282), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1269), .A2(G2897), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT123), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1305), .A2(new_n1307), .A3(KEYINPUT123), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1299), .B(new_n1303), .C1(new_n1312), .C2(new_n1278), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1273), .A2(new_n1272), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1277), .B1(new_n1315), .B2(G375), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1269), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1285), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1314), .B1(new_n1318), .B2(new_n1267), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1313), .A2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(KEYINPUT122), .B(new_n1267), .C1(new_n1286), .C2(new_n1291), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1294), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1318), .A2(new_n1289), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT62), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1316), .A2(KEYINPUT121), .A3(new_n1317), .A4(new_n1285), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT124), .B1(new_n1329), .B2(KEYINPUT61), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT124), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1331), .B(new_n1314), .C1(new_n1278), .C2(new_n1328), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1326), .A2(new_n1327), .A3(new_n1330), .A4(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1299), .A2(new_n1303), .A3(KEYINPUT125), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT125), .B1(new_n1299), .B2(new_n1303), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1333), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1322), .A2(new_n1338), .ZN(G405));
  OAI211_X1 g1139(.A(new_n1274), .B(KEYINPUT126), .C1(new_n1170), .C2(new_n1260), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1290), .A2(KEYINPUT127), .ZN(new_n1341));
  OR3_X1    g1141(.A1(new_n1260), .A2(KEYINPUT126), .A3(new_n1170), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1340), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1290), .A2(KEYINPUT127), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1335), .A2(new_n1336), .A3(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1344), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT125), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1297), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1348));
  NOR3_X1   g1148(.A1(new_n1295), .A2(new_n1302), .A3(new_n1300), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1347), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1346), .B1(new_n1350), .B2(new_n1334), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1343), .B1(new_n1345), .B2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1344), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1343), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1350), .A2(new_n1334), .A3(new_n1346), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1353), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1352), .A2(new_n1356), .ZN(G402));
endmodule


