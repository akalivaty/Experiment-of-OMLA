//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(new_n452));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n467), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n471), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G101), .ZN(new_n479));
  OR3_X1    g054(.A1(new_n466), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT71), .B1(new_n466), .B2(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n474), .A2(new_n478), .A3(new_n482), .ZN(G160));
  AND4_X1   g058(.A1(G2105), .A2(new_n467), .A3(new_n471), .A4(new_n469), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n470), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n472), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G136), .B2(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(new_n475), .A2(new_n471), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(new_n470), .A3(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT72), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(new_n475), .A4(new_n471), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n495), .A2(G2105), .ZN(new_n499));
  AND4_X1   g074(.A1(new_n467), .A2(new_n469), .A3(new_n499), .A4(new_n471), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n494), .B(new_n498), .C1(new_n500), .C2(new_n492), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n484), .B2(G126), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT75), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n515), .A2(new_n517), .B1(KEYINPUT5), .B2(new_n514), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(KEYINPUT74), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT6), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT76), .B(G88), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n514), .B1(new_n527), .B2(new_n529), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G50), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n523), .A2(new_n534), .A3(new_n536), .ZN(G166));
  NAND2_X1  g112(.A1(new_n532), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(G51), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n538), .A2(new_n539), .A3(new_n541), .A4(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  AOI22_X1  g119(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n526), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n535), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n531), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n526), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n535), .A2(G43), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n531), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT77), .Z(G176));
  XOR2_X1   g134(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n560));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n535), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n532), .A2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n524), .A2(G65), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n526), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  XNOR2_X1  g148(.A(G171), .B(new_n573), .ZN(G301));
  NAND3_X1  g149(.A1(new_n523), .A2(new_n534), .A3(new_n536), .ZN(G303));
  OAI21_X1  g150(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n524), .A2(G87), .A3(new_n530), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n535), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n524), .A2(G86), .A3(new_n530), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n535), .A2(G48), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n526), .ZN(G305));
  AOI22_X1  g158(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n526), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n535), .A2(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n531), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(new_n532), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT80), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n520), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n535), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  MUX2_X1   g174(.A(new_n599), .B(G301), .S(G868), .Z(G321));
  XNOR2_X1  g175(.A(G321), .B(KEYINPUT81), .ZN(G284));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n571), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n571), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(new_n599), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(new_n556), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n599), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n480), .A2(new_n481), .ZN(new_n614));
  INV_X1    g189(.A(new_n491), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n621));
  INV_X1    g196(.A(new_n484), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G135), .B2(new_n489), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT83), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT82), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT84), .Z(G401));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n659), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n659), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G229));
  XOR2_X1   g251(.A(KEYINPUT87), .B(G16), .Z(new_n677));
  MUX2_X1   g252(.A(G303), .B(G22), .S(new_n677), .Z(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G23), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n681), .A2(G16), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(G288), .B2(G16), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT33), .B(G1976), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT32), .B(G1981), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n683), .B2(new_n684), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n680), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  MUX2_X1   g270(.A(G290), .B(G24), .S(new_n677), .Z(new_n696));
  XOR2_X1   g271(.A(KEYINPUT88), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n489), .A2(G131), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT86), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G107), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n484), .B2(G119), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n700), .B1(new_n708), .B2(new_n699), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n698), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n694), .A2(new_n695), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT36), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT90), .B(KEYINPUT36), .Z(new_n718));
  NOR2_X1   g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(new_n608), .B(G19), .S(new_n677), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT91), .B(G1341), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT26), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G105), .B2(new_n614), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n489), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n484), .A2(G129), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G29), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n729), .B(new_n730), .C1(G29), .C2(G32), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT27), .B(G1996), .Z(new_n733));
  AND2_X1   g308(.A1(new_n699), .A2(G33), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n489), .A2(G139), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n615), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n736), .B(new_n739), .C1(new_n470), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2072), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n732), .A2(new_n733), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n722), .B(new_n744), .C1(new_n733), .C2(new_n732), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(G28), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n699), .B1(new_n747), .B2(G28), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G160), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n699), .B1(new_n752), .B2(G34), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(G34), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n753), .B2(KEYINPUT94), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n751), .A2(new_n699), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n750), .B(new_n759), .C1(G29), .C2(new_n625), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  INV_X1    g336(.A(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G168), .B2(new_n762), .ZN(new_n764));
  INV_X1    g339(.A(G1966), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n760), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n677), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G1956), .Z(new_n771));
  NOR3_X1   g346(.A1(new_n745), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n762), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n762), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  INV_X1    g354(.A(G2090), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n699), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n699), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT29), .Z(new_n783));
  OAI211_X1 g358(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n742), .A2(new_n743), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT95), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n699), .A2(G26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT28), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n484), .A2(G128), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n470), .A2(G116), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n489), .A2(KEYINPUT92), .A3(G140), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n794));
  INV_X1    g369(.A(G140), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n472), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n788), .B1(new_n797), .B2(new_n699), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n762), .A2(G4), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n605), .B2(new_n762), .ZN(new_n802));
  INV_X1    g377(.A(G1348), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n786), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n773), .A2(new_n784), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n783), .A2(KEYINPUT98), .A3(new_n780), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n808));
  INV_X1    g383(.A(new_n783), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G2090), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n699), .A2(G27), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G164), .B2(new_n699), .ZN(new_n812));
  INV_X1    g387(.A(G2078), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n806), .A2(new_n807), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n717), .A2(new_n719), .A3(new_n815), .ZN(G311));
  OR3_X1    g391(.A1(new_n717), .A2(new_n719), .A3(new_n815), .ZN(G150));
  AOI22_X1  g392(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(new_n526), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n535), .A2(G55), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n531), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n819), .B2(KEYINPUT99), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n608), .A2(KEYINPUT100), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n556), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n820), .A2(new_n824), .A3(new_n827), .A4(new_n556), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n605), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n836), .A2(new_n837), .A3(G860), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n825), .A2(G860), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n625), .B(new_n751), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G162), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n506), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT102), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n797), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n741), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n728), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n728), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n707), .B(new_n617), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n489), .A2(G142), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n484), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n470), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n854), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n851), .B2(new_n852), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n844), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n844), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT103), .B1(new_n853), .B2(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n853), .A2(KEYINPUT103), .A3(new_n861), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n842), .B(new_n864), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g445(.A1(G166), .A2(KEYINPUT105), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  NOR2_X1   g447(.A1(G303), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G290), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n589), .B1(new_n871), .B2(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G305), .B(G288), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(KEYINPUT107), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(KEYINPUT107), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n831), .B(new_n611), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n605), .A2(KEYINPUT104), .A3(G299), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT104), .B1(new_n599), .B2(new_n571), .ZN(new_n889));
  NAND3_X1  g464(.A1(G299), .A2(new_n593), .A3(new_n598), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n599), .A2(new_n571), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n887), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n886), .A2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(G868), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n825), .A2(new_n609), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(G295));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(G331));
  NOR2_X1   g479(.A1(G301), .A2(G286), .ZN(new_n905));
  NOR2_X1   g480(.A1(G168), .A2(G171), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n830), .B(new_n829), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G171), .B(KEYINPUT79), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n908), .B2(G168), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n831), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n891), .A2(new_n888), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n893), .A2(new_n896), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n879), .B(new_n913), .C1(new_n914), .C2(new_n911), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n842), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n907), .A2(new_n910), .B1(new_n888), .B2(new_n891), .ZN(new_n920));
  INV_X1    g495(.A(new_n911), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n897), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(new_n879), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n915), .A2(KEYINPUT108), .A3(new_n842), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n918), .A2(new_n919), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n912), .B1(new_n911), .B2(new_n895), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n890), .A2(new_n894), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n907), .A2(new_n910), .A3(KEYINPUT41), .A4(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n879), .A3(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n930), .B(new_n842), .C1(new_n922), .C2(new_n879), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n926), .B1(new_n931), .B2(KEYINPUT43), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n925), .A2(KEYINPUT109), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT109), .B1(new_n925), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n918), .A2(new_n923), .A3(new_n924), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n936), .B2(KEYINPUT43), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n933), .A2(new_n934), .B1(KEYINPUT44), .B2(new_n937), .ZN(G397));
  XNOR2_X1  g513(.A(new_n797), .B(G2067), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n728), .B(G1996), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n708), .A2(new_n710), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n711), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT102), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT102), .B1(new_n501), .B2(new_n505), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  XOR2_X1   g524(.A(KEYINPUT110), .B(G40), .Z(new_n950));
  NOR4_X1   g525(.A1(new_n474), .A2(new_n478), .A3(new_n482), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n943), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT127), .Z(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(G1986), .A3(G290), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT48), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n939), .A2(new_n940), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(new_n941), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n799), .B2(new_n797), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n954), .A2(new_n956), .B1(new_n952), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n952), .A2(G1996), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT46), .Z(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n952), .B1(new_n728), .B2(new_n939), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT126), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT47), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OR3_X1    g541(.A1(new_n963), .A2(KEYINPUT47), .A3(new_n965), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n510), .B2(new_n947), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n949), .A2(G1384), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n846), .A2(new_n847), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n951), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n679), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n501), .B2(new_n505), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n951), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT73), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT73), .B1(new_n501), .B2(new_n505), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n947), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n979), .B(new_n780), .C1(new_n982), .C2(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n970), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT55), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n969), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n508), .B2(new_n509), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n951), .B(new_n973), .C1(new_n989), .C2(KEYINPUT45), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n978), .B1(new_n989), .B2(new_n977), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n990), .A2(new_n679), .B1(new_n991), .B2(new_n780), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT115), .B(new_n986), .C1(new_n992), .C2(new_n970), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n976), .A2(new_n951), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1981), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n580), .A2(new_n581), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n524), .A2(G61), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G73), .A2(G543), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G651), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n998), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(G305), .B2(G1981), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1000), .A2(new_n1004), .A3(KEYINPUT112), .A4(new_n998), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n997), .B1(new_n1009), .B2(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1005), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(KEYINPUT49), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  OR2_X1    g593(.A1(G288), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n995), .A2(new_n1019), .A3(G8), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(KEYINPUT111), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n995), .A2(G8), .A3(new_n1019), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(KEYINPUT52), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT116), .B1(new_n1017), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n996), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1009), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT113), .B1(new_n1009), .B2(KEYINPUT49), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1025), .A2(new_n1021), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1022), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1027), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n506), .A2(new_n977), .A3(new_n947), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n951), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(KEYINPUT50), .B2(new_n982), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n780), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n975), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(G8), .A3(new_n987), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT110), .B(G40), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G160), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n977), .B2(new_n976), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n758), .B(new_n1048), .C1(new_n989), .C2(new_n977), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT117), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT45), .B(new_n947), .C1(new_n980), .C2(new_n981), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n506), .A2(new_n947), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1047), .B1(new_n1052), .B2(new_n949), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n765), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n758), .A4(new_n1048), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(G8), .A3(G168), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n994), .A2(new_n1039), .A3(new_n1045), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT63), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1044), .A2(G8), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n986), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(KEYINPUT63), .A3(new_n1045), .A4(new_n1061), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1047), .B1(new_n946), .B2(new_n972), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n982), .A2(new_n949), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n813), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1048), .B1(new_n989), .B2(new_n977), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1072), .A2(new_n1073), .B1(new_n777), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1073), .A2(G2078), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1051), .A2(new_n1053), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AND4_X1   g653(.A1(new_n1039), .A2(new_n994), .A3(new_n1045), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1058), .A2(new_n1055), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1057), .B1(new_n1042), .B2(new_n758), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G286), .A2(G8), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT51), .B1(new_n1083), .B2(KEYINPUT124), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  OAI211_X1 g662(.A(G8), .B(new_n1084), .C1(new_n1059), .C2(G286), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1059), .A2(G8), .A3(G286), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1079), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1033), .A2(new_n1094), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1095), .A2(new_n996), .B1(new_n1045), .B2(new_n1065), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT114), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1069), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1074), .A2(new_n777), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n948), .A2(new_n949), .ZN(new_n1102));
  AND3_X1   g677(.A1(G160), .A2(G40), .A3(new_n1076), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n973), .A3(new_n1103), .ZN(new_n1104));
  AND4_X1   g679(.A1(G301), .A2(new_n1100), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1099), .B1(new_n1105), .B2(new_n1078), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n970), .B(new_n986), .C1(new_n1043), .C2(new_n975), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n988), .B2(new_n993), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1108), .A3(new_n1039), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1075), .A2(G301), .A3(new_n1077), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT54), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1100), .A2(new_n1104), .A3(new_n1101), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G171), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1109), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n571), .B(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n991), .A2(G1956), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1070), .A2(new_n1071), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1122), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n995), .A2(G2067), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1074), .B2(new_n803), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n599), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1126), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1042), .A2(G1348), .B1(G2067), .B2(new_n995), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI211_X1 g710(.A(KEYINPUT122), .B(new_n599), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n1137));
  AOI21_X1  g712(.A(G1348), .B1(new_n1056), .B2(new_n1048), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1133), .B1(new_n1138), .B2(new_n1128), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1139), .B2(new_n605), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n605), .B1(new_n1129), .B2(KEYINPUT60), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT122), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1137), .A3(new_n605), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1134), .A3(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n995), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n990), .B2(G1996), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n556), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT120), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(new_n556), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1148), .A2(new_n1154), .A3(new_n556), .A4(new_n1149), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1141), .A2(new_n1145), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1127), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1127), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1120), .B(new_n1131), .C1(new_n1157), .C2(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1119), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1131), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT123), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1098), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n589), .B(G1986), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n952), .B1(new_n943), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n968), .B1(new_n1166), .B2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g744(.A1(G227), .A2(new_n463), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n644), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G229), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n869), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1174), .A2(new_n937), .ZN(G308));
  OR2_X1    g749(.A1(new_n1174), .A2(new_n937), .ZN(G225));
endmodule


