//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1370, new_n1371;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT66), .B(G77), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n211), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n211), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n228), .A2(G50), .A3(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n209), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AND4_X1   g0034(.A1(new_n222), .A2(new_n226), .A3(new_n227), .A4(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n259), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n257), .B1(new_n258), .B2(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n265), .B(new_n268), .C1(new_n212), .C2(new_n257), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(new_n267), .A3(G274), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(G226), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G200), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT10), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n232), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n209), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n289), .A2(new_n291), .B1(G150), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n286), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n208), .A2(G20), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(G50), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G50), .B2(new_n296), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n283), .A2(new_n284), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n281), .A3(new_n303), .A4(new_n282), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n309), .B2(new_n279), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G179), .B2(new_n279), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(new_n291), .B1(new_n212), .B2(G20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n289), .A2(new_n292), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n287), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n298), .A2(G77), .A3(new_n299), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n212), .B2(new_n296), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n273), .B1(new_n214), .B2(new_n276), .ZN(new_n320));
  INV_X1    g0120(.A(G232), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n255), .B2(new_n256), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n259), .B1(new_n255), .B2(new_n256), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G238), .ZN(new_n328));
  AND2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G107), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n320), .B1(new_n333), .B2(new_n268), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n319), .B(new_n336), .C1(G169), .C2(new_n334), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(G190), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n316), .A2(new_n318), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n334), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n308), .A2(new_n311), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT70), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n308), .A2(KEYINPUT70), .A3(new_n311), .A4(new_n342), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n288), .B1(new_n208), .B2(G20), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n298), .B1(new_n297), .B2(new_n288), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n255), .A2(new_n209), .A3(new_n256), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n331), .B2(new_n209), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(G58), .A2(G68), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n355), .B2(new_n201), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n292), .A2(G159), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n287), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  INV_X1    g0161(.A(G68), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n350), .A2(new_n351), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n356), .A2(new_n357), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n349), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n261), .B(new_n262), .C1(new_n329), .C2(new_n330), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n258), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G226), .A2(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G87), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n331), .A2(new_n371), .B1(new_n254), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n268), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n267), .A2(G232), .A3(new_n275), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n273), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(G190), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n377), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G200), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n368), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n273), .A2(new_n375), .A3(new_n335), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n374), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n371), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n257), .A2(new_n388), .B1(G33), .B2(G87), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n257), .A2(new_n325), .A3(G223), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n267), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT75), .B1(new_n391), .B2(new_n385), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n387), .A2(new_n392), .B1(new_n379), .B2(new_n309), .ZN(new_n393));
  INV_X1    g0193(.A(new_n366), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT16), .B1(new_n354), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n286), .B1(new_n365), .B2(new_n358), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n348), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(KEYINPUT18), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT18), .B1(new_n393), .B2(new_n397), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n383), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n345), .A2(new_n346), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G226), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT71), .B1(new_n369), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n322), .B2(G1698), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT71), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n257), .A2(new_n325), .A3(new_n409), .A4(G226), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n268), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n276), .A2(KEYINPUT73), .ZN(new_n414));
  INV_X1    g0214(.A(G238), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n276), .B2(KEYINPUT73), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT72), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n273), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n272), .A2(new_n267), .A3(KEYINPUT72), .A4(G274), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n414), .A2(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n412), .A2(new_n413), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n413), .B1(new_n412), .B2(new_n420), .ZN(new_n422));
  OAI21_X1  g0222(.A(G200), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(G232), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n406), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n257), .A2(new_n325), .A3(G226), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(KEYINPUT71), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n267), .B1(new_n427), .B2(new_n410), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n414), .A2(new_n416), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(new_n419), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT13), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n412), .A2(new_n413), .A3(new_n420), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(G190), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n362), .ZN(new_n435));
  INV_X1    g0235(.A(G77), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n290), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(new_n286), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n438), .A2(KEYINPUT11), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n297), .A2(new_n362), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(KEYINPUT11), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n298), .A2(G68), .A3(new_n299), .ZN(new_n443));
  AND4_X1   g0243(.A1(new_n439), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n423), .A2(new_n434), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(G169), .C1(new_n421), .C2(new_n422), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n432), .A2(G179), .A3(new_n433), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT74), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n309), .B1(new_n432), .B2(new_n433), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n446), .ZN(new_n452));
  OAI21_X1  g0252(.A(G169), .B1(new_n421), .B2(new_n422), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n449), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n445), .B1(new_n455), .B2(new_n444), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n403), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n327), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n214), .B1(new_n255), .B2(new_n256), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n325), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT4), .ZN(new_n462));
  OAI21_X1  g0262(.A(G244), .B1(new_n329), .B2(new_n330), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n263), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n268), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n208), .B(G45), .C1(new_n270), .C2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  OAI211_X1 g0269(.A(G257), .B(new_n267), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n267), .A2(G274), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT76), .B1(new_n468), .B2(G41), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT76), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n270), .A3(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n271), .A2(G1), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n470), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n309), .ZN(new_n481));
  XNOR2_X1  g0281(.A(G97), .B(G107), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n204), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n482), .A2(new_n483), .B1(new_n205), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n292), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n485), .A2(new_n209), .B1(new_n436), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n205), .B1(new_n363), .B2(new_n364), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n286), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n296), .A2(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n208), .A2(G33), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n296), .A2(new_n491), .A3(new_n232), .A4(new_n285), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n478), .B1(new_n465), .B2(new_n268), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n335), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n481), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n494), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n482), .A2(new_n483), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n484), .A2(new_n205), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n503));
  OAI21_X1  g0303(.A(G107), .B1(new_n352), .B2(new_n353), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n499), .B1(new_n505), .B2(new_n286), .ZN(new_n506));
  AOI21_X1  g0306(.A(G200), .B1(new_n466), .B2(new_n479), .ZN(new_n507));
  AOI211_X1 g0307(.A(G190), .B(new_n478), .C1(new_n465), .C2(new_n268), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT77), .B1(new_n369), .B2(new_n415), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n460), .B2(G1698), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT77), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n257), .A2(new_n325), .A3(new_n514), .A4(G238), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n510), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n268), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n476), .A2(G250), .ZN(new_n518));
  INV_X1    g0318(.A(G274), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n476), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n267), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(new_n335), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n209), .B1(new_n406), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G87), .B2(new_n206), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n209), .B(G68), .C1(new_n329), .C2(new_n330), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n523), .B1(new_n290), .B2(new_n204), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(new_n286), .B1(new_n297), .B2(new_n312), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n493), .A2(new_n313), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n521), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n516), .B2(new_n268), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n522), .B(new_n531), .C1(G169), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n517), .A2(G190), .A3(new_n521), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n286), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n312), .A2(new_n297), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n493), .A2(G87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n535), .B(new_n540), .C1(new_n340), .C2(new_n533), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n498), .A2(new_n509), .A3(new_n534), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n257), .A2(new_n209), .A3(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT22), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n257), .A2(new_n545), .A3(new_n209), .A4(G87), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT79), .B1(new_n511), .B2(G20), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT79), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(new_n209), .A3(G33), .A4(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n205), .A2(G20), .ZN(new_n554));
  AND2_X1   g0354(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n209), .A2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n551), .A3(new_n552), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n550), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n550), .A2(new_n556), .A3(KEYINPUT81), .A4(new_n558), .ZN(new_n562));
  AOI221_X4 g0362(.A(KEYINPUT24), .B1(new_n544), .B2(new_n546), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n544), .A2(new_n546), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n286), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n208), .A2(G13), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT82), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT25), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n554), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  OAI211_X1 g0373(.A(KEYINPUT82), .B(KEYINPUT25), .C1(new_n554), .C2(new_n569), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n205), .C2(new_n492), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n477), .A2(new_n471), .ZN(new_n577));
  OAI211_X1 g0377(.A(G264), .B(new_n267), .C1(new_n467), .C2(new_n469), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n261), .A2(G250), .A3(new_n262), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G257), .A2(G1698), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n257), .B1(G33), .B2(G294), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n577), .B(new_n578), .C1(new_n582), .C2(new_n267), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n340), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(G190), .B2(new_n583), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n568), .A2(new_n576), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n587));
  NAND2_X1  g0387(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n557), .B2(new_n588), .ZN(new_n589));
  NOR4_X1   g0389(.A1(new_n209), .A2(KEYINPUT80), .A3(KEYINPUT23), .A4(G107), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT81), .B1(new_n591), .B2(new_n550), .ZN(new_n592));
  INV_X1    g0392(.A(new_n562), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n566), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n565), .A2(new_n564), .A3(new_n566), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n287), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n582), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n268), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(G179), .A3(new_n577), .A4(new_n578), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n583), .A2(KEYINPUT83), .A3(G169), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT83), .B1(new_n583), .B2(G169), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n597), .A2(new_n575), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G264), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT78), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT78), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n257), .A2(new_n607), .A3(G264), .A4(G1698), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n257), .A2(new_n325), .A3(G257), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n331), .A2(G303), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n606), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n268), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n267), .B1(new_n467), .B2(new_n469), .ZN(new_n613));
  INV_X1    g0413(.A(G270), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(new_n477), .B2(new_n471), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n492), .A2(G116), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n296), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n285), .A2(new_n232), .B1(G20), .B2(new_n619), .ZN(new_n622));
  AOI21_X1  g0422(.A(G20), .B1(G33), .B2(G283), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(G33), .B2(new_n204), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT20), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n622), .A2(new_n624), .A3(KEYINPUT20), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n617), .A2(KEYINPUT21), .A3(G169), .A4(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(G169), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n615), .B1(new_n611), .B2(new_n268), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n627), .A3(G179), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n628), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G190), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n617), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n627), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n631), .B2(new_n340), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n542), .A2(new_n586), .A3(new_n604), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n458), .A2(new_n641), .ZN(G372));
  AND3_X1   g0442(.A1(new_n536), .A2(new_n537), .A3(new_n530), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n517), .A2(new_n521), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n309), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n539), .B1(new_n533), .B2(G190), .ZN(new_n646));
  OAI211_X1 g0446(.A(G244), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n511), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n257), .A2(new_n325), .A3(G238), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(KEYINPUT77), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n267), .B1(new_n650), .B2(new_n515), .ZN(new_n651));
  OAI21_X1  g0451(.A(G200), .B1(new_n651), .B2(new_n532), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n645), .A2(new_n522), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n498), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT26), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT26), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n466), .A2(new_n635), .A3(new_n479), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(G200), .B2(new_n496), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n335), .A2(new_n496), .B1(new_n489), .B2(new_n494), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n659), .A2(new_n506), .B1(new_n660), .B2(new_n481), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n653), .A3(new_n586), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n568), .A2(new_n576), .ZN(new_n663));
  INV_X1    g0463(.A(new_n603), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n600), .A3(new_n601), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n634), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n534), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n457), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n311), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT18), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n309), .B1(new_n391), .B2(new_n376), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n384), .B1(new_n374), .B2(new_n386), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n391), .A2(KEYINPUT75), .A3(new_n385), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n675), .A2(new_n368), .A3(KEYINPUT84), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT84), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n393), .B2(new_n397), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n671), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT84), .B1(new_n675), .B2(new_n368), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n393), .A2(new_n677), .A3(new_n397), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(KEYINPUT18), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n447), .A2(new_n448), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n451), .A2(new_n450), .A3(new_n446), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT74), .B1(new_n453), .B2(KEYINPUT14), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n444), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n334), .A2(G169), .B1(new_n318), .B2(new_n316), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n334), .A2(new_n335), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n687), .A2(new_n688), .B1(new_n445), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n683), .B1(new_n692), .B2(new_n383), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n670), .B1(new_n693), .B2(new_n308), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n669), .A2(new_n694), .ZN(G369));
  INV_X1    g0495(.A(new_n586), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT85), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n569), .B2(G20), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT85), .A4(G13), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(G213), .A3(G343), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n568), .B2(new_n576), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n604), .B1(new_n696), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n703), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n604), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n634), .A2(new_n703), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n708), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n637), .A2(new_n703), .ZN(new_n712));
  MUX2_X1   g0512(.A(new_n640), .B(new_n634), .S(new_n712), .Z(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n706), .A2(new_n708), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(G399));
  NAND2_X1  g0517(.A1(new_n223), .A2(new_n270), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n230), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(new_n578), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n598), .B2(new_n268), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(new_n496), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n631), .A2(G179), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n727), .A3(KEYINPUT30), .A4(new_n533), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n533), .A3(new_n496), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n496), .A2(G179), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n583), .A3(new_n644), .A4(new_n617), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n707), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT86), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n641), .B2(new_n707), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n640), .A2(new_n604), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n662), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(KEYINPUT86), .A4(new_n703), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n739), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G330), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT87), .B(KEYINPUT29), .Z(new_n749));
  NAND3_X1  g0549(.A1(new_n668), .A2(new_n703), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n668), .A2(new_n703), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT87), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT29), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n748), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n722), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n713), .A2(G330), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT88), .ZN(new_n758));
  INV_X1    g0558(.A(new_n718), .ZN(new_n759));
  INV_X1    g0559(.A(G13), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n208), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n758), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n718), .A2(KEYINPUT88), .A3(new_n762), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n757), .B(new_n714), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n223), .A2(new_n257), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n223), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n223), .A2(new_n331), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n231), .B2(new_n271), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n251), .A2(G45), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n232), .B1(G20), .B2(new_n309), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n768), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n209), .A2(new_n635), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(new_n340), .A3(G179), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n257), .B1(new_n785), .B2(G303), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT93), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n209), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n789), .A2(G179), .A3(new_n340), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT92), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n335), .A2(new_n340), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT91), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n789), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n791), .A2(G283), .B1(G329), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(G20), .B1(new_n793), .B2(new_n635), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G294), .ZN(new_n797));
  NAND3_X1  g0597(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n635), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G326), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n335), .A2(G200), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n783), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n788), .A2(new_n803), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n798), .A2(G190), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT33), .B(G317), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n802), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n787), .A2(new_n795), .A3(new_n797), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n791), .A2(G107), .ZN(new_n813));
  INV_X1    g0613(.A(new_n809), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n362), .ZN(new_n815));
  INV_X1    g0615(.A(new_n785), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n372), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n813), .A2(new_n331), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n794), .A2(G159), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT32), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n796), .A2(G97), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G50), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n213), .A2(new_n806), .B1(new_n800), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n804), .B(KEYINPUT89), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n824), .B1(new_n826), .B2(G58), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT90), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n812), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n782), .B1(new_n829), .B2(new_n779), .ZN(new_n830));
  INV_X1    g0630(.A(new_n778), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n713), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT94), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n766), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  NAND2_X1  g0635(.A1(new_n791), .A2(G68), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n331), .B1(new_n785), .B2(G50), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  INV_X1    g0638(.A(new_n794), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G58), .B2(new_n796), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT96), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(new_n806), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n845), .A2(G159), .B1(G137), .B2(new_n799), .ZN(new_n846));
  INV_X1    g0646(.A(G150), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n814), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G143), .B2(new_n826), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT34), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n843), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n791), .A2(G87), .B1(G311), .B2(new_n794), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT95), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n816), .A2(new_n205), .B1(new_n806), .B2(new_n619), .ZN(new_n854));
  INV_X1    g0654(.A(new_n804), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n257), .B(new_n854), .C1(G294), .C2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n809), .A2(G283), .B1(new_n799), .B2(G303), .ZN(new_n857));
  AND4_X1   g0657(.A1(new_n821), .A2(new_n853), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n779), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n779), .A2(new_n776), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n859), .B(new_n768), .C1(G77), .C2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n337), .B(new_n341), .C1(new_n339), .C2(new_n703), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT97), .B1(new_n691), .B2(new_n707), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT97), .ZN(new_n865));
  NOR4_X1   g0665(.A1(new_n689), .A2(new_n690), .A3(new_n703), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT98), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT98), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n863), .B(new_n869), .C1(new_n864), .C2(new_n866), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n862), .B1(new_n776), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n751), .A2(new_n872), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n871), .B(new_n703), .C1(new_n657), .C2(new_n667), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n748), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n764), .B2(new_n765), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n748), .A3(new_n875), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  NOR2_X1   g0680(.A1(new_n761), .A2(new_n208), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n457), .A2(new_n754), .A3(new_n750), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n694), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT103), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n397), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n383), .B2(new_n401), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n393), .A2(new_n397), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n381), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n381), .A2(new_n891), .A3(new_n894), .A4(new_n888), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n890), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n381), .B(KEYINPUT17), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n683), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n889), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n380), .A2(new_n378), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n680), .A2(new_n681), .B1(new_n368), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT101), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n889), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n680), .A2(new_n681), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n381), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT101), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n894), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n895), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n902), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n899), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n399), .A2(new_n400), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n888), .B1(new_n915), .B2(new_n900), .ZN(new_n916));
  INV_X1    g0716(.A(new_n896), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n898), .B1(new_n918), .B2(new_n897), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n885), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n897), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT39), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n888), .B1(new_n683), .B2(new_n900), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n905), .B(new_n381), .C1(new_n676), .C2(new_n678), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n888), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n905), .B1(new_n907), .B2(new_n381), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n927), .B2(new_n895), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(KEYINPUT38), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n922), .B(KEYINPUT102), .C1(new_n929), .C2(new_n899), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n920), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n687), .A2(new_n688), .A3(new_n703), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n691), .A2(new_n703), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n875), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n684), .B(new_n445), .C1(new_n685), .C2(new_n686), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n444), .A2(new_n703), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT100), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n938), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n445), .B(new_n942), .C1(new_n455), .C2(new_n444), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n937), .A2(KEYINPUT100), .A3(new_n938), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n936), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n921), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n946), .A2(new_n947), .B1(new_n683), .B2(new_n887), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n934), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n884), .B(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n737), .A2(new_n738), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n742), .A2(new_n662), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT86), .B1(new_n953), .B2(new_n703), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n742), .A2(new_n662), .A3(new_n740), .A4(new_n707), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n945), .A2(new_n956), .A3(new_n921), .A4(new_n871), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT40), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n897), .B1(new_n928), .B2(KEYINPUT38), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n741), .A2(new_n745), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n872), .B1(new_n961), .B2(new_n952), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n960), .A2(new_n962), .A3(KEYINPUT40), .A4(new_n945), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n458), .A2(new_n746), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n747), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n965), .B2(new_n964), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n881), .B1(new_n951), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n951), .B2(new_n967), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(G116), .A3(new_n233), .A4(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n230), .A2(new_n213), .A3(new_n355), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n362), .A2(G50), .ZN(new_n976));
  OAI211_X1 g0776(.A(G1), .B(new_n760), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n969), .A2(new_n974), .A3(new_n977), .ZN(G367));
  OAI21_X1  g0778(.A(new_n661), .B1(new_n506), .B2(new_n703), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n498), .B2(new_n703), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n710), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT42), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n979), .A2(new_n604), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n707), .B1(new_n983), .B2(new_n498), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n981), .B2(KEYINPUT42), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n653), .B1(new_n540), .B2(new_n703), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n645), .A2(new_n522), .A3(new_n539), .A4(new_n707), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n982), .A2(new_n985), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n716), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n980), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n991), .B(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n718), .B(KEYINPUT41), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n711), .A2(new_n980), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT104), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT104), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n711), .A2(new_n998), .A3(new_n980), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n711), .A2(new_n980), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n997), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n992), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n715), .B(new_n709), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n755), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1002), .A2(new_n1004), .A3(new_n716), .A4(new_n1005), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1007), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n995), .B1(new_n1016), .B2(new_n755), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n994), .B1(new_n1017), .B2(new_n763), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n243), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n780), .B1(new_n223), .B2(new_n312), .C1(new_n1019), .C2(new_n772), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n768), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n816), .A2(new_n619), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(KEYINPUT46), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G294), .B2(new_n809), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1022), .A2(KEYINPUT46), .B1(new_n799), .B2(G311), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n796), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1025), .C1(new_n205), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(G283), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n790), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n331), .B1(new_n1028), .B2(new_n806), .C1(new_n1029), .C2(new_n204), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G317), .B2(new_n794), .ZN(new_n1031));
  INV_X1    g0831(.A(G303), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n825), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n794), .A2(G137), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n331), .B1(new_n785), .B2(G58), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n790), .A2(new_n212), .B1(new_n855), .B2(G150), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n799), .A2(G143), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n796), .A2(G68), .ZN(new_n1039));
  INV_X1    g0839(.A(G159), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n814), .A2(new_n1040), .B1(new_n806), .B2(new_n823), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT106), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT106), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1027), .A2(new_n1033), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT47), .Z(new_n1046));
  INV_X1    g0846(.A(new_n779), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1021), .B1(new_n831), .B2(new_n988), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1018), .A2(new_n1048), .ZN(G387));
  INV_X1    g0849(.A(new_n1014), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n718), .B(KEYINPUT113), .Z(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1012), .A2(new_n762), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n778), .B1(new_n706), .B2(new_n708), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n769), .A2(new_n719), .B1(G107), .B2(new_n223), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n719), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT107), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n271), .B1(new_n362), .B2(new_n436), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n288), .A2(G50), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n772), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT109), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1064), .A2(new_n1065), .B1(G45), .B2(new_n240), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1056), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n768), .B1(new_n1068), .B2(new_n781), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n791), .A2(G97), .B1(G150), .B2(new_n794), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n796), .A2(new_n313), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n816), .A2(new_n213), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n804), .A2(new_n823), .B1(new_n806), .B2(new_n362), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n331), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n289), .A2(new_n809), .B1(G159), .B2(new_n799), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n826), .A2(G317), .B1(G303), .B2(new_n845), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(KEYINPUT111), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(KEYINPUT111), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n809), .A2(G311), .B1(new_n799), .B2(G322), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT112), .Z(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT48), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n796), .A2(G283), .B1(G294), .B2(new_n785), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT110), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1083), .B2(new_n1082), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1088), .A3(KEYINPUT49), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n257), .B1(new_n790), .B2(G116), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n801), .C2(new_n839), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT49), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1076), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1069), .B1(new_n1093), .B2(new_n779), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1054), .B1(new_n1055), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1053), .A2(new_n1095), .ZN(G393));
  NAND3_X1  g0896(.A1(new_n1007), .A2(new_n763), .A3(new_n1015), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n248), .A2(new_n223), .A3(new_n331), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n780), .B1(new_n204), .B2(new_n223), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n768), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n257), .B1(new_n845), .B2(G294), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n1032), .B2(new_n814), .C1(new_n816), .C2(new_n1028), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1102), .B(new_n813), .C1(G322), .C2(new_n794), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n855), .A2(G311), .B1(G317), .B2(new_n799), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(new_n619), .C2(new_n1026), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1106), .A2(KEYINPUT114), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(KEYINPUT114), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n257), .B1(new_n806), .B2(new_n288), .C1(new_n816), .C2(new_n362), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G50), .B2(new_n809), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n800), .A2(new_n847), .B1(new_n804), .B2(new_n1040), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT51), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n796), .A2(G77), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n791), .A2(G87), .B1(G143), .B2(new_n794), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1107), .A2(new_n1108), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1100), .B1(new_n1116), .B2(new_n779), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n831), .B2(new_n980), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1016), .A2(new_n1052), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1014), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1097), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(G390));
  NAND2_X1  g0921(.A1(new_n946), .A2(new_n932), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n920), .A2(new_n1122), .A3(new_n930), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n945), .A2(new_n956), .A3(G330), .A4(new_n871), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n960), .A2(new_n932), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n943), .A2(new_n944), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT100), .B1(new_n937), .B2(new_n938), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT115), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT115), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n941), .A2(new_n1130), .A3(new_n943), .A4(new_n944), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1126), .B1(new_n936), .B2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1123), .A2(new_n1125), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1133), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n920), .A2(new_n1122), .A3(new_n930), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1124), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n920), .A2(new_n930), .A3(new_n776), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n768), .B1(new_n289), .B2(new_n861), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n804), .A2(new_n619), .B1(new_n806), .B2(new_n204), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n814), .A2(new_n205), .B1(new_n800), .B2(new_n1028), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n817), .A2(new_n257), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n794), .A2(G294), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1143), .A2(new_n836), .A3(new_n1113), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n809), .A2(G137), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n816), .A2(new_n847), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT53), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G128), .B2(new_n799), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n804), .A2(new_n838), .B1(new_n806), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(new_n1153), .C1(new_n1040), .C2(new_n1026), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n794), .A2(G125), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n257), .C1(new_n823), .C2(new_n1029), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT117), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1145), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1140), .B1(new_n1158), .B2(new_n779), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1138), .A2(new_n763), .B1(new_n1139), .B2(new_n1159), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n746), .A2(new_n747), .A3(new_n872), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT116), .B1(new_n1132), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n956), .A2(G330), .A3(new_n871), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT116), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n936), .B1(new_n1161), .B2(new_n945), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n945), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1124), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n936), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n457), .A2(new_n748), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n882), .A2(new_n694), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1125), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1174), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1135), .A2(new_n1136), .A3(new_n1124), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1177), .A2(new_n1052), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT118), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1160), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n1160), .B2(new_n1182), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(G378));
  NAND3_X1  g0987(.A1(new_n959), .A2(new_n963), .A3(G330), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n308), .A2(new_n311), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n302), .A2(new_n886), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1188), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1193), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1195), .A2(new_n959), .A3(new_n963), .A4(G330), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n950), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT120), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n948), .B1(new_n931), .B2(new_n933), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1200), .A2(new_n1194), .A3(KEYINPUT120), .A4(new_n1196), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n763), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n331), .A2(new_n270), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n823), .C1(G33), .C2(G41), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n804), .A2(new_n205), .B1(new_n806), .B2(new_n312), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(new_n1205), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n839), .B2(new_n1028), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1072), .B1(G58), .B2(new_n790), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n204), .B2(new_n814), .C1(new_n619), .C2(new_n800), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(G68), .C2(new_n796), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1206), .B1(new_n1212), .B2(KEYINPUT58), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT119), .Z(new_n1214));
  NAND2_X1  g1014(.A1(new_n855), .A2(G128), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n816), .B2(new_n1151), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G137), .B2(new_n845), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n809), .A2(G132), .B1(new_n799), .B2(G125), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n847), .C2(new_n1026), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n790), .C2(G159), .ZN(new_n1221));
  INV_X1    g1021(.A(G124), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1222), .B2(new_n839), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1219), .B2(KEYINPUT59), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1212), .A2(KEYINPUT58), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1047), .B1(new_n1214), .B2(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n767), .B(new_n1226), .C1(new_n823), .C2(new_n860), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1195), .B2(new_n777), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1204), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1181), .A2(new_n1175), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT121), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1198), .A2(new_n1235), .A3(new_n1201), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1200), .A2(new_n1194), .A3(KEYINPUT121), .A4(new_n1196), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1231), .A2(new_n1236), .A3(KEYINPUT57), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1052), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1230), .B1(new_n1234), .B2(new_n1239), .ZN(G375));
  NAND3_X1  g1040(.A1(new_n1129), .A2(new_n776), .A3(new_n1131), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n768), .B1(G68), .B2(new_n861), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n785), .A2(G97), .B1(G107), .B2(new_n845), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n257), .B1(new_n855), .B2(G283), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n809), .A2(G116), .B1(new_n799), .B2(G294), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n791), .A2(G77), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n794), .A2(G303), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1071), .A4(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n826), .A2(G137), .B1(G128), .B2(new_n794), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n331), .B1(new_n790), .B2(G58), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n785), .A2(G159), .B1(G150), .B2(new_n845), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1151), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1253), .A2(new_n809), .B1(G132), .B2(new_n799), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1026), .A2(new_n823), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1249), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1257), .A2(KEYINPUT122), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1047), .B1(new_n1257), .B2(KEYINPUT122), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1242), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1241), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n936), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1169), .B2(new_n1124), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1124), .A2(new_n1262), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1132), .A2(new_n1161), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n1164), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1263), .B1(new_n1266), .B2(new_n1162), .ZN(new_n1267));
  OAI211_X1 g1067(.A(KEYINPUT123), .B(new_n1261), .C1(new_n1267), .C2(new_n762), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT123), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n762), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1261), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n995), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1167), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1176), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT124), .ZN(G381));
  INV_X1    g1078(.A(G390), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1053), .A2(new_n834), .A3(new_n1095), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n879), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1160), .A2(new_n1182), .ZN(new_n1283));
  NOR4_X1   g1083(.A1(new_n1282), .A2(G381), .A3(G387), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1052), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1233), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1229), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1284), .A2(new_n1290), .ZN(G407));
  INV_X1    g1091(.A(new_n1283), .ZN(new_n1292));
  INV_X1    g1092(.A(G343), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(G213), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1290), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G407), .A2(G213), .A3(new_n1296), .ZN(G409));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1018), .A2(new_n1048), .A3(G390), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G390), .B1(new_n1018), .B2(new_n1048), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n834), .B1(new_n1053), .B2(new_n1095), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n1300), .A2(new_n1301), .B1(new_n1281), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1301), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1281), .A2(new_n1302), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1299), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1275), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1167), .A2(new_n1171), .A3(new_n1174), .A4(KEYINPUT60), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1310), .A2(new_n1176), .A3(new_n1052), .A4(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1273), .A2(G384), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G384), .B1(new_n1273), .B2(new_n1312), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1289), .A2(new_n1052), .A3(new_n1238), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1283), .A2(KEYINPUT118), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n1184), .A4(new_n1230), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1231), .A2(new_n1202), .A3(new_n1274), .A4(new_n1203), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1236), .A2(new_n763), .A3(new_n1237), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1228), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1292), .ZN(new_n1323));
  AOI211_X1 g1123(.A(new_n1295), .B(new_n1316), .C1(new_n1319), .C2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1308), .B1(new_n1324), .B2(KEYINPUT63), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1273), .A2(new_n1312), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n879), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1273), .A2(G384), .A3(new_n1312), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(KEYINPUT125), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1295), .A2(G2897), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1327), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1332), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1315), .A2(KEYINPUT125), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1321), .A2(new_n1228), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1283), .B1(new_n1337), .B2(new_n1320), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1338), .B1(new_n1290), .B2(G378), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1336), .B1(new_n1339), .B2(new_n1295), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1318), .A2(new_n1184), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1323), .B1(G375), .B2(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1342), .A2(KEYINPUT63), .A3(new_n1294), .A4(new_n1315), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT61), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1340), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1298), .B1(new_n1325), .B2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1342), .A2(new_n1294), .A3(new_n1315), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT63), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1307), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1342), .A2(new_n1294), .ZN(new_n1350));
  AOI21_X1  g1150(.A(KEYINPUT61), .B1(new_n1350), .B2(new_n1336), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1349), .A2(new_n1351), .A3(KEYINPUT126), .A4(new_n1343), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1346), .A2(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1295), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1354));
  NOR4_X1   g1154(.A1(new_n1313), .A2(new_n1314), .A3(new_n1326), .A4(new_n1332), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1334), .B1(new_n1315), .B2(KEYINPUT125), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1355), .B1(new_n1356), .B2(new_n1327), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1344), .B1(new_n1354), .B2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1347), .A2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1354), .A2(KEYINPUT62), .A3(new_n1315), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1358), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT127), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1307), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1361), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT62), .B1(new_n1354), .B2(new_n1315), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1363), .B(new_n1351), .C1(new_n1365), .C2(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1367), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1353), .B1(new_n1364), .B2(new_n1368), .ZN(G405));
  OAI21_X1  g1169(.A(new_n1319), .B1(new_n1283), .B2(new_n1290), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1370), .B(new_n1315), .ZN(new_n1371));
  XNOR2_X1  g1171(.A(new_n1371), .B(new_n1307), .ZN(G402));
endmodule


