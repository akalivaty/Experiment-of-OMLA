//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT65), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G113), .A3(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n469), .A2(new_n471), .A3(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(G101), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n469), .A2(new_n471), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n462), .B2(G114), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n496), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n489), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n507), .B(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(G50), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n515), .B(new_n517), .C1(new_n511), .C2(new_n512), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n510), .A2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n511), .A2(new_n512), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(new_n505), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n505), .A2(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n504), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(G52), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n518), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n504), .ZN(new_n542));
  OAI211_X1 g117(.A(G43), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n518), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n515), .A2(new_n517), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(KEYINPUT68), .A3(G651), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n542), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n548), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n518), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(G651), .B1(new_n563), .B2(G91), .ZN(new_n564));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(G299));
  AOI22_X1  g142(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n536), .B1(new_n537), .B2(new_n518), .C1(new_n568), .C2(new_n504), .ZN(G301));
  OR2_X1    g144(.A1(new_n510), .A2(new_n520), .ZN(G303));
  NAND2_X1  g145(.A1(new_n563), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n527), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n548), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n563), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n527), .A2(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n563), .A2(G85), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n527), .A2(G47), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n504), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n584), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n518), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n592));
  XNOR2_X1  g167(.A(KEYINPUT69), .B(G66), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n505), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g169(.A1(G79), .A2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n505), .A2(new_n593), .B1(G79), .B2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT70), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(G651), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n527), .A2(G54), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n591), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND4_X1  g185(.A1(new_n591), .A2(new_n599), .A3(new_n609), .A4(new_n600), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n553), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT71), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g190(.A1(new_n468), .A2(G2105), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n493), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n479), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT72), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n621), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2430), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n632), .A2(G2435), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n633), .B2(new_n634), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT14), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n640), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n641), .B2(new_n644), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n631), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n649), .A2(new_n630), .A3(new_n645), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n650), .A3(G14), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT75), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT74), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n659), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  INV_X1    g239(.A(new_n653), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n661), .A2(new_n653), .A3(new_n658), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT73), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n668), .A2(G2096), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G2096), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n661), .A2(new_n660), .B1(new_n663), .B2(new_n666), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n675), .B2(new_n671), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n620), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(G2096), .B1(new_n668), .B2(new_n672), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n674), .A3(new_n671), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n679), .A3(G2100), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT79), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n686), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(KEYINPUT77), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT76), .B(KEYINPUT20), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n694), .B1(new_n693), .B2(new_n697), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n683), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n693), .A2(new_n697), .ZN(new_n701));
  INV_X1    g276(.A(new_n694), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n704));
  INV_X1    g279(.A(new_n683), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT78), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1981), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n700), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n700), .B2(new_n706), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G4), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n602), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G1348), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G33), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n481), .A2(G139), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n721), .B(new_n722), .C1(new_n462), .C2(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT88), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT88), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n718), .B1(new_n727), .B2(new_n717), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(G2072), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT89), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  NOR2_X1   g306(.A1(G27), .A2(G29), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G164), .B2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT93), .B(G2078), .Z(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  NAND3_X1  g310(.A1(new_n712), .A2(KEYINPUT23), .A3(G20), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT23), .ZN(new_n737));
  INV_X1    g312(.A(G20), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G16), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n739), .C1(new_n606), .C2(new_n712), .ZN(new_n740));
  INV_X1    g315(.A(G1956), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n717), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n717), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n744), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n748));
  INV_X1    g323(.A(G26), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G29), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n479), .A2(G128), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n481), .A2(G140), .ZN(new_n753));
  OR2_X1    g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(new_n756), .B2(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n750), .B1(new_n757), .B2(new_n748), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT86), .B(G2067), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n742), .A2(new_n747), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G2072), .B2(new_n728), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n730), .A2(new_n731), .A3(new_n735), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(G160), .A2(G29), .ZN(new_n764));
  AND2_X1   g339(.A1(KEYINPUT24), .A2(G34), .ZN(new_n765));
  NOR2_X1   g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n717), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n758), .A2(new_n759), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  NAND2_X1  g348(.A1(G168), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G16), .B2(G21), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n770), .B(new_n772), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n773), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n626), .A2(new_n717), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n712), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n712), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1961), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT30), .B(G28), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n717), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n763), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n712), .A2(G22), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT83), .B(G1971), .Z(new_n788));
  OAI211_X1 g363(.A(new_n787), .B(new_n788), .C1(G166), .C2(new_n712), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(G166), .B2(new_n712), .ZN(new_n790));
  INV_X1    g365(.A(new_n788), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n712), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G288), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT33), .B(G1976), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT82), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n797), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n794), .B(new_n799), .C1(G288), .C2(G16), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n789), .B(new_n792), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  NAND2_X1  g377(.A1(G305), .A2(G16), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n712), .A2(G6), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n803), .A2(new_n804), .A3(new_n802), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT84), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n792), .A2(new_n789), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n803), .A2(new_n804), .A3(new_n802), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n805), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n795), .B(new_n797), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n810), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G25), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT80), .B1(new_n819), .B2(G29), .ZN(new_n820));
  OR3_X1    g395(.A1(new_n819), .A2(KEYINPUT80), .A3(G29), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n479), .A2(G119), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n481), .A2(G131), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n820), .B(new_n821), .C1(new_n827), .C2(new_n717), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G24), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(G16), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(KEYINPUT81), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(G16), .B1(new_n584), .B2(new_n586), .ZN(new_n836));
  INV_X1    g411(.A(new_n833), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT81), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G1986), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(G1986), .B(new_n835), .C1(new_n838), .C2(new_n839), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n818), .A2(new_n831), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT85), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n830), .B1(new_n816), .B2(new_n817), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT85), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n845), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n809), .A2(new_n815), .A3(KEYINPUT34), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n786), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n849), .B1(new_n848), .B2(new_n845), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT34), .B1(new_n809), .B2(new_n815), .ZN(new_n855));
  NOR4_X1   g430(.A1(new_n855), .A2(new_n844), .A3(KEYINPUT85), .A4(new_n830), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n786), .B(new_n852), .C1(new_n854), .C2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n716), .B(new_n785), .C1(new_n853), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n717), .A2(G32), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n469), .A2(new_n471), .A3(G141), .A4(new_n462), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT90), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n493), .A2(KEYINPUT90), .A3(G141), .A4(new_n462), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n469), .A2(new_n471), .A3(G129), .A4(G2105), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT91), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT91), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n493), .A2(new_n868), .A3(G129), .A4(G2105), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT26), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g448(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n616), .A2(G105), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n865), .A2(new_n870), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n860), .B1(new_n880), .B2(new_n717), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT27), .B(G1996), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT92), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n881), .B(new_n883), .Z(new_n884));
  NOR2_X1   g459(.A1(new_n553), .A2(new_n712), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n712), .B2(G19), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G1341), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n859), .A2(new_n884), .A3(new_n888), .ZN(G311));
  INV_X1    g464(.A(new_n785), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n851), .A2(new_n852), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT36), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n892), .B2(new_n857), .ZN(new_n893));
  INV_X1    g468(.A(new_n884), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n887), .A4(new_n716), .ZN(G150));
  OR2_X1    g470(.A1(new_n511), .A2(new_n512), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(G55), .A3(G543), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT95), .B(G93), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n505), .A3(new_n898), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n897), .B(new_n899), .C1(new_n900), .C2(new_n504), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n552), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n901), .A2(new_n546), .A3(new_n542), .A4(new_n551), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n602), .A2(G559), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n910));
  AOI21_X1  g485(.A(G860), .B1(new_n908), .B2(KEYINPUT39), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n908), .B2(KEYINPUT39), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT97), .Z(new_n914));
  NAND2_X1  g489(.A1(new_n901), .A2(G860), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT37), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(G145));
  NAND2_X1  g492(.A1(new_n479), .A2(G130), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n481), .A2(G142), .ZN(new_n919));
  NOR2_X1   g494(.A1(G106), .A2(G2105), .ZN(new_n920));
  OAI21_X1  g495(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n918), .B(new_n919), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G162), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n626), .B(G160), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n923), .B(new_n924), .Z(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n879), .A2(G164), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n877), .B1(new_n867), .B2(new_n869), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n502), .B1(new_n928), .B2(new_n865), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n756), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n879), .A2(G164), .ZN(new_n931));
  INV_X1    g506(.A(new_n756), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n502), .A3(new_n865), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n930), .A2(new_n724), .A3(new_n934), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n930), .A2(new_n934), .B1(new_n725), .B2(new_n726), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n618), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n934), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n727), .ZN(new_n939));
  INV_X1    g514(.A(new_n618), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n930), .A2(new_n724), .A3(new_n934), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n937), .A2(new_n942), .A3(new_n826), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n826), .B1(new_n937), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n926), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n935), .A2(new_n936), .A3(new_n618), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n827), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n937), .A2(new_n942), .A3(new_n826), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n925), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT98), .B(G37), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n945), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT99), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n945), .A2(new_n950), .A3(new_n955), .A4(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n902), .B2(G868), .ZN(new_n960));
  INV_X1    g535(.A(new_n600), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n597), .B(new_n592), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(G651), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n964));
  NAND2_X1  g539(.A1(G299), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n564), .A2(KEYINPUT100), .A3(new_n566), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n591), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n601), .A2(new_n964), .A3(G299), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n905), .B(new_n611), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(KEYINPUT41), .A3(new_n968), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT101), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n972), .A2(new_n969), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT101), .A4(new_n973), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  XNOR2_X1  g555(.A(G303), .B(G288), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(G305), .ZN(new_n982));
  INV_X1    g557(.A(G290), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(G305), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n982), .B2(new_n984), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n976), .A2(new_n989), .A3(new_n977), .A4(new_n978), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n980), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n980), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n960), .B1(new_n993), .B2(G868), .ZN(new_n994));
  INV_X1    g569(.A(G868), .ZN(new_n995));
  NOR4_X1   g570(.A1(new_n991), .A2(new_n992), .A3(new_n959), .A4(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(G295));
  NOR2_X1   g572(.A1(new_n994), .A2(new_n996), .ZN(G331));
  NAND2_X1  g573(.A1(new_n971), .A2(new_n973), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n525), .A2(new_n505), .B1(new_n527), .B2(G51), .ZN(new_n1000));
  NAND3_X1  g575(.A1(G301), .A2(new_n1000), .A3(new_n530), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G286), .A2(G171), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT104), .B1(new_n905), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n905), .A2(new_n1003), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n903), .A2(new_n1001), .A3(new_n904), .A4(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1007), .B2(KEYINPUT104), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT105), .B1(new_n999), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1006), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n903), .A2(new_n904), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT104), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1004), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n973), .A4(new_n971), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1007), .A2(new_n969), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1009), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n988), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1008), .A2(new_n968), .A3(new_n967), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n971), .A2(new_n973), .A3(new_n1007), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1020), .B(new_n1021), .C1(new_n986), .C2(new_n987), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1019), .A2(new_n952), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT44), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n988), .ZN(new_n1027));
  INV_X1    g602(.A(G37), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1022), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(KEYINPUT43), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1019), .A2(new_n1024), .A3(new_n952), .A4(new_n1022), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(KEYINPUT43), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n1035));
  OAI22_X1  g610(.A1(new_n1025), .A2(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(G397));
  XNOR2_X1  g611(.A(KEYINPUT106), .B(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n502), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n464), .A2(new_n466), .ZN(new_n1042));
  OAI21_X1  g617(.A(G2105), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n474), .A2(new_n475), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n462), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1045), .A3(G40), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n756), .B(G2067), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT107), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1050), .B2(new_n880), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1996), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT46), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT47), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n879), .B(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n826), .A2(new_n829), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n1063), .B(KEYINPUT124), .Z(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2067), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n932), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1048), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G290), .A2(G1986), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1047), .ZN(new_n1070));
  XOR2_X1   g645(.A(new_n1070), .B(KEYINPUT48), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n826), .A2(new_n829), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1062), .A2(new_n1072), .A3(new_n1063), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n1073), .B2(new_n1047), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1059), .A2(new_n1068), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n1076));
  INV_X1    g651(.A(G1384), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n502), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT50), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n502), .A2(new_n1080), .A3(new_n1077), .ZN(new_n1081));
  INV_X1    g656(.A(G40), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n473), .A2(new_n1082), .A3(new_n476), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1079), .A2(new_n769), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1077), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT45), .B1(new_n502), .B2(new_n1077), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1046), .ZN(new_n1087));
  OAI211_X1 g662(.A(G168), .B(new_n1084), .C1(new_n1087), .C2(G1966), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(KEYINPUT118), .A3(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT51), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(KEYINPUT118), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1084), .B1(new_n1087), .B2(G1966), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G286), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1091), .A2(new_n1097), .A3(KEYINPUT62), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n498), .A2(new_n500), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1100), .A2(new_n496), .B1(new_n493), .B2(new_n492), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1384), .B1(new_n1101), .B2(new_n489), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1083), .B(new_n1099), .C1(new_n1102), .C2(KEYINPUT45), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT109), .B(G1971), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1079), .A2(new_n1106), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1107));
  INV_X1    g682(.A(G2090), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1046), .B1(new_n1078), .B2(KEYINPUT50), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1106), .B1(new_n1110), .B2(new_n1081), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1105), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(G303), .A2(G8), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT55), .Z(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1103), .B2(G2078), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT119), .B(G1961), .Z(new_n1120));
  OAI21_X1  g695(.A(new_n1083), .B1(new_n1102), .B2(new_n1080), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n502), .A2(new_n1080), .A3(new_n1077), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1085), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1078), .A2(new_n1039), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1083), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1127), .A2(G2078), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1119), .B(new_n1123), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT110), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1105), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1080), .B1(new_n502), .B2(new_n1077), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1122), .A2(new_n1134), .A3(new_n1046), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1108), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1103), .A2(KEYINPUT110), .A3(new_n1104), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(G8), .A3(new_n1115), .ZN(new_n1139));
  NAND2_X1  g714(.A1(G305), .A2(G1981), .ZN(new_n1140));
  INV_X1    g715(.A(G1981), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(KEYINPUT111), .A2(KEYINPUT49), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1078), .A2(new_n1046), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1092), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1140), .A2(new_n1142), .B1(KEYINPUT111), .B2(KEYINPUT49), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1145), .B(new_n1147), .C1(new_n1148), .C2(new_n1144), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1102), .A2(new_n1083), .ZN(new_n1150));
  INV_X1    g725(.A(G1976), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1150), .B(G8), .C1(new_n1151), .C2(G288), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT52), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT52), .B1(G288), .B2(new_n1151), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1147), .B(new_n1154), .C1(new_n1151), .C2(G288), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1149), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1117), .A2(new_n1131), .A3(new_n1139), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1076), .B1(new_n1098), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1117), .A2(new_n1139), .A3(new_n1156), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(G8), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(new_n1163), .A3(new_n1090), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1160), .A2(new_n1164), .A3(KEYINPUT123), .A4(new_n1131), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT62), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1158), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1082), .B(new_n473), .C1(KEYINPUT121), .C2(new_n1045), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1128), .B1(new_n476), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1168), .A2(new_n1099), .A3(new_n1170), .A4(new_n1040), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1119), .A2(new_n1123), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(G171), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1129), .A2(G171), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1159), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1172), .A2(G171), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT54), .B1(new_n1181), .B2(new_n1130), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1162), .B2(new_n1090), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g759(.A1(G299), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n564), .A2(KEYINPUT57), .A3(new_n566), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(KEYINPUT56), .B(G2072), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1125), .A2(new_n1083), .A3(new_n1099), .A4(new_n1188), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1187), .B(new_n1189), .C1(new_n1135), .C2(G1956), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(G1348), .B1(new_n1110), .B2(new_n1081), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1150), .A2(G2067), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT115), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n715), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT115), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1146), .A2(new_n1066), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1194), .A2(new_n1198), .A3(new_n602), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1187), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1189), .ZN(new_n1201));
  AOI21_X1  g776(.A(G1956), .B1(new_n1110), .B2(new_n1081), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1191), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT116), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n741), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1187), .B1(new_n1207), .B2(new_n1189), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1191), .B2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1125), .A2(new_n1054), .A3(new_n1083), .A4(new_n1099), .ZN(new_n1210));
  XOR2_X1   g785(.A(KEYINPUT58), .B(G1341), .Z(new_n1211));
  NAND2_X1  g786(.A1(new_n1150), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT59), .B1(new_n1213), .B2(new_n553), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT59), .ZN(new_n1215));
  AOI211_X1 g790(.A(new_n1215), .B(new_n552), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1191), .A2(KEYINPUT117), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1206), .A2(KEYINPUT117), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1203), .A2(new_n1190), .A3(new_n1219), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1209), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n602), .B1(new_n1222), .B2(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(KEYINPUT60), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1222), .A2(KEYINPUT60), .A3(new_n602), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1221), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g802(.A(new_n1180), .B(new_n1183), .C1(new_n1205), .C2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1167), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1138), .A2(G8), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1230), .A2(new_n1116), .ZN(new_n1231));
  NAND4_X1  g806(.A1(new_n1095), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1232), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1231), .A2(new_n1139), .A3(new_n1156), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1234), .A2(KEYINPUT113), .ZN(new_n1235));
  AOI22_X1  g810(.A1(new_n1126), .A2(new_n773), .B1(new_n1135), .B2(new_n769), .ZN(new_n1236));
  NOR3_X1   g811(.A1(new_n1236), .A2(new_n1092), .A3(G286), .ZN(new_n1237));
  NAND4_X1  g812(.A1(new_n1117), .A2(new_n1139), .A3(new_n1156), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT63), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g815(.A(new_n1232), .B1(new_n1230), .B2(new_n1116), .ZN(new_n1241));
  INV_X1    g816(.A(KEYINPUT113), .ZN(new_n1242));
  NAND4_X1  g817(.A1(new_n1241), .A2(new_n1242), .A3(new_n1139), .A4(new_n1156), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n1235), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g819(.A(KEYINPUT114), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1139), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1247));
  OAI21_X1  g822(.A(new_n1142), .B1(new_n1247), .B2(G288), .ZN(new_n1248));
  AOI22_X1  g823(.A1(new_n1246), .A2(new_n1156), .B1(new_n1248), .B2(new_n1147), .ZN(new_n1249));
  NAND3_X1  g824(.A1(new_n1244), .A2(new_n1245), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1251), .A2(KEYINPUT114), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1229), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1073), .A2(new_n1047), .ZN(new_n1254));
  NOR2_X1   g829(.A1(new_n983), .A2(new_n841), .ZN(new_n1255));
  OAI21_X1  g830(.A(new_n1047), .B1(new_n1255), .B2(new_n1069), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  XOR2_X1   g832(.A(new_n1257), .B(KEYINPUT108), .Z(new_n1258));
  OAI21_X1  g833(.A(new_n1075), .B1(new_n1253), .B2(new_n1258), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g834(.A(KEYINPUT126), .ZN(new_n1261));
  INV_X1    g835(.A(new_n710), .ZN(new_n1262));
  NAND3_X1  g836(.A1(new_n700), .A2(new_n706), .A3(new_n708), .ZN(new_n1263));
  AOI21_X1  g837(.A(new_n460), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AND3_X1   g838(.A1(new_n651), .A2(new_n677), .A3(new_n680), .ZN(new_n1265));
  AOI21_X1  g839(.A(new_n1261), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g840(.A(G319), .B1(new_n709), .B2(new_n710), .ZN(new_n1267));
  NAND3_X1  g841(.A1(new_n651), .A2(new_n677), .A3(new_n680), .ZN(new_n1268));
  NOR3_X1   g842(.A1(new_n1267), .A2(new_n1268), .A3(KEYINPUT126), .ZN(new_n1269));
  NOR2_X1   g843(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g844(.A1(new_n957), .A2(new_n1033), .A3(new_n1270), .ZN(G225));
  NAND2_X1  g845(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1272));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1273));
  NAND4_X1  g847(.A1(new_n957), .A2(new_n1033), .A3(new_n1270), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g848(.A1(new_n1272), .A2(new_n1274), .ZN(G308));
endmodule


