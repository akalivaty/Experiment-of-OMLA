//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NOR2_X1   g0008(.A1(G58), .A2(G68), .ZN(new_n209));
  AND2_X1   g0009(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  NOR3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(G20), .A3(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n208), .B(new_n216), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G58), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  AOI21_X1  g0042(.A(KEYINPUT67), .B1(new_n242), .B2(new_n214), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n242), .A2(KEYINPUT67), .A3(new_n214), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G13), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G1), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  INV_X1    g0053(.A(G58), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT8), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(new_n255), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n250), .A2(new_n258), .B1(new_n260), .B2(new_n249), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G20), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT7), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  NOR4_X1   g0067(.A1(new_n262), .A2(new_n263), .A3(new_n267), .A4(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(G68), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G68), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n254), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(G20), .B1(new_n271), .B2(new_n209), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G159), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT16), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n246), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n269), .A2(KEYINPUT16), .A3(new_n276), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n261), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n284));
  OR3_X1    g0084(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n215), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(KEYINPUT66), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT66), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n290), .B(new_n256), .C1(G41), .C2(G45), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n288), .A2(new_n289), .A3(G232), .A4(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G223), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G1698), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT3), .B(G33), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n295), .A2(new_n296), .B1(G33), .B2(G87), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n285), .B(new_n292), .C1(new_n297), .C2(new_n288), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n296), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G87), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n282), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT70), .A2(G179), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT70), .A2(G179), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n304), .A2(new_n307), .A3(new_n292), .A4(new_n285), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT18), .B1(new_n281), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n298), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n304), .A2(new_n313), .A3(new_n292), .A4(new_n285), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n265), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n267), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n265), .A4(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n270), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n278), .B1(new_n321), .B2(new_n275), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n242), .A2(KEYINPUT67), .A3(new_n214), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n243), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n280), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n261), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n315), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT17), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n326), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n300), .A2(new_n308), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT18), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n315), .A2(new_n325), .A3(KEYINPUT17), .A4(new_n326), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n310), .A2(new_n329), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT80), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(G1698), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n296), .A2(G222), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n296), .A2(G223), .A3(G1698), .ZN(new_n341));
  INV_X1    g0141(.A(G77), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n296), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n282), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(G226), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n348), .A2(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT69), .B1(new_n201), .B2(new_n265), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n273), .A2(G150), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n201), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n252), .A2(new_n265), .A3(G33), .A4(new_n255), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n324), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n247), .A2(new_n265), .A3(G1), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n324), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n257), .A2(G50), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(new_n361), .B1(new_n212), .B2(new_n358), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n348), .A2(new_n307), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n349), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n311), .B1(new_n344), .B2(new_n347), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G190), .B2(new_n348), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT9), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n357), .A2(new_n368), .A3(new_n362), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n246), .B1(new_n354), .B2(new_n355), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n250), .A2(new_n360), .B1(G50), .B2(new_n249), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT9), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT10), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n367), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n373), .B2(new_n367), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n365), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(KEYINPUT71), .A2(G107), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT71), .A2(G107), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n288), .B1(new_n264), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G232), .A2(G1698), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n339), .A2(G238), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n296), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n288), .A2(new_n289), .A3(G244), .A4(new_n291), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n285), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n299), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G20), .A2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n265), .A2(G33), .ZN(new_n392));
  INV_X1    g0192(.A(new_n273), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n390), .B1(new_n391), .B2(new_n392), .C1(new_n393), .C2(new_n251), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n324), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n246), .A2(G77), .A3(new_n249), .A4(new_n257), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n249), .B2(G77), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n358), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n389), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT76), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n386), .A2(new_n307), .A3(new_n285), .A4(new_n387), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n345), .B1(new_n382), .B2(new_n385), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n408), .A2(KEYINPUT75), .A3(new_n307), .A4(new_n387), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n389), .A2(new_n401), .A3(KEYINPUT76), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n404), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n386), .A2(G190), .A3(new_n285), .A4(new_n387), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT72), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n388), .A2(G200), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT74), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n394), .A2(new_n324), .B1(new_n398), .B2(new_n399), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n396), .A4(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n311), .B1(new_n408), .B2(new_n387), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT74), .B1(new_n419), .B2(new_n401), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n337), .A2(new_n338), .A3(new_n377), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n294), .A2(new_n339), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n227), .A2(G1698), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n262), .C2(new_n263), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n427), .A2(KEYINPUT77), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT77), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n282), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT78), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(KEYINPUT78), .B(new_n282), .C1(new_n429), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n346), .A2(G238), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n285), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n424), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g0239(.A(KEYINPUT13), .B(new_n437), .C1(new_n433), .C2(new_n434), .ZN(new_n440));
  OAI21_X1  g0240(.A(G200), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n427), .A2(new_n428), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n427), .A2(KEYINPUT77), .A3(new_n428), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT78), .B1(new_n446), .B2(new_n282), .ZN(new_n447));
  INV_X1    g0247(.A(new_n434), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n438), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT13), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n435), .A2(new_n424), .A3(new_n438), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(G190), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n270), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n342), .B2(new_n392), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n324), .A2(new_n454), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(KEYINPUT11), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n358), .A2(new_n270), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT12), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(KEYINPUT11), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n359), .A2(G68), .A3(new_n257), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n456), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n441), .A2(new_n452), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT79), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n439), .A2(new_n440), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(G190), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT79), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(new_n441), .ZN(new_n468));
  OAI21_X1  g0268(.A(G169), .B1(new_n439), .B2(new_n440), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT14), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n450), .A2(G179), .A3(new_n451), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT14), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(G169), .C1(new_n439), .C2(new_n440), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n464), .A2(new_n468), .B1(new_n474), .B2(new_n461), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n423), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT85), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n242), .A2(new_n214), .B1(G20), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n265), .C1(G33), .C2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT20), .B1(new_n479), .B2(new_n482), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n483), .A2(new_n484), .B1(G116), .B2(new_n249), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n256), .A2(G33), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n249), .B(new_n486), .C1(new_n323), .C2(new_n243), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n478), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n477), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n249), .A2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n479), .A2(new_n482), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n246), .A2(G116), .A3(new_n249), .A4(new_n486), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(KEYINPUT85), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n256), .B(G45), .C1(new_n287), .C2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT81), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G41), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n256), .A4(G45), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G270), .A3(new_n288), .ZN(new_n507));
  OAI211_X1 g0307(.A(G264), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(new_n339), .C1(new_n262), .C2(new_n263), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n316), .A2(G303), .A3(new_n317), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n282), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n499), .A2(new_n500), .B1(KEYINPUT5), .B2(new_n287), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(G274), .A3(new_n288), .A4(new_n504), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n507), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(G169), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n498), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT21), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(KEYINPUT21), .A3(G169), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n507), .A2(new_n512), .A3(G179), .A4(new_n514), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n498), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n515), .A2(G200), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n507), .A2(new_n512), .A3(G190), .A4(new_n514), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(new_n489), .A3(new_n497), .A4(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n519), .B(new_n523), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n265), .B(G87), .C1(new_n262), .C2(new_n263), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n296), .A2(new_n532), .A3(new_n265), .A4(G87), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  INV_X1    g0335(.A(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(G20), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n478), .B2(new_n392), .ZN(new_n538));
  INV_X1    g0338(.A(new_n380), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(G20), .A3(new_n378), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(KEYINPUT23), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n534), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n534), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n324), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n248), .A2(G20), .A3(new_n536), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT25), .ZN(new_n547));
  INV_X1    g0347(.A(new_n487), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(G107), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n506), .A2(G264), .A3(new_n288), .ZN(new_n551));
  OAI211_X1 g0351(.A(G257), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n552));
  OAI211_X1 g0352(.A(G250), .B(new_n339), .C1(new_n262), .C2(new_n263), .ZN(new_n553));
  AND2_X1   g0353(.A1(KEYINPUT87), .A2(G294), .ZN(new_n554));
  NOR2_X1   g0354(.A1(KEYINPUT87), .A2(G294), .ZN(new_n555));
  OAI21_X1  g0355(.A(G33), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n282), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n551), .A2(new_n558), .A3(new_n514), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT88), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(G169), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n282), .B1(new_n513), .B2(new_n504), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(G264), .B1(new_n282), .B2(new_n557), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(G179), .A3(new_n514), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n560), .B1(new_n559), .B2(G169), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n550), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(G200), .B1(new_n563), .B2(new_n514), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n313), .A2(new_n551), .A3(new_n514), .A4(new_n558), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n545), .B(new_n549), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G244), .B(new_n339), .C1(new_n262), .C2(new_n263), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n480), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G250), .A2(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(KEYINPUT4), .A2(G244), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n575), .B1(new_n296), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n282), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n506), .A2(G257), .A3(new_n288), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n514), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT82), .B1(new_n583), .B2(G200), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n273), .A2(G77), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n536), .A2(KEYINPUT6), .A3(G97), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT6), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n586), .B1(new_n591), .B2(new_n265), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n381), .B1(new_n319), .B2(new_n320), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n324), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n548), .A2(G97), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n249), .A2(G97), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n583), .A2(KEYINPUT82), .A3(G200), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n581), .A2(G190), .A3(new_n514), .A4(new_n582), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n585), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G87), .A2(G97), .ZN(new_n602));
  NAND3_X1  g0402(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n381), .A2(new_n602), .B1(new_n265), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n265), .B(G68), .C1(new_n262), .C2(new_n263), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n392), .B2(new_n481), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n324), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n391), .A2(new_n358), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n609), .B(new_n610), .C1(new_n487), .C2(new_n391), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT83), .ZN(new_n612));
  INV_X1    g0412(.A(G45), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(G250), .C1(new_n613), .C2(G1), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n256), .A2(G45), .ZN(new_n615));
  AOI21_X1  g0415(.A(G274), .B1(KEYINPUT83), .B2(G250), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n288), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT84), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g0420(.A1(G238), .A2(G1698), .ZN(new_n621));
  INV_X1    g0421(.A(G244), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G1698), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n623), .C1(new_n262), .C2(new_n263), .ZN(new_n624));
  NAND2_X1  g0424(.A1(G33), .A2(G116), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n288), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n617), .A2(KEYINPUT84), .A3(new_n288), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n620), .A2(new_n627), .A3(new_n628), .A4(new_n307), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n617), .A2(KEYINPUT84), .A3(new_n288), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT84), .B1(new_n617), .B2(new_n288), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n630), .A2(new_n631), .A3(new_n626), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n611), .B(new_n629), .C1(new_n632), .C2(G169), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n620), .A2(new_n627), .A3(new_n628), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n246), .A2(G87), .A3(new_n249), .A4(new_n486), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n609), .A2(new_n636), .A3(new_n610), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n620), .A2(new_n627), .A3(G190), .A4(new_n628), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n381), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n266), .B2(new_n268), .ZN(new_n642));
  AND2_X1   g0442(.A1(G97), .A2(G107), .ZN(new_n643));
  NOR2_X1   g0443(.A1(G97), .A2(G107), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n589), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n587), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(G20), .B1(G77), .B2(new_n273), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n596), .B1(new_n648), .B2(new_n324), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n595), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n583), .A2(new_n299), .ZN(new_n651));
  INV_X1    g0451(.A(new_n514), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n288), .B1(new_n574), .B2(new_n579), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n307), .A3(new_n582), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n601), .A2(new_n640), .A3(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n476), .A2(new_n529), .A3(new_n571), .A4(new_n657), .ZN(G372));
  INV_X1    g0458(.A(new_n365), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT91), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n330), .A2(new_n332), .A3(new_n331), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n332), .B1(new_n330), .B2(new_n331), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n310), .A2(KEYINPUT91), .A3(new_n333), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n412), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n474), .A2(new_n461), .B1(new_n667), .B2(new_n463), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n329), .A2(new_n334), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n375), .A2(new_n376), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n659), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT89), .B1(new_n632), .B2(new_n311), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n634), .A2(new_n675), .A3(G200), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n638), .A3(new_n637), .A4(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n649), .A2(new_n595), .B1(new_n299), .B2(new_n583), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n633), .A3(new_n678), .A4(new_n655), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n640), .A2(KEYINPUT26), .A3(new_n655), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n567), .A2(new_n519), .A3(new_n523), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n570), .A2(new_n677), .A3(new_n633), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n600), .A2(new_n595), .A3(new_n594), .A4(new_n597), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n584), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n687), .A2(new_n599), .B1(new_n655), .B2(new_n678), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n633), .B(KEYINPUT90), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n683), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n423), .A2(new_n475), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n673), .A2(new_n692), .ZN(G369));
  XNOR2_X1  g0493(.A(KEYINPUT93), .B(G343), .ZN(new_n694));
  INV_X1    g0494(.A(G213), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n247), .A2(G1), .A3(G20), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n697), .B2(KEYINPUT27), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT92), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n696), .B2(new_n699), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n694), .B(new_n698), .C1(new_n701), .C2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT94), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT94), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n498), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n519), .A2(new_n523), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n529), .B2(new_n709), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n550), .A2(new_n707), .ZN(new_n715));
  INV_X1    g0515(.A(new_n707), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n571), .A2(new_n715), .B1(new_n567), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n710), .A2(new_n716), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(new_n571), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n567), .B2(new_n707), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n719), .A2(new_n722), .ZN(G399));
  INV_X1    g0523(.A(new_n206), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G41), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n256), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n381), .A2(new_n478), .A3(new_n602), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n726), .A2(new_n728), .B1(new_n213), .B2(new_n725), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n657), .A2(new_n571), .ZN(new_n732));
  INV_X1    g0532(.A(new_n529), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(new_n716), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n654), .A2(new_n632), .A3(new_n563), .A4(new_n582), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n521), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n632), .A2(new_n563), .ZN(new_n738));
  INV_X1    g0538(.A(new_n521), .ZN(new_n739));
  INV_X1    g0539(.A(new_n583), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT30), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n307), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n632), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n515), .A3(new_n559), .A4(new_n583), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n737), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n745), .B2(new_n707), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n731), .B1(new_n734), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT96), .ZN(new_n751));
  INV_X1    g0551(.A(new_n690), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n601), .A2(new_n656), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n570), .A2(new_n677), .A3(new_n633), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n755), .B2(new_n684), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n707), .B1(new_n756), .B2(new_n683), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n751), .B1(new_n757), .B2(KEYINPUT29), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n691), .A2(new_n716), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT29), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(KEYINPUT96), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n633), .A2(new_n639), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n763), .A2(new_n656), .A3(KEYINPUT26), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(KEYINPUT26), .B2(new_n679), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n689), .A3(new_n690), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(KEYINPUT29), .A3(new_n716), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n750), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n730), .B1(new_n768), .B2(G1), .ZN(G364));
  NAND2_X1  g0569(.A1(new_n265), .A2(G13), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G45), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n726), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n714), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G330), .B2(new_n712), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n724), .A2(new_n264), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G355), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G116), .B2(new_n206), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n237), .A2(new_n613), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n724), .A2(new_n296), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n213), .B2(new_n613), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n779), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n214), .B1(G20), .B2(new_n299), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n774), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n265), .A2(new_n311), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n742), .A2(G190), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(KEYINPUT99), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(KEYINPUT99), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G326), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n265), .A2(new_n313), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n742), .A2(new_n311), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(KEYINPUT98), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(KEYINPUT98), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G322), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n265), .A2(G190), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n311), .A2(G179), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G179), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G283), .A2(new_n809), .B1(new_n812), .B2(G329), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n554), .A2(new_n555), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n265), .B1(new_n810), .B2(G190), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n806), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n307), .A2(new_n817), .A3(G200), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(G311), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n799), .A2(new_n807), .ZN(new_n820));
  INV_X1    g0620(.A(G303), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n264), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT100), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n742), .A2(new_n313), .A3(new_n792), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n798), .A2(new_n805), .A3(new_n819), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G87), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n296), .B1(new_n808), .B2(new_n536), .C1(new_n829), .C2(new_n820), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G77), .B2(new_n818), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n270), .B2(new_n824), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n815), .A2(new_n481), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n811), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT32), .Z(new_n836));
  OR3_X1    g0636(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n212), .A2(new_n796), .B1(new_n803), .B2(new_n254), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n828), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n791), .B1(new_n839), .B2(new_n788), .ZN(new_n840));
  INV_X1    g0640(.A(new_n787), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n712), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n776), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  AND3_X1   g0644(.A1(new_n411), .A2(new_n407), .A3(new_n409), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n705), .A2(new_n706), .B1(new_n396), .B2(new_n417), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n845), .A2(KEYINPUT102), .A3(new_n404), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n412), .A2(new_n421), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n404), .A2(new_n410), .A3(new_n411), .A4(new_n846), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT102), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n847), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n759), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n847), .A2(new_n849), .A3(new_n852), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n691), .A2(new_n716), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n750), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n774), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  INV_X1    g0660(.A(new_n818), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n861), .A2(new_n478), .B1(new_n862), .B2(new_n824), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n264), .B1(new_n808), .B2(new_n829), .ZN(new_n864));
  INV_X1    g0664(.A(G311), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n820), .A2(new_n536), .B1(new_n811), .B2(new_n865), .ZN(new_n866));
  NOR4_X1   g0666(.A1(new_n863), .A2(new_n833), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(G294), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n867), .B1(new_n868), .B2(new_n803), .C1(new_n821), .C2(new_n796), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n825), .A2(G150), .B1(G159), .B2(new_n818), .ZN(new_n870));
  INV_X1    g0670(.A(G143), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n803), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G137), .B2(new_n797), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT34), .Z(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n875));
  INV_X1    g0675(.A(new_n815), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(G58), .ZN(new_n877));
  INV_X1    g0677(.A(new_n820), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n264), .B1(new_n878), .B2(G50), .ZN(new_n879));
  AOI22_X1  g0679(.A1(G68), .A2(new_n809), .B1(new_n812), .B2(G132), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n875), .A2(new_n877), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n869), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n788), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n788), .A2(new_n785), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n773), .B1(new_n342), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n884), .B(new_n886), .C1(new_n786), .C2(new_n855), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n860), .A2(new_n887), .ZN(G384));
  NOR3_X1   g0688(.A1(new_n214), .A2(new_n265), .A3(new_n478), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n646), .B(KEYINPUT103), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT35), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n213), .B(G77), .C1(new_n254), .C2(new_n270), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n897), .A2(KEYINPUT104), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n897), .A2(KEYINPUT104), .B1(new_n212), .B2(G68), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n256), .B(G13), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n701), .A2(new_n703), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n904), .A2(new_n698), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n330), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n335), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n330), .A2(new_n331), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n906), .A3(new_n327), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n909), .A2(new_n906), .A3(new_n912), .A4(new_n327), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n903), .B1(new_n335), .B2(new_n907), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n902), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n335), .A2(new_n907), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n919), .A2(KEYINPUT38), .A3(new_n914), .A4(new_n908), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n473), .A2(new_n471), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n450), .A2(new_n451), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n472), .B1(new_n923), .B2(G169), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n461), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n461), .A2(new_n707), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n466), .B2(new_n441), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n474), .B1(new_n468), .B2(new_n464), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n926), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n853), .B1(new_n734), .B2(new_n749), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n921), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n663), .A2(new_n669), .A3(new_n664), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n907), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n914), .ZN(new_n938));
  XOR2_X1   g0738(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n920), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n941), .A2(KEYINPUT40), .A3(new_n931), .A4(new_n932), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n476), .B1(new_n734), .B2(new_n749), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n731), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n412), .A2(new_n707), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n856), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n921), .A2(new_n931), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT39), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n915), .A2(new_n902), .A3(new_n916), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n940), .B1(new_n937), .B2(new_n914), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n920), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n474), .A2(new_n461), .A3(new_n716), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n950), .B1(new_n666), .B2(new_n905), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n463), .A2(new_n667), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n670), .B1(new_n925), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n672), .B1(new_n960), .B2(new_n665), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n365), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n767), .A2(new_n423), .A3(new_n475), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n962), .B1(new_n762), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n958), .B(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n946), .A2(new_n966), .B1(new_n256), .B2(new_n771), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT107), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n946), .A2(new_n966), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n967), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n901), .B1(new_n969), .B2(new_n971), .ZN(G367));
  NAND2_X1  g0772(.A1(new_n233), .A2(new_n781), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n973), .B(new_n789), .C1(new_n206), .C2(new_n391), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT109), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n774), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n974), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT110), .Z(new_n978));
  AOI22_X1  g0778(.A1(new_n825), .A2(G159), .B1(G50), .B2(new_n818), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT112), .B(G137), .Z(new_n980));
  OAI22_X1  g0780(.A1(new_n980), .A2(new_n811), .B1(new_n820), .B2(new_n254), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n808), .A2(new_n342), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n815), .A2(new_n270), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n264), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(G150), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n985), .B1(new_n871), .B2(new_n796), .C1(new_n986), .C2(new_n803), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G303), .A2(new_n804), .B1(new_n797), .B2(G311), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT111), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n878), .A2(KEYINPUT46), .A3(G116), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n820), .B2(new_n478), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(new_n824), .C2(new_n814), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n988), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n989), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n264), .B1(new_n811), .B2(new_n996), .C1(new_n481), .C2(new_n808), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n641), .B2(new_n876), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n995), .B(new_n998), .C1(new_n862), .C2(new_n861), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n987), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT47), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n788), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n978), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n677), .A2(new_n633), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n716), .A2(new_n637), .ZN(new_n1007));
  MUX2_X1   g0807(.A(new_n690), .B(new_n1006), .S(new_n1007), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1005), .B1(new_n841), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n772), .A2(G1), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT108), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n688), .B1(new_n598), .B2(new_n716), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n678), .A2(new_n655), .A3(new_n707), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n722), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT44), .Z(new_n1017));
  NOR2_X1   g0817(.A1(new_n722), .A2(new_n1015), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n719), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(new_n718), .A3(new_n1019), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n720), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n721), .B1(new_n717), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n713), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n768), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n725), .B(KEYINPUT41), .Z(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1012), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1015), .A2(new_n721), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT42), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n656), .B1(new_n1013), .B2(new_n567), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1031), .A2(KEYINPUT42), .B1(new_n716), .B2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1032), .A2(new_n1034), .B1(KEYINPUT43), .B2(new_n1009), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n718), .A2(new_n1015), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1010), .B1(new_n1030), .B2(new_n1039), .ZN(G387));
  INV_X1    g0840(.A(new_n1026), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n768), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n725), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n768), .B2(new_n1041), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n717), .A2(new_n841), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n230), .A2(new_n613), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1048), .A2(new_n781), .B1(new_n727), .B2(new_n777), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n251), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT114), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1051), .A2(KEYINPUT50), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(KEYINPUT50), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n728), .B(new_n613), .C1(new_n270), .C2(new_n342), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n536), .B2(new_n724), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n774), .B1(new_n1057), .B2(new_n790), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n861), .A2(new_n270), .B1(new_n259), .B2(new_n824), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n815), .A2(new_n391), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n296), .B1(new_n808), .B2(new_n481), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n820), .A2(new_n342), .B1(new_n811), .B2(new_n986), .ZN(new_n1062));
  NOR4_X1   g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n212), .B2(new_n803), .C1(new_n834), .C2(new_n796), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n296), .B1(new_n812), .B2(G326), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n820), .A2(new_n814), .B1(new_n815), .B2(new_n862), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n825), .A2(G311), .B1(G303), .B2(new_n818), .ZN(new_n1067));
  INV_X1    g0867(.A(G322), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n796), .B2(new_n1068), .C1(new_n996), .C2(new_n803), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1065), .B1(new_n478), .B2(new_n808), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1064), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1047), .B(new_n1058), .C1(new_n1076), .C2(new_n788), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1041), .A2(KEYINPUT113), .A3(new_n1012), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT113), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1012), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1026), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1046), .A2(new_n1082), .ZN(G393));
  INV_X1    g0883(.A(new_n1023), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1044), .B1(new_n1084), .B2(new_n1043), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1043), .B2(new_n1084), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1080), .B1(new_n1023), .B2(KEYINPUT115), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(KEYINPUT115), .B2(new_n1023), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1015), .A2(new_n787), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n789), .B1(new_n481), .B2(new_n206), .C1(new_n240), .C2(new_n782), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n774), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT116), .Z(new_n1092));
  OAI22_X1  g0892(.A1(new_n865), .A2(new_n803), .B1(new_n796), .B2(new_n996), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n878), .A2(G283), .B1(new_n812), .B2(G322), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n264), .C1(new_n536), .C2(new_n808), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT117), .Z(new_n1097));
  NAND2_X1  g0897(.A1(new_n818), .A2(G294), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n825), .A2(G303), .B1(G116), .B2(new_n876), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n986), .A2(new_n796), .B1(new_n803), .B2(new_n834), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT51), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n878), .A2(G68), .B1(new_n812), .B2(G143), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n296), .C1(new_n829), .C2(new_n808), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n861), .A2(new_n251), .B1(new_n212), .B2(new_n824), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n815), .A2(new_n342), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1094), .A2(new_n1100), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1089), .B(new_n1092), .C1(new_n1108), .C2(new_n1003), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1086), .A2(new_n1088), .A3(new_n1109), .ZN(G390));
  NOR4_X1   g0910(.A1(new_n529), .A2(new_n657), .A3(new_n571), .A4(new_n707), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n748), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n746), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n855), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n474), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n467), .B1(new_n466), .B2(new_n441), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n463), .A2(KEYINPUT79), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n927), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1114), .B1(new_n1119), .B2(new_n929), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n931), .A2(new_n949), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n957), .A2(new_n1121), .B1(new_n954), .B2(new_n955), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n957), .B1(new_n952), .B2(new_n953), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n707), .B1(new_n756), .B2(new_n765), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n855), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n948), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1126), .B2(new_n931), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n731), .B(new_n853), .C1(new_n734), .C2(new_n749), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n931), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n947), .B1(new_n1124), .B2(new_n855), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1118), .A2(new_n927), .B1(new_n925), .B2(new_n928), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n941), .B(new_n957), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n954), .A2(new_n955), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n957), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n931), .B2(new_n949), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1130), .B(new_n1133), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1128), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n750), .A2(new_n423), .A3(new_n475), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT96), .B1(new_n759), .B2(new_n760), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n751), .B(KEYINPUT29), .C1(new_n691), .C2(new_n716), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n767), .A2(new_n423), .A3(new_n475), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n673), .B(new_n1140), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1129), .A2(new_n931), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n949), .B1(new_n1146), .B2(new_n1120), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1119), .A2(new_n1114), .A3(new_n929), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1130), .A2(new_n1148), .A3(new_n1131), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1044), .B1(new_n1139), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT119), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT118), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1138), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1128), .A2(new_n1137), .A3(KEYINPUT118), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1130), .A2(new_n1148), .A3(new_n1131), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n949), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1130), .B2(new_n1148), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n964), .B(new_n1140), .C1(new_n1156), .C2(new_n1158), .ZN(new_n1159));
  AND4_X1   g0959(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .A4(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1150), .B1(new_n1138), .B2(new_n1153), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1152), .B1(new_n1161), .B2(new_n1155), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1151), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1139), .A2(new_n1012), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n885), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n264), .B1(new_n812), .B2(G125), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n212), .B2(new_n808), .C1(new_n834), .C2(new_n815), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n820), .A2(new_n986), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n824), .B2(new_n980), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT120), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1167), .B(new_n1170), .C1(new_n818), .C2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G128), .A2(new_n797), .B1(new_n804), .B2(G132), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n808), .A2(new_n270), .B1(new_n811), .B2(new_n868), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n264), .B1(new_n820), .B2(new_n829), .ZN(new_n1176));
  OR3_X1    g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n1106), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n861), .A2(new_n481), .B1(new_n381), .B2(new_n824), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n797), .C2(G283), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n804), .A2(G116), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1173), .A2(new_n1174), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n774), .B1(new_n260), .B2(new_n1165), .C1(new_n1181), .C2(new_n1003), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n956), .B2(new_n785), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT121), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n1164), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1163), .A2(new_n1186), .ZN(G378));
  OAI21_X1  g0987(.A(new_n774), .B1(G50), .B2(new_n1165), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n363), .A2(new_n905), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n672), .A2(new_n365), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n377), .A2(new_n363), .A3(new_n905), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(new_n786), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n861), .A2(new_n391), .B1(new_n481), .B2(new_n824), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n287), .B(new_n264), .C1(new_n820), .C2(new_n342), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n808), .A2(new_n254), .B1(new_n811), .B2(new_n862), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1198), .A2(new_n983), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n796), .B2(new_n478), .C1(new_n536), .C2(new_n803), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n264), .A2(new_n287), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G50), .B1(new_n286), .B2(new_n287), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1202), .A2(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G125), .A2(new_n797), .B1(new_n804), .B2(G128), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n818), .A2(G137), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n825), .A2(G132), .B1(G150), .B2(new_n876), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1172), .A2(new_n878), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT122), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT123), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n286), .B(new_n287), .C1(new_n808), .C2(new_n834), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G124), .B2(new_n812), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1206), .B1(new_n1203), .B2(new_n1202), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1188), .B(new_n1197), .C1(new_n788), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n731), .B1(new_n933), .B2(new_n934), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1221), .A2(new_n942), .A3(new_n1196), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1196), .B1(new_n1221), .B2(new_n942), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n958), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n935), .A2(new_n942), .A3(G330), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1196), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n950), .B1(new_n666), .B2(new_n905), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1135), .B2(new_n1134), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1221), .A2(new_n942), .A3(new_n1196), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1224), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1220), .B1(new_n1232), .B2(new_n1012), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1145), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1138), .B2(new_n1159), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(KEYINPUT57), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n725), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1233), .B1(new_n1237), .B2(new_n1238), .ZN(G375));
  NAND3_X1  g1039(.A1(new_n1145), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1159), .A2(new_n1029), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G128), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n820), .A2(new_n834), .B1(new_n811), .B2(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n861), .A2(new_n986), .B1(KEYINPUT124), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n825), .A2(new_n1172), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n264), .B1(new_n809), .B2(G58), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n212), .C2(new_n815), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1244), .B(new_n1247), .C1(KEYINPUT124), .C2(new_n1243), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n980), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G132), .A2(new_n797), .B1(new_n804), .B2(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n861), .A2(new_n381), .B1(new_n478), .B2(new_n824), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n820), .A2(new_n481), .B1(new_n811), .B2(new_n821), .ZN(new_n1252));
  OR4_X1    g1052(.A1(new_n296), .A2(new_n1252), .A3(new_n982), .A4(new_n1060), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1251), .B(new_n1253), .C1(new_n797), .C2(G294), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n804), .A2(G283), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1248), .A2(new_n1250), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n774), .B1(G68), .B2(new_n1165), .C1(new_n1256), .C2(new_n1003), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1132), .B2(new_n785), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n1012), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1241), .A2(new_n1260), .ZN(G381));
  NOR2_X1   g1061(.A1(G393), .A2(G396), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1260), .A3(new_n1241), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(G387), .A2(new_n1263), .A3(G390), .A4(G384), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1154), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT119), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1161), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1185), .B1(new_n1268), .B2(new_n1151), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT57), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n725), .A3(new_n1236), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1233), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1264), .A2(new_n1275), .ZN(G407));
  NOR2_X1   g1076(.A1(new_n694), .A2(new_n695), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(KEYINPUT125), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1240), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n725), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1159), .B2(new_n1240), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1260), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G384), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1286), .A2(KEYINPUT126), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(KEYINPUT126), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1285), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1145), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT60), .B1(new_n1290), .B2(new_n1150), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1044), .B1(new_n1240), .B2(new_n1281), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(KEYINPUT126), .A3(new_n1286), .A4(new_n1260), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1277), .A2(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1289), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT127), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1295), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1289), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1299), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1232), .A2(new_n1029), .A3(new_n1235), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1233), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1277), .B1(new_n1269), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G378), .A2(G375), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1305), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n843), .B1(new_n1046), .B2(new_n1082), .ZN(new_n1312));
  OAI221_X1 g1112(.A(new_n1010), .B1(new_n1039), .B2(new_n1030), .C1(new_n1262), .C2(new_n1312), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1262), .A2(new_n1312), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(G387), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1316), .A2(G390), .ZN(new_n1317));
  INV_X1    g1117(.A(G390), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1277), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1307), .A2(new_n1163), .A3(new_n1186), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1309), .A2(new_n1321), .A3(new_n1300), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  OR2_X1    g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1311), .A2(new_n1320), .A3(new_n1325), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1322), .A2(new_n1321), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1273), .A2(new_n1233), .B1(new_n1163), .B2(new_n1186), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1299), .B(new_n1304), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1308), .A2(new_n1333), .A3(new_n1300), .A4(new_n1309), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1328), .A2(new_n1329), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1316), .B(G390), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1327), .A2(new_n1337), .ZN(G405));
  INV_X1    g1138(.A(new_n1300), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1275), .A2(new_n1331), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1300), .B1(new_n1274), .B2(new_n1309), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1320), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1336), .B1(new_n1341), .B2(new_n1340), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(G402));
endmodule


