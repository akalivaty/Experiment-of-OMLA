//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(new_n192), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(new_n187), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT69), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  OR3_X1    g016(.A1(new_n202), .A2(KEYINPUT67), .A3(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(G134), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT67), .B1(new_n205), .B2(G137), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n203), .B(G131), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT64), .B1(new_n208), .B2(G143), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(G143), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT68), .A2(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT68), .A2(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n213), .A2(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n214), .A2(new_n220), .A3(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n207), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n202), .B2(G134), .ZN(new_n225));
  OAI22_X1  g039(.A1(new_n205), .A2(G137), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n202), .A4(G134), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n225), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n226), .ZN(new_n234));
  INV_X1    g048(.A(new_n225), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n223), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n230), .A2(new_n232), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n237), .B2(new_n233), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT0), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n221), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n213), .A2(new_n214), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT0), .B(G128), .Z(new_n245));
  AOI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n239), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n230), .A2(new_n232), .ZN(new_n249));
  AND4_X1   g063(.A1(new_n231), .A2(new_n234), .A3(new_n232), .A4(new_n235), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT70), .A3(new_n246), .ZN(new_n253));
  AOI211_X1 g067(.A(new_n201), .B(new_n238), .C1(new_n248), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n246), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n217), .A2(new_n218), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n244), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(new_n207), .C1(new_n250), .C2(new_n251), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n255), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n238), .B1(new_n248), .B2(new_n253), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n254), .B1(new_n264), .B2(new_n201), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G210), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n267), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n271), .B(new_n272), .Z(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n255), .A2(new_n261), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n201), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n276), .B2(new_n201), .ZN(new_n279));
  INV_X1    g093(.A(new_n201), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n263), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n277), .B(new_n279), .C1(new_n281), .C2(new_n278), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n274), .B(new_n275), .C1(new_n273), .C2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT74), .B(G902), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n241), .A2(new_n247), .A3(new_n239), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT70), .B1(new_n252), .B2(new_n246), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n261), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n201), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n281), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT28), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n291), .A2(new_n279), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n273), .A2(new_n275), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n285), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n283), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G472), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n264), .A2(new_n201), .ZN(new_n297));
  INV_X1    g111(.A(new_n273), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT73), .B(KEYINPUT31), .Z(new_n299));
  NAND4_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n281), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n282), .A2(new_n273), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n273), .B(new_n254), .C1(new_n264), .C2(new_n201), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT31), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT72), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n262), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n288), .B2(KEYINPUT30), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n298), .B(new_n281), .C1(new_n307), .C2(new_n280), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT31), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n302), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G472), .A2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n311), .A2(KEYINPUT32), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT32), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n279), .A2(new_n277), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n298), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n303), .B2(new_n299), .ZN(new_n319));
  AOI211_X1 g133(.A(KEYINPUT72), .B(new_n304), .C1(new_n265), .C2(new_n298), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n309), .B1(new_n308), .B2(KEYINPUT31), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n322), .B2(new_n312), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n296), .B1(new_n314), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n284), .B2(G234), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n217), .A2(new_n189), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT75), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n329));
  INV_X1    g143(.A(G128), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(G119), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n328), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n327), .A2(KEYINPUT23), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT23), .B1(new_n330), .B2(G119), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n189), .B2(G128), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n332), .A2(new_n334), .B1(new_n338), .B2(G110), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n340), .A2(KEYINPUT16), .A3(G140), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n208), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n339), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n332), .A2(new_n334), .B1(new_n338), .B2(G110), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n343), .B(new_n208), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n353), .A3(new_n357), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT25), .B1(new_n362), .B2(new_n284), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n361), .A2(new_n364), .A3(new_n285), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n326), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n326), .A2(G902), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G214), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n371), .A2(G237), .A3(G953), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G143), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT84), .B(G143), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT18), .A3(G131), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n375), .A2(new_n372), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT18), .A2(G131), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  OR3_X1    g194(.A1(new_n342), .A2(KEYINPUT85), .A3(new_n208), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT85), .B1(new_n342), .B2(new_n208), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n377), .B(new_n380), .C1(new_n347), .C2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n342), .B(KEYINPUT19), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n208), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n374), .B(new_n232), .C1(new_n372), .C2(new_n375), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n232), .B1(new_n378), .B2(new_n374), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n386), .B(new_n344), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n376), .A2(G131), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n387), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n389), .A2(KEYINPUT17), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n351), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n394), .A3(new_n384), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(G475), .A2(G902), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT20), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  INV_X1    g222(.A(G902), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n401), .A2(new_n394), .A3(new_n384), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n394), .B1(new_n401), .B2(new_n384), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT86), .B(G475), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n406), .A2(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n415));
  INV_X1    g229(.A(G122), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G116), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n191), .A2(G122), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT77), .B(G107), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n215), .A2(G143), .A3(new_n216), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n211), .A2(G128), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n205), .A3(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n422), .A2(KEYINPUT13), .A3(new_n423), .ZN(new_n425));
  OAI21_X1  g239(.A(G134), .B1(new_n423), .B2(KEYINPUT13), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n421), .B(new_n424), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n419), .A2(new_n420), .ZN(new_n428));
  INV_X1    g242(.A(new_n424), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n205), .B1(new_n422), .B2(new_n423), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G107), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n191), .A2(G122), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n418), .B1(new_n434), .B2(KEYINPUT14), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(KEYINPUT87), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(new_n418), .C1(new_n434), .C2(KEYINPUT14), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n432), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n427), .B1(new_n431), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT9), .B(G234), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n441), .A2(new_n325), .A3(G953), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n415), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n431), .A2(new_n439), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(KEYINPUT88), .A3(new_n427), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n443), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G478), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(KEYINPUT15), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n284), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n448), .B2(new_n284), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G952), .ZN(new_n456));
  AOI211_X1 g270(.A(G953), .B(new_n456), .C1(G234), .C2(G237), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n269), .B(new_n284), .C1(G234), .C2(G237), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(KEYINPUT21), .B(G898), .Z(new_n461));
  OAI21_X1  g275(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n414), .A2(new_n455), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n432), .A2(G104), .ZN(new_n464));
  OR2_X1    g278(.A1(KEYINPUT77), .A2(G107), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT77), .A2(G107), .ZN(new_n466));
  AOI21_X1  g280(.A(G104), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT78), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n420), .A2(new_n468), .A3(new_n393), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G101), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT1), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(G143), .B2(new_n208), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n211), .A2(G146), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n208), .A2(G143), .ZN(new_n476));
  OAI22_X1  g290(.A1(new_n474), .A2(new_n330), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n214), .A2(new_n220), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT79), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n479), .B(new_n480), .C1(new_n330), .C2(new_n474), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n259), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT3), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n432), .B2(G104), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n464), .ZN(new_n485));
  INV_X1    g299(.A(G101), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(G104), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n485), .B(new_n486), .C1(new_n420), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n472), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n485), .B1(new_n420), .B2(new_n487), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G101), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n488), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n495), .A3(G101), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n246), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n472), .A2(new_n260), .A3(KEYINPUT10), .A4(new_n488), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n491), .A2(new_n241), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G110), .B(G140), .ZN(new_n500));
  INV_X1    g314(.A(G227), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G953), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n500), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT80), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n499), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n497), .A2(new_n498), .ZN(new_n509));
  INV_X1    g323(.A(new_n488), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n420), .A2(new_n393), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT78), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n464), .A3(new_n470), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n513), .B2(G101), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT10), .B1(new_n514), .B2(new_n482), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n252), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n508), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n489), .B1(new_n514), .B2(new_n260), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT12), .B1(new_n518), .B2(new_n252), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n219), .A2(new_n222), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n393), .A2(G107), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n511), .B2(KEYINPUT78), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n486), .B1(new_n523), .B2(new_n470), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n521), .B1(new_n524), .B2(new_n510), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n520), .B(new_n241), .C1(new_n525), .C2(new_n489), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n499), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n503), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n409), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G469), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n516), .A2(new_n499), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n503), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n499), .B(new_n504), .C1(new_n519), .C2(new_n526), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n285), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT81), .ZN(new_n536));
  INV_X1    g350(.A(G469), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n531), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G221), .B1(new_n441), .B2(G902), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n494), .A2(new_n200), .A3(new_n199), .A4(new_n496), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT5), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n546), .B(G113), .C1(new_n547), .C2(new_n195), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n472), .A2(new_n194), .A3(new_n488), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G110), .B(G122), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n549), .A3(new_n551), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT6), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n521), .A2(new_n556), .A3(new_n340), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT82), .B1(new_n260), .B2(G125), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n246), .A2(new_n340), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G224), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G953), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n562), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT6), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n550), .A2(new_n565), .A3(new_n552), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n555), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT7), .B1(new_n561), .B2(G953), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n557), .B(new_n568), .C1(new_n558), .C2(new_n559), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n554), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n568), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n560), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n551), .B(KEYINPUT8), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n548), .A2(new_n194), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(new_n524), .B2(new_n510), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n575), .B2(new_n549), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT83), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI211_X1 g392(.A(KEYINPUT83), .B(new_n573), .C1(new_n575), .C2(new_n549), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n570), .B(new_n572), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n567), .A2(new_n580), .A3(new_n409), .ZN(new_n581));
  OAI21_X1  g395(.A(G210), .B1(G237), .B2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n576), .B(new_n577), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n572), .A2(new_n554), .A3(new_n569), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n582), .A3(new_n567), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n544), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  AND4_X1   g403(.A1(new_n463), .A2(new_n541), .A3(new_n542), .A4(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n324), .A2(new_n370), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  OR2_X1    g406(.A1(new_n442), .A2(KEYINPUT89), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n440), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n440), .A2(new_n593), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT33), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n448), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n597), .A2(new_n599), .A3(G478), .A4(new_n284), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n448), .A2(new_n284), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT90), .B1(new_n601), .B2(new_n449), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT90), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n603), .B(G478), .C1(new_n448), .C2(new_n284), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n600), .B(KEYINPUT91), .C1(new_n602), .C2(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n412), .A2(new_n413), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n611));
  INV_X1    g425(.A(new_n404), .ZN(new_n612));
  AOI211_X1 g426(.A(KEYINPUT20), .B(new_n612), .C1(new_n396), .C2(new_n402), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n581), .A2(new_n583), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n582), .B1(new_n587), .B2(new_n567), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n462), .B(new_n543), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n322), .A2(new_n312), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n533), .A2(new_n534), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n537), .A3(new_n284), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT81), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n623), .A2(new_n538), .B1(new_n530), .B2(G469), .ZN(new_n624));
  INV_X1    g438(.A(new_n542), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n624), .A2(new_n369), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n311), .B2(new_n285), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n619), .A2(new_n620), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n620), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n611), .A2(new_n613), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n454), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n452), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n618), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n632), .A2(new_n626), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND2_X1  g457(.A1(new_n623), .A2(new_n538), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n625), .B1(new_n644), .B2(new_n531), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n354), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n367), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n366), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g463(.A1(new_n463), .A2(new_n645), .A3(new_n589), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n632), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n283), .B2(new_n294), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT32), .B1(new_n311), .B2(new_n313), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n322), .A2(new_n315), .A3(new_n312), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT93), .B(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n459), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n458), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n455), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n645), .A2(new_n663), .A3(new_n589), .A4(new_n649), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n330), .ZN(G30));
  NAND2_X1  g480(.A1(new_n656), .A2(new_n657), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n290), .A2(new_n298), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n266), .B2(new_n298), .ZN(new_n669));
  AOI21_X1  g483(.A(G902), .B1(new_n669), .B2(KEYINPUT94), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(KEYINPUT94), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G472), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n667), .A2(KEYINPUT95), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT95), .B1(new_n667), .B2(new_n672), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n661), .B(KEYINPUT39), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n645), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n616), .A2(new_n617), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT38), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n414), .A2(new_n455), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n682), .A2(new_n544), .A3(new_n649), .A4(new_n684), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n676), .A2(new_n679), .A3(new_n680), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n211), .ZN(G45));
  INV_X1    g501(.A(new_n661), .ZN(new_n688));
  AOI211_X1 g502(.A(new_n414), .B(new_n688), .C1(new_n607), .C2(new_n608), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n645), .A3(new_n589), .A4(new_n649), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n658), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n208), .ZN(G48));
  NOR2_X1   g506(.A1(new_n658), .A2(new_n369), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT96), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n518), .A2(new_n252), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n520), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n518), .A2(KEYINPUT12), .A3(new_n252), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n505), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n698), .A2(new_n699), .B1(new_n532), .B2(new_n503), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n694), .B1(new_n700), .B2(new_n285), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n621), .A2(KEYINPUT96), .A3(new_n284), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(G469), .A3(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n703), .B(new_n542), .C1(new_n539), .C2(new_n540), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT97), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n644), .A2(KEYINPUT97), .A3(new_n542), .A4(new_n703), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n693), .A2(new_n619), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND3_X1  g525(.A1(new_n693), .A2(new_n640), .A3(new_n708), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  AND2_X1   g527(.A1(new_n649), .A2(new_n463), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n589), .A2(new_n706), .A3(new_n707), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n324), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NOR2_X1   g531(.A1(new_n618), .A2(new_n684), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n706), .A2(new_n707), .A3(new_n718), .ZN(new_n719));
  OAI221_X1 g533(.A(new_n300), .B1(new_n304), .B2(new_n303), .C1(new_n292), .C2(new_n298), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n312), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n627), .A2(new_n721), .A3(new_n370), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n416), .ZN(G24));
  NAND4_X1  g538(.A1(new_n706), .A2(new_n589), .A3(new_n689), .A4(new_n707), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n627), .A2(new_n721), .A3(new_n649), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n340), .ZN(G27));
  OAI21_X1  g542(.A(KEYINPUT99), .B1(new_n658), .B2(new_n369), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n324), .A2(new_n730), .A3(new_n370), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT98), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n584), .A2(new_n588), .A3(new_n732), .A4(new_n543), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n584), .A2(new_n588), .A3(new_n543), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT98), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n645), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n689), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n729), .A2(new_n731), .A3(new_n739), .ZN(new_n740));
  AND4_X1   g554(.A1(new_n542), .A2(new_n541), .A3(new_n733), .A4(new_n735), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n324), .A2(new_n370), .A3(new_n741), .A4(new_n689), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n738), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NOR3_X1   g559(.A1(new_n658), .A2(new_n736), .A3(new_n369), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n663), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT100), .B(G134), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G36));
  INV_X1    g563(.A(new_n529), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n750), .B2(KEYINPUT45), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT101), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(KEYINPUT45), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT102), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT103), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n537), .A2(new_n409), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n644), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n542), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n677), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n614), .B1(new_n607), .B2(new_n608), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(KEYINPUT43), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n631), .A3(new_n649), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT44), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n735), .A2(new_n733), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT105), .Z(new_n777));
  NAND4_X1  g591(.A1(new_n766), .A2(new_n774), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  XNOR2_X1  g593(.A(new_n764), .B(KEYINPUT47), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n324), .A2(new_n370), .A3(new_n737), .A4(new_n776), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT106), .Z(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NAND2_X1  g599(.A1(new_n644), .A2(new_n703), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT49), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n682), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n767), .A2(new_n370), .A3(new_n542), .A4(new_n543), .ZN(new_n789));
  OAI221_X1 g603(.A(new_n788), .B1(KEYINPUT107), .B2(new_n789), .C1(KEYINPUT49), .C2(new_n786), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(KEYINPUT107), .B2(new_n789), .ZN(new_n791));
  INV_X1    g605(.A(new_n676), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n658), .B1(new_n664), .B2(new_n690), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n727), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n645), .A2(new_n589), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n796), .A2(new_n649), .A3(new_n688), .A4(new_n684), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n674), .B2(new_n675), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n795), .A2(new_n798), .A3(KEYINPUT52), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI211_X1 g616(.A(KEYINPUT111), .B(KEYINPUT52), .C1(new_n795), .C2(new_n798), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n689), .A2(new_n627), .A3(new_n721), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n636), .A2(new_n455), .A3(new_n661), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n658), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n736), .B1(new_n366), .B2(new_n648), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n663), .A2(new_n746), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n744), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n591), .A2(new_n813), .A3(new_n628), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n813), .B1(new_n591), .B2(new_n628), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n715), .A2(new_n324), .B1(new_n632), .B2(new_n650), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n455), .A2(new_n614), .A3(KEYINPUT109), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT109), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n414), .B2(new_n638), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n618), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n626), .A2(new_n620), .A3(new_n627), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n719), .B2(new_n722), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n817), .A2(new_n825), .A3(new_n709), .A4(new_n712), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n812), .A2(new_n816), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n804), .B2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n709), .A2(new_n817), .A3(new_n712), .A4(new_n825), .ZN(new_n829));
  INV_X1    g643(.A(new_n815), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n591), .A2(new_n813), .A3(new_n628), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n744), .A3(new_n832), .A4(new_n811), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n795), .A2(new_n798), .A3(KEYINPUT52), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n799), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT54), .B1(new_n828), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n838), .A2(KEYINPUT112), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n827), .B(KEYINPUT53), .C1(new_n802), .C2(new_n803), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n836), .B1(new_n833), .B2(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n838), .A2(new_n843), .A3(KEYINPUT112), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n708), .A2(new_n457), .A3(new_n733), .A4(new_n735), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n792), .A2(new_n370), .A3(new_n847), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n848), .A2(new_n614), .A3(new_n609), .ZN(new_n849));
  INV_X1    g663(.A(new_n722), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n771), .A3(new_n457), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n544), .A2(new_n852), .A3(new_n682), .A4(new_n708), .ZN(new_n853));
  XOR2_X1   g667(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n854));
  OR2_X1    g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(KEYINPUT114), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n847), .A2(new_n771), .ZN(new_n858));
  INV_X1    g672(.A(new_n726), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n849), .A2(new_n855), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT47), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n764), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n764), .A2(new_n864), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n644), .A2(new_n625), .A3(new_n703), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(KEYINPUT115), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n777), .A3(new_n852), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT115), .B1(new_n780), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n852), .A2(new_n777), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n867), .B(KEYINPUT113), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n780), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n862), .B1(new_n874), .B2(new_n861), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n729), .A2(new_n731), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n858), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT48), .Z(new_n878));
  NOR2_X1   g692(.A1(new_n456), .A2(G953), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n708), .A2(new_n589), .ZN(new_n880));
  OAI221_X1 g694(.A(new_n879), .B1(new_n880), .B2(new_n851), .C1(new_n848), .C2(new_n615), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n871), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n845), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(G952), .A2(G953), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n793), .B1(new_n884), .B2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n269), .A2(G952), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT117), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n555), .A2(new_n566), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n563), .A2(new_n564), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n567), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT55), .Z(new_n894));
  AOI21_X1  g708(.A(new_n284), .B1(new_n840), .B2(new_n841), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n582), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT116), .B(new_n894), .C1(new_n897), .C2(KEYINPUT56), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n889), .B1(new_n901), .B2(new_n902), .ZN(G51));
  NOR2_X1   g717(.A1(new_n896), .A2(new_n756), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT119), .Z(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n843), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n842), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n757), .B(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n621), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n887), .B1(new_n905), .B2(new_n912), .ZN(G54));
  INV_X1    g727(.A(new_n887), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n403), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n403), .B2(new_n915), .ZN(G60));
  AND2_X1   g731(.A1(new_n597), .A2(new_n599), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT59), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n845), .B2(new_n920), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n918), .A2(new_n908), .A3(new_n909), .A4(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n889), .A3(new_n922), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n325), .A2(new_n409), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n840), .B2(new_n841), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n647), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n842), .A2(new_n927), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n889), .B1(new_n933), .B2(new_n361), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n930), .A2(new_n931), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n924), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n888), .A2(KEYINPUT61), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n929), .B2(new_n647), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT122), .B1(new_n933), .B2(new_n361), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n929), .A2(new_n942), .A3(new_n362), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n938), .B(new_n940), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n933), .A2(KEYINPUT122), .A3(new_n361), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n929), .B2(new_n362), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n938), .B1(new_n948), .B2(new_n940), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n937), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT124), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n937), .B(new_n952), .C1(new_n945), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(G66));
  AOI21_X1  g768(.A(new_n269), .B1(new_n461), .B2(G224), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n816), .A2(new_n826), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(new_n269), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n890), .B1(G898), .B2(new_n269), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(G69));
  NOR2_X1   g774(.A1(new_n780), .A2(new_n783), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n686), .A2(new_n727), .A3(new_n794), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n765), .B1(new_n615), .B2(new_n821), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n746), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT125), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT126), .B1(new_n778), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n778), .A2(KEYINPUT126), .A3(new_n967), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n307), .B(new_n385), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n269), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n501), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n269), .B1(new_n973), .B2(G900), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n766), .A2(new_n589), .A3(new_n683), .A4(new_n876), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n744), .A2(new_n747), .A3(new_n795), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n778), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n269), .B1(new_n977), .B2(new_n961), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n971), .B1(new_n501), .B2(G953), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n972), .A2(new_n980), .ZN(G72));
  OAI211_X1 g795(.A(new_n964), .B(new_n956), .C1(new_n968), .C2(new_n969), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  AOI211_X1 g798(.A(new_n273), .B(new_n265), .C1(new_n982), .C2(new_n984), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n977), .A2(new_n961), .A3(new_n957), .ZN(new_n986));
  INV_X1    g800(.A(new_n984), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n273), .B(new_n265), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n274), .B(KEYINPUT127), .Z(new_n989));
  OAI221_X1 g803(.A(new_n984), .B1(new_n303), .B2(new_n989), .C1(new_n828), .C2(new_n837), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n988), .A2(new_n914), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n985), .A2(new_n991), .ZN(G57));
endmodule


