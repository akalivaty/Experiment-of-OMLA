//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT65), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n463), .ZN(new_n476));
  NAND3_X1  g051(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  NAND2_X1  g054(.A1(G101), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n473), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n478), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n485), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n476), .B2(new_n477), .ZN(new_n494));
  NAND2_X1  g069(.A1(G102), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n473), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n476), .B2(new_n477), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(G114), .B2(G2104), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n467), .B2(new_n470), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n497), .B(new_n503), .C1(new_n505), .C2(KEYINPUT4), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(KEYINPUT67), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n508));
  AND3_X1   g083(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n510));
  OAI211_X1 g085(.A(KEYINPUT4), .B(G138), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(G2105), .B1(new_n511), .B2(new_n495), .ZN(new_n512));
  OAI21_X1  g087(.A(G126), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n473), .B1(new_n513), .B2(new_n501), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT65), .ZN(new_n516));
  AOI21_X1  g091(.A(KEYINPUT65), .B1(new_n468), .B2(new_n469), .ZN(new_n517));
  OAI21_X1  g092(.A(G138), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n500), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n508), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n507), .A2(new_n520), .ZN(G164));
  NAND2_X1  g096(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(G543), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(G62), .ZN(new_n534));
  NAND2_X1  g109(.A1(G75), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n532), .A2(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  INV_X1    g113(.A(new_n528), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(new_n531), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n540), .A2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  INV_X1    g123(.A(G52), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n528), .A2(new_n548), .B1(new_n549), .B2(new_n531), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n526), .A2(G64), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n533), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n528), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n526), .A2(G56), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n533), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n531), .ZN(new_n560));
  AOI211_X1 g135(.A(new_n556), .B(new_n559), .C1(G43), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT69), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(KEYINPUT70), .A2(G53), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n531), .A2(KEYINPUT9), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n531), .B2(new_n568), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n569), .A2(new_n570), .B1(G91), .B2(new_n539), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n533), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n528), .A2(new_n576), .B1(new_n577), .B2(new_n531), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n578), .A2(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n533), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n528), .A2(new_n584), .B1(new_n585), .B2(new_n531), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  XNOR2_X1  g163(.A(KEYINPUT72), .B(G85), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n539), .A2(new_n589), .B1(G47), .B2(new_n560), .ZN(new_n590));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n523), .A2(new_n525), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n526), .A2(G92), .A3(new_n527), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT73), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n592), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n560), .B2(G54), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT74), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n602), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n602), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XOR2_X1   g200(.A(KEYINPUT75), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT76), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n465), .A2(G2105), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n471), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT77), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n487), .A2(G123), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT78), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n484), .A2(G135), .ZN(new_n637));
  NOR2_X1   g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G2096), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n633), .A2(new_n634), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT79), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n649), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT80), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(G2072), .A2(G2078), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n442), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n662), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT83), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n664), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n661), .B(new_n670), .C1(new_n667), .C2(new_n665), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT82), .Z(new_n672));
  NOR3_X1   g247(.A1(new_n661), .A2(new_n667), .A3(new_n664), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n641), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n680), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT84), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n689), .B(new_n691), .Z(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT85), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G4), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n613), .B2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT91), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(G1348), .Z(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(G32), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT26), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n708), .A2(new_n709), .B1(G105), .B2(new_n628), .ZN(new_n710));
  INV_X1    g285(.A(G141), .ZN(new_n711));
  INV_X1    g286(.A(G129), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n710), .B1(new_n483), .B2(new_n711), .C1(new_n712), .C2(new_n486), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n699), .A2(G5), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G171), .B2(new_n699), .ZN(new_n718));
  AND2_X1   g293(.A1(KEYINPUT24), .A2(G34), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n704), .B1(KEYINPUT24), .B2(G34), .ZN(new_n720));
  OAI22_X1  g295(.A1(G160), .A2(new_n704), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n716), .B1(G1961), .B2(new_n718), .C1(new_n721), .C2(G2084), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT98), .Z(new_n723));
  NOR2_X1   g298(.A1(G27), .A2(G29), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G164), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2078), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(G168), .A2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT96), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G21), .ZN(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n704), .A2(G35), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G162), .B2(new_n704), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT29), .Z(new_n735));
  OAI22_X1  g310(.A1(new_n730), .A2(new_n731), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G28), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT30), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n737), .B2(KEYINPUT30), .ZN(new_n739));
  OR2_X1    g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n640), .B2(new_n704), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n718), .B2(G1961), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n699), .A2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n561), .B2(new_n699), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT92), .B(G1341), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n484), .A2(G140), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n487), .A2(G128), .ZN(new_n750));
  NOR2_X1   g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(new_n473), .B2(G116), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n704), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n721), .A2(G2084), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n744), .A2(new_n748), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n735), .A2(new_n732), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n699), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1956), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n714), .A2(new_n715), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT95), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n762), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n736), .A2(new_n761), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n730), .A2(new_n731), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(new_n473), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  INV_X1    g351(.A(G139), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n483), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT93), .Z(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT94), .B(G2072), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n772), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n703), .A2(new_n727), .A3(new_n770), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n699), .A2(G22), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G166), .B2(new_n699), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1971), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n699), .A2(G6), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n587), .B2(new_n699), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n788), .B1(G1981), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G1981), .B2(new_n791), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n699), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(G288), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n699), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT87), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT34), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n793), .A2(KEYINPUT34), .A3(new_n799), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n699), .A2(G24), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n600), .B2(new_n699), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1986), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT86), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n484), .A2(G131), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n487), .A2(G119), .ZN(new_n808));
  NOR2_X1   g383(.A1(G95), .A2(G2105), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(G29), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n805), .A2(KEYINPUT86), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n806), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n802), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(KEYINPUT88), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT88), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n802), .B2(new_n817), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n800), .B(new_n801), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n800), .B1(new_n819), .B2(new_n821), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n822), .A2(KEYINPUT90), .B1(new_n823), .B2(KEYINPUT36), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(KEYINPUT88), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n825), .A2(new_n826), .A3(new_n800), .A4(new_n801), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n785), .B1(new_n824), .B2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n822), .A2(KEYINPUT90), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n785), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(G150));
  NOR2_X1   g408(.A1(new_n612), .A2(new_n620), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n539), .A2(G93), .B1(G55), .B2(new_n560), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT100), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n533), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(new_n561), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n836), .B(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n845), .A2(new_n846), .A3(G860), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(G860), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n506), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n515), .A2(KEYINPUT101), .A3(new_n519), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(new_n753), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n780), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n713), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n487), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(G106), .A2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(G142), .B2(new_n484), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n811), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n630), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n640), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n864), .B(KEYINPUT102), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n865), .B(new_n868), .C1(new_n857), .C2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(KEYINPUT103), .B(G37), .Z(new_n871));
  XOR2_X1   g446(.A(new_n857), .B(new_n869), .Z(new_n872));
  OAI211_X1 g447(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n868), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g449(.A(new_n600), .B(new_n795), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G305), .B(G303), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n877), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(KEYINPUT108), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT42), .Z(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n612), .A2(new_n617), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT104), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n613), .A2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n612), .A2(new_n891), .A3(new_n617), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n886), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT41), .A4(new_n892), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n842), .B(new_n622), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n890), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n900), .A2(KEYINPUT106), .A3(KEYINPUT41), .A4(new_n892), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n892), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n898), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT105), .Z(new_n905));
  AND3_X1   g480(.A1(new_n885), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n885), .B1(new_n905), .B2(new_n902), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n841), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(G868), .B2(new_n909), .ZN(G295));
  OAI21_X1  g485(.A(new_n908), .B1(G868), .B2(new_n909), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  XNOR2_X1  g487(.A(G286), .B(G171), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n842), .A2(KEYINPUT109), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n843), .A2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n842), .A2(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n897), .A2(new_n901), .A3(new_n915), .A4(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n916), .A2(new_n918), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n903), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n883), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n883), .B1(new_n920), .B2(new_n922), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n912), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n921), .B1(new_n894), .B2(new_n895), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n919), .A2(new_n915), .B1(new_n892), .B2(new_n900), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n882), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(new_n923), .A3(KEYINPUT43), .A4(new_n871), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT44), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n925), .B2(new_n926), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n930), .A2(new_n923), .A3(new_n912), .A4(new_n871), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n938), .ZN(G397));
  NOR2_X1   g514(.A1(new_n854), .A2(G1384), .ZN(new_n940));
  INV_X1    g515(.A(new_n481), .ZN(new_n941));
  OAI211_X1 g516(.A(G40), .B(new_n941), .C1(new_n472), .C2(new_n473), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n940), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n753), .B(new_n758), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT110), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n713), .B(G1996), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n813), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n811), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n753), .A2(G2067), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n811), .B(new_n813), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(G290), .A2(G1986), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n943), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n959));
  AOI22_X1  g534(.A1(new_n955), .A2(new_n943), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n953), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n943), .B1(new_n946), .B2(new_n713), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n944), .A2(G1996), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(KEYINPUT46), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(KEYINPUT46), .B2(new_n964), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT125), .Z(new_n967));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n962), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n968), .B2(new_n967), .ZN(new_n970));
  INV_X1    g545(.A(new_n942), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT45), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n497), .A2(new_n503), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT4), .B1(new_n471), .B2(G138), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT67), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n515), .A2(new_n508), .A3(new_n519), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n971), .B(new_n973), .C1(new_n978), .C2(KEYINPUT45), .ZN(new_n979));
  INV_X1    g554(.A(G1971), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n506), .A2(new_n972), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n942), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n972), .B1(new_n507), .B2(new_n520), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT111), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n978), .A2(new_n988), .A3(new_n984), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n981), .B1(new_n990), .B2(G2090), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n942), .A2(new_n982), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT112), .B(G8), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT113), .B(G1981), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n587), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(G1981), .B1(new_n583), .B2(new_n586), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1001), .A2(KEYINPUT114), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT114), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n995), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n795), .A2(G1976), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(G288), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n995), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n995), .A2(new_n1006), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1005), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT55), .Z(new_n1014));
  NAND3_X1  g589(.A1(new_n992), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1005), .A2(new_n1007), .A3(new_n795), .ZN(new_n1016));
  INV_X1    g591(.A(new_n998), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n995), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT63), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n991), .A2(G8), .A3(new_n1014), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1014), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n942), .B1(KEYINPUT50), .B2(new_n982), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1026), .A2(new_n732), .B1(new_n979), .B2(new_n980), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1022), .B1(new_n1027), .B2(new_n994), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1021), .A2(new_n1028), .A3(new_n1012), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2084), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(new_n985), .C1(new_n987), .C2(new_n989), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n942), .B1(new_n1033), .B2(new_n982), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n986), .B2(new_n1033), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n731), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n994), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G168), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1020), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1021), .A2(new_n1012), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1038), .A2(new_n1020), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1040), .B(new_n1041), .C1(new_n1014), .C2(new_n992), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1019), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G168), .A2(new_n994), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1046), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT120), .B(new_n1049), .C1(new_n1032), .C2(new_n1036), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1047), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OR3_X1    g629(.A1(new_n1037), .A2(KEYINPUT51), .A3(new_n1046), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT62), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(KEYINPUT62), .A3(new_n1055), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n979), .B2(G2078), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT122), .B(new_n1058), .C1(new_n979), .C2(G2078), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1961), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1035), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n990), .A2(new_n1064), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G301), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1057), .A2(new_n1069), .A3(new_n1029), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1043), .B1(new_n1056), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n617), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G299), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n973), .A2(new_n971), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n986), .A2(new_n1033), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1080), .A2(new_n1084), .A3(KEYINPUT116), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT116), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1078), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n985), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n986), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n988), .B1(new_n978), .B2(new_n984), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(G1348), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n993), .A2(new_n758), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1087), .B1(new_n612), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1078), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1080), .A2(new_n1097), .A3(new_n1084), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT60), .B(new_n1093), .C1(new_n1091), .C2(G1348), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(KEYINPUT118), .A3(new_n612), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT60), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1100), .A2(KEYINPUT118), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n612), .B1(new_n1100), .B2(KEYINPUT118), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1083), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n979), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n978), .A2(new_n984), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1956), .B1(new_n1110), .B2(new_n1024), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1078), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT61), .B1(new_n1112), .B2(new_n1098), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1098), .A2(KEYINPUT61), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1087), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n979), .B2(G1996), .ZN(new_n1117));
  INV_X1    g692(.A(G1996), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1081), .A2(KEYINPUT117), .A3(new_n1082), .A4(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n942), .B2(new_n982), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n561), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT59), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1125), .A3(new_n561), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1115), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1099), .B1(new_n1107), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT119), .B(new_n1099), .C1(new_n1107), .C2(new_n1128), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1054), .A2(new_n1055), .A3(new_n1029), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1063), .A2(new_n1068), .A3(G301), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n990), .A2(new_n1064), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1081), .B(new_n1067), .C1(KEYINPUT45), .C2(new_n940), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1062), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1082), .A2(new_n1066), .A3(new_n971), .A4(new_n973), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT122), .B1(new_n1140), .B2(new_n1058), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1137), .B(new_n1138), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1135), .A2(new_n1136), .B1(new_n1142), .B2(G171), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1063), .A2(new_n1068), .A3(KEYINPUT123), .A4(G301), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1134), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1142), .A2(G171), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1146), .A2(KEYINPUT54), .A3(new_n1069), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1133), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1131), .A2(new_n1132), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1071), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(G290), .A2(G1986), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n955), .A2(new_n956), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n944), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n970), .B1(new_n1152), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g731(.A1(G227), .A2(new_n460), .A3(G401), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n1158), .A2(new_n697), .ZN(new_n1159));
  XOR2_X1   g733(.A(new_n1159), .B(KEYINPUT127), .Z(new_n1160));
  NAND3_X1  g734(.A1(new_n936), .A2(new_n1160), .A3(new_n873), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


