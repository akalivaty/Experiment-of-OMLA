//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(G50), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n215), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G169), .ZN(new_n245));
  AND2_X1   g0045(.A1(G1), .A2(G13), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G264), .A3(G1698), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G303), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT85), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  OAI211_X1 g0061(.A(G257), .B(new_n261), .C1(new_n256), .C2(new_n257), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n255), .B(new_n259), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n262), .A2(new_n260), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n249), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT5), .B(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G274), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n249), .B1(new_n266), .B2(new_n268), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(G270), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n245), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT67), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n276), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n218), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n209), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G116), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n209), .B2(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n281), .A2(new_n284), .A3(new_n282), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT86), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n281), .A2(KEYINPUT86), .A3(new_n284), .A4(new_n282), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n283), .A2(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(G20), .B1(G33), .B2(G283), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n251), .A2(G97), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n291), .A2(new_n292), .B1(G20), .B2(new_n284), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n278), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n278), .A2(new_n293), .A3(KEYINPUT20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n290), .A2(KEYINPUT87), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT87), .B1(new_n290), .B2(new_n298), .ZN(new_n300));
  OAI211_X1 g0100(.A(KEYINPUT21), .B(new_n273), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n265), .A2(G179), .A3(new_n272), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n283), .A2(new_n285), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n288), .A2(new_n289), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT87), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n290), .A2(KEYINPUT87), .A3(new_n298), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n265), .A2(new_n272), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n265), .B2(new_n272), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n311), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT21), .B1(new_n311), .B2(new_n273), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n304), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n275), .A2(new_n277), .A3(new_n321), .A4(new_n218), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  INV_X1    g0124(.A(G50), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n210), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT69), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n210), .A2(G33), .ZN(new_n329));
  INV_X1    g0129(.A(G150), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G20), .A2(G33), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n323), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n323), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n209), .A2(G20), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT70), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n335), .A2(G50), .A3(new_n279), .A4(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n334), .B(new_n339), .C1(G50), .C2(new_n279), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT9), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n267), .A2(KEYINPUT66), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT66), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G45), .ZN(new_n344));
  INV_X1    g0144(.A(G41), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n209), .A2(G274), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n267), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n209), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n248), .ZN(new_n351));
  INV_X1    g0151(.A(G226), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n258), .A2(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G222), .ZN(new_n355));
  INV_X1    g0155(.A(G77), .ZN(new_n356));
  INV_X1    g0156(.A(G223), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n254), .A2(G1698), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n355), .B1(new_n356), .B2(new_n254), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n353), .B1(new_n359), .B2(new_n249), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n315), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(G190), .B2(new_n360), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n341), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(G190), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(KEYINPUT72), .C1(new_n315), .C2(new_n360), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n341), .B(new_n362), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n360), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n371), .B(new_n340), .C1(G169), .C2(new_n360), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n337), .A2(new_n202), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT74), .B(KEYINPUT12), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n281), .A2(new_n282), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(G68), .ZN(new_n377));
  INV_X1    g0177(.A(G13), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(G1), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT12), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(G20), .A4(new_n202), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n283), .A2(new_n374), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n331), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n356), .B2(new_n329), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n323), .A2(KEYINPUT11), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT11), .B1(new_n323), .B2(new_n384), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G238), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n348), .B1(new_n351), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n352), .A2(new_n261), .ZN(new_n391));
  INV_X1    g0191(.A(G232), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n391), .B(new_n393), .C1(new_n256), .C2(new_n257), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G97), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n248), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT13), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT73), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT73), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(KEYINPUT13), .C1(new_n390), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n395), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n249), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n209), .A2(new_n349), .B1(new_n246), .B2(new_n247), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(G238), .B1(new_n346), .B2(new_n347), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n398), .A2(G179), .A3(new_n400), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n397), .A2(new_n406), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT14), .B1(new_n408), .B2(G169), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT14), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n410), .B(new_n245), .C1(new_n397), .C2(new_n406), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT75), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT75), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n407), .C1(new_n409), .C2(new_n411), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n388), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n328), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n331), .B1(G20), .B2(G77), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n329), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n376), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n420), .A2(new_n278), .B1(new_n356), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n283), .A2(G77), .A3(new_n338), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G244), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n348), .B1(new_n351), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n354), .A2(G232), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n427), .B1(new_n206), .B2(new_n254), .C1(new_n389), .C2(new_n358), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n428), .B2(new_n249), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n424), .B1(new_n429), .B2(G190), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n315), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n370), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n424), .C1(G169), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n398), .A2(G190), .A3(new_n400), .A4(new_n406), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n408), .A2(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n388), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n416), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g0239(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n440));
  NAND3_X1  g0240(.A1(new_n252), .A2(new_n210), .A3(new_n253), .ZN(new_n441));
  AND2_X1   g0241(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n442));
  NOR2_X1   g0242(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n253), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n202), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G58), .A2(G68), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT78), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G58), .A3(G68), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n451), .A3(new_n203), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G20), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n331), .A2(G159), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n440), .B1(new_n447), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n452), .A2(G20), .B1(G159), .B2(new_n331), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n458), .A2(KEYINPUT16), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n202), .B1(new_n441), .B2(KEYINPUT7), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n256), .A2(new_n257), .A3(G20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n444), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n460), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n440), .C1(new_n447), .C2(new_n455), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n457), .A2(new_n466), .A3(new_n278), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n337), .A2(new_n328), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(new_n279), .A3(new_n320), .A4(new_n322), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n279), .B2(new_n417), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n404), .A2(G232), .B1(new_n346), .B2(new_n347), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n352), .A2(G1698), .ZN(new_n476));
  OAI221_X1 g0276(.A(new_n476), .B1(G223), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G87), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G179), .B(new_n475), .C1(new_n479), .C2(new_n248), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n348), .B1(new_n351), .B2(new_n392), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n248), .B1(new_n477), .B2(new_n478), .ZN(new_n482));
  OAI21_X1  g0282(.A(G169), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n474), .A2(KEYINPUT18), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n484), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n469), .B2(new_n473), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(KEYINPUT81), .A3(KEYINPUT18), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n474), .A2(new_n484), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT18), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n481), .A2(new_n482), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n313), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G200), .B2(new_n495), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n469), .A2(new_n473), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT17), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n373), .A2(new_n439), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n258), .A2(G20), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT22), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(G87), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n254), .A2(new_n210), .A3(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT22), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n329), .A2(new_n284), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT88), .B1(new_n210), .B2(G107), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n511), .A2(KEYINPUT23), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(KEYINPUT23), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n508), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n508), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n278), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n279), .A2(G107), .ZN(new_n518));
  XOR2_X1   g0318(.A(new_n518), .B(KEYINPUT25), .Z(new_n519));
  NAND2_X1  g0319(.A1(new_n209), .A2(G33), .ZN(new_n520));
  AND4_X1   g0320(.A1(new_n279), .A2(new_n320), .A3(new_n520), .A4(new_n322), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n521), .B2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n271), .A2(G264), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(new_n261), .C1(new_n256), .C2(new_n257), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n526));
  XOR2_X1   g0326(.A(KEYINPUT89), .B(G294), .Z(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n251), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n249), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(new_n529), .A3(new_n269), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n245), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n524), .A2(new_n529), .A3(new_n370), .A4(new_n269), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n523), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n315), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G190), .B2(new_n530), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n517), .A3(new_n522), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n521), .A2(G97), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT6), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT6), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n206), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n207), .A2(new_n543), .A3(new_n545), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(G20), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n331), .A2(G77), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n206), .B1(new_n445), .B2(new_n446), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n278), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n279), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n205), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n541), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G244), .B(new_n261), .C1(new_n256), .C2(new_n257), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n249), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n270), .B1(new_n271), .B2(G257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n245), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n370), .A3(new_n567), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n558), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n210), .B1(new_n395), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G87), .B2(new_n207), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n329), .B2(new_n205), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n254), .A2(new_n210), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n202), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n278), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n421), .A2(new_n419), .ZN(new_n579));
  INV_X1    g0379(.A(new_n521), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n419), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n347), .A2(G45), .ZN(new_n582));
  OAI21_X1  g0382(.A(G250), .B1(new_n267), .B2(G1), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n249), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G116), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n389), .A2(G1698), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n256), .B2(new_n257), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n254), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n249), .B1(new_n594), .B2(KEYINPUT84), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  INV_X1    g0396(.A(new_n588), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT84), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n370), .B(new_n585), .C1(new_n595), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n597), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT84), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n248), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n594), .A2(KEYINPUT84), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n584), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n581), .B(new_n599), .C1(new_n604), .C2(G169), .ZN(new_n605));
  OAI211_X1 g0405(.A(G190), .B(new_n585), .C1(new_n595), .C2(new_n598), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n578), .A2(new_n579), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(G87), .B2(new_n521), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n606), .B(new_n608), .C1(new_n604), .C2(new_n315), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n445), .A2(new_n446), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n552), .B(new_n551), .C1(new_n610), .C2(new_n206), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n278), .B1(new_n205), .B2(new_n556), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n566), .A2(new_n313), .A3(new_n567), .ZN(new_n613));
  AOI21_X1  g0413(.A(G200), .B1(new_n566), .B2(new_n567), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n612), .B(new_n541), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n571), .A2(new_n605), .A3(new_n609), .A4(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n319), .A2(new_n502), .A3(new_n540), .A4(new_n616), .ZN(G372));
  NOR2_X1   g0417(.A1(new_n304), .A2(new_n318), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n535), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n538), .A3(new_n616), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n558), .A2(new_n569), .A3(new_n570), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n605), .A2(new_n609), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT90), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n605), .A2(new_n609), .A3(new_n621), .A4(KEYINPUT26), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(KEYINPUT90), .A3(new_n623), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n620), .A2(new_n627), .A3(new_n605), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n502), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT91), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n438), .A2(new_n433), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n499), .B1(new_n416), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n493), .A2(new_n485), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n369), .A3(new_n368), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n372), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n631), .A2(new_n637), .ZN(G369));
  NAND2_X1  g0438(.A1(new_n379), .A2(new_n210), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n311), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n319), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n618), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n644), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n517), .B2(new_n522), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n539), .A2(new_n651), .B1(new_n535), .B2(new_n650), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n618), .A2(new_n644), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n540), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n533), .B1(new_n517), .B2(new_n522), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n650), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n213), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G41), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G1), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n217), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(new_n662), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n319), .A2(new_n616), .A3(new_n540), .A4(new_n650), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n524), .A2(new_n566), .A3(new_n529), .A4(new_n567), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n604), .A2(new_n669), .A3(new_n302), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT30), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n604), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n530), .A2(new_n370), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n312), .A4(new_n568), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n604), .A2(new_n669), .A3(new_n302), .A4(KEYINPUT30), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n644), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n668), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n615), .A2(new_n571), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n538), .A3(new_n605), .A4(new_n609), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n304), .A2(new_n318), .A3(new_n656), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n605), .B(new_n628), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n650), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  XNOR2_X1  g0490(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n689), .B2(new_n692), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n605), .B1(new_n685), .B2(new_n686), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n624), .A2(new_n626), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n644), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n683), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n667), .B1(new_n701), .B2(G1), .ZN(G364));
  NOR2_X1   g0502(.A1(new_n647), .A2(G330), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT94), .Z(new_n704));
  NOR2_X1   g0504(.A1(new_n378), .A2(G20), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n209), .B1(new_n705), .B2(G45), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n662), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n648), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n707), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n213), .A2(new_n254), .ZN(new_n710));
  INV_X1    g0510(.A(G355), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n710), .A2(new_n711), .B1(G116), .B2(new_n213), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n240), .A2(new_n267), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n213), .A2(new_n258), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n342), .A2(new_n344), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n217), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n712), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n218), .B1(G20), .B2(new_n245), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n709), .B1(new_n717), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n313), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n370), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n205), .ZN(new_n729));
  NOR4_X1   g0529(.A1(new_n210), .A2(new_n370), .A3(new_n315), .A4(G190), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(G68), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT96), .Z(new_n732));
  NOR2_X1   g0532(.A1(new_n210), .A2(G179), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(G190), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(G87), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n210), .A2(new_n370), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n313), .A3(G200), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n738), .A2(new_n325), .B1(new_n739), .B2(new_n206), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G190), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G159), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n736), .B(new_n740), .C1(KEYINPUT32), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n737), .A2(new_n741), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n254), .B1(new_n356), .B2(new_n747), .C1(new_n745), .C2(KEYINPUT32), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n737), .A2(new_n725), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT95), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n748), .B1(G58), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n732), .A2(new_n746), .A3(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n734), .B(KEYINPUT97), .Z(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G329), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n258), .B1(new_n742), .B2(new_n762), .C1(new_n763), .C2(new_n747), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n755), .B2(G322), .ZN(new_n765));
  INV_X1    g0565(.A(new_n738), .ZN(new_n766));
  INV_X1    g0566(.A(new_n739), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G326), .A2(new_n766), .B1(new_n767), .B2(G283), .ZN(new_n768));
  INV_X1    g0568(.A(new_n730), .ZN(new_n769));
  OR2_X1    g0569(.A1(KEYINPUT33), .A2(G317), .ZN(new_n770));
  NAND2_X1  g0570(.A1(KEYINPUT33), .A2(G317), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n527), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n727), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n765), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n757), .B1(new_n761), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n724), .B1(new_n776), .B2(new_n721), .ZN(new_n777));
  INV_X1    g0577(.A(new_n720), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n647), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n708), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT98), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n780), .B(new_n781), .ZN(G396));
  NOR2_X1   g0582(.A1(new_n721), .A2(new_n718), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n709), .B1(G77), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n769), .A2(new_n786), .B1(new_n739), .B2(new_n735), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n729), .B(new_n787), .C1(G303), .C2(new_n766), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n258), .B1(new_n742), .B2(new_n763), .C1(new_n284), .C2(new_n747), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n755), .B2(G294), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n790), .C1(new_n206), .C2(new_n759), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT99), .Z(new_n792));
  INV_X1    g0592(.A(new_n747), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n766), .A2(G137), .B1(new_n793), .B2(G159), .ZN(new_n794));
  INV_X1    g0594(.A(G143), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n330), .B2(new_n769), .C1(new_n754), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT34), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n254), .B1(new_n742), .B2(new_n800), .C1(new_n202), .C2(new_n739), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G58), .B2(new_n727), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n799), .B(new_n802), .C1(new_n325), .C2(new_n759), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n792), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n785), .B1(new_n804), .B2(new_n721), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n424), .A2(new_n644), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n431), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n433), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n433), .A2(new_n644), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n805), .B1(new_n811), .B2(new_n719), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT100), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n689), .A2(new_n810), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n434), .A2(new_n644), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n687), .B2(new_n688), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n814), .A2(new_n683), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n707), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT101), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n683), .B1(new_n816), .B2(new_n814), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n818), .B2(KEYINPUT101), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n813), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G384));
  NAND2_X1  g0623(.A1(new_n548), .A2(new_n550), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT102), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT35), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(KEYINPUT35), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(G116), .A4(new_n219), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT36), .Z(new_n829));
  NAND4_X1  g0629(.A1(new_n217), .A2(G77), .A3(new_n451), .A4(new_n449), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n325), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n209), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G330), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n466), .A2(new_n323), .ZN(new_n836));
  INV_X1    g0636(.A(new_n440), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT7), .ZN(new_n838));
  OAI21_X1  g0638(.A(G68), .B1(new_n462), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n441), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT77), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n460), .A2(new_n463), .A3(new_n461), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n837), .B1(new_n844), .B2(new_n458), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n473), .B1(new_n836), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n642), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n484), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n498), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT37), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT103), .ZN(new_n852));
  INV_X1    g0652(.A(new_n468), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n458), .A2(KEYINPUT16), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n842), .B2(new_n843), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n278), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n456), .B2(KEYINPUT80), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n472), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n852), .B1(new_n859), .B2(new_n488), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT37), .B1(new_n859), .B2(new_n497), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n642), .B1(new_n469), .B2(new_n473), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n489), .A2(KEYINPUT103), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n860), .A2(new_n861), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n851), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(KEYINPUT38), .B(new_n866), .C1(new_n500), .C2(new_n848), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n848), .B1(new_n494), .B2(new_n499), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n489), .B(new_n852), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n498), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n862), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n870), .A2(new_n873), .B1(new_n850), .B2(KEYINPUT37), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n868), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n413), .A2(new_n415), .ZN(new_n877));
  INV_X1    g0677(.A(new_n388), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n644), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n437), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n878), .B(new_n644), .C1(new_n877), .C2(new_n438), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n682), .A2(new_n883), .A3(new_n811), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n835), .B1(new_n876), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n863), .B1(new_n634), .B2(new_n499), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n863), .A2(new_n498), .A3(new_n491), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n865), .A2(KEYINPUT105), .B1(KEYINPUT37), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n873), .A2(new_n889), .A3(new_n860), .A4(new_n864), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n867), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n892));
  AND4_X1   g0692(.A1(KEYINPUT40), .A2(new_n682), .A3(new_n883), .A4(new_n811), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n885), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n502), .A2(new_n682), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n834), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n501), .B1(new_n699), .B2(KEYINPUT29), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n693), .B2(new_n694), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n637), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n860), .A2(new_n864), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n863), .A2(new_n871), .A3(new_n498), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT105), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n890), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n886), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n869), .A2(new_n874), .A3(new_n868), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n416), .A2(new_n650), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT104), .Z(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n867), .A2(new_n875), .A3(KEYINPUT39), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n634), .A2(new_n847), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n881), .A2(new_n882), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n816), .B2(new_n809), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n919), .B2(new_n876), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n901), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n898), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n209), .B2(new_n705), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n898), .A2(new_n922), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n833), .B1(new_n924), .B2(new_n925), .ZN(G367));
  NAND2_X1  g0726(.A1(new_n558), .A2(new_n644), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n684), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n621), .A2(new_n644), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n655), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n571), .B1(new_n928), .B2(new_n535), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n933), .A2(KEYINPUT42), .B1(new_n650), .B2(new_n935), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n605), .A2(new_n608), .A3(new_n650), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n605), .B(new_n609), .C1(new_n608), .C2(new_n650), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n934), .A2(new_n936), .B1(KEYINPUT43), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n653), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n930), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n661), .B(new_n946), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n655), .A2(new_n657), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n931), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT45), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n931), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n943), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n653), .A3(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT108), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n655), .B1(new_n652), .B2(new_n654), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n648), .B(new_n959), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n701), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n957), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n701), .A2(KEYINPUT108), .A3(new_n960), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n947), .B1(new_n964), .B2(new_n701), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n706), .B(KEYINPUT109), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n945), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n722), .B1(new_n213), .B2(new_n419), .C1(new_n236), .C2(new_n714), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n738), .A2(new_n795), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n728), .A2(new_n202), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(G159), .C2(new_n730), .ZN(new_n972));
  INV_X1    g0772(.A(new_n742), .ZN(new_n973));
  AOI22_X1  g0773(.A1(G50), .A2(new_n793), .B1(new_n973), .B2(G137), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n201), .B2(new_n734), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G150), .B2(new_n755), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n254), .B1(new_n739), .B2(new_n356), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n972), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n739), .A2(new_n205), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n769), .A2(new_n527), .B1(new_n763), .B2(new_n738), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(G107), .C2(new_n727), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n734), .B2(new_n284), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n258), .B1(new_n742), .B2(new_n986), .C1(new_n786), .C2(new_n747), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n755), .B2(G303), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n758), .A2(KEYINPUT46), .A3(G116), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n983), .A2(new_n985), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  INV_X1    g0792(.A(new_n721), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n709), .B(new_n969), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT111), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n778), .B2(new_n939), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n968), .A2(new_n996), .ZN(G387));
  NOR2_X1   g0797(.A1(new_n233), .A2(new_n715), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n998), .A2(new_n714), .B1(new_n663), .B2(new_n710), .ZN(new_n999));
  AOI21_X1  g0799(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n417), .A2(KEYINPUT50), .A3(new_n325), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT50), .B1(new_n417), .B2(new_n325), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n663), .B(new_n1000), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n999), .A2(new_n1003), .B1(new_n206), .B2(new_n660), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n709), .B1(new_n1004), .B2(new_n723), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G303), .A2(new_n793), .B1(new_n730), .B2(G311), .ZN(new_n1006));
  INV_X1    g0806(.A(G322), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n738), .C1(new_n754), .C2(new_n986), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT48), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n734), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n773), .A2(new_n1012), .B1(new_n727), .B2(G283), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT49), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n739), .A2(new_n284), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n254), .B(new_n1018), .C1(G326), .C2(new_n973), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n254), .B1(new_n742), .B2(new_n330), .C1(new_n202), .C2(new_n747), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n981), .B(new_n1021), .C1(G159), .C2(new_n766), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n730), .A2(new_n417), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n728), .A2(new_n419), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G77), .B2(new_n1012), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n755), .A2(G50), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1005), .B1(new_n1028), .B2(new_n721), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n652), .B2(new_n778), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n960), .B2(new_n967), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n961), .A2(new_n661), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n701), .A2(new_n960), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(G393));
  INV_X1    g0835(.A(KEYINPUT113), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n957), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n955), .A2(KEYINPUT113), .A3(new_n956), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n967), .A3(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n722), .B1(new_n205), .B2(new_n213), .C1(new_n243), .C2(new_n714), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n709), .A2(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n754), .A2(new_n743), .B1(new_n330), .B2(new_n738), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT51), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n728), .A2(new_n356), .B1(new_n734), .B2(new_n202), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n769), .A2(new_n325), .B1(new_n739), .B2(new_n735), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n254), .B1(new_n742), .B2(new_n795), .C1(new_n328), .C2(new_n747), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n754), .A2(new_n763), .B1(new_n986), .B2(new_n738), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT52), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n728), .A2(new_n284), .B1(new_n769), .B2(new_n760), .ZN(new_n1050));
  INV_X1    g0850(.A(G294), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n258), .B1(new_n742), .B2(new_n1007), .C1(new_n1051), .C2(new_n747), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n206), .A2(new_n739), .B1(new_n734), .B2(new_n786), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1043), .A2(new_n1047), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1041), .B1(new_n993), .B2(new_n1055), .C1(new_n930), .C2(new_n778), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1039), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n662), .B1(new_n957), .B2(new_n961), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(new_n964), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(G390));
  NAND4_X1  g0860(.A1(new_n682), .A2(new_n883), .A3(new_n811), .A4(G330), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n816), .A2(new_n809), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n883), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n911), .A2(new_n915), .B1(new_n1064), .B2(new_n913), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n909), .A2(new_n910), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n698), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n650), .B(new_n808), .C1(new_n696), .C2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n918), .B1(new_n1068), .B2(new_n809), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1066), .A2(new_n1069), .A3(new_n914), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1062), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n911), .A2(new_n915), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n809), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n629), .B2(new_n815), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n913), .B1(new_n1074), .B2(new_n918), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1068), .A2(new_n809), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n892), .B(new_n913), .C1(new_n1077), .C2(new_n918), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1078), .A3(new_n1061), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1071), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n502), .A2(new_n683), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n900), .A2(new_n637), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n682), .A2(new_n811), .A3(G330), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n918), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n1061), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1063), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1077), .A2(new_n1084), .A3(new_n1061), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1082), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1080), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1071), .A2(new_n1079), .A3(new_n1082), .A4(new_n1088), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n661), .A3(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1071), .A2(new_n1079), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1072), .A2(new_n718), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n709), .B1(new_n417), .B2(new_n784), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n755), .A2(G132), .B1(G128), .B2(new_n766), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT116), .Z(new_n1097));
  INV_X1    g0897(.A(G125), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n254), .B1(new_n742), .B2(new_n1098), .C1(new_n325), .C2(new_n739), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT115), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1012), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT53), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n734), .B2(new_n330), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1101), .A2(new_n1103), .B1(G159), .B2(new_n727), .ZN(new_n1104));
  INV_X1    g0904(.A(G137), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n769), .A2(new_n1105), .B1(new_n747), .B2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT114), .Z(new_n1108));
  NAND4_X1  g0908(.A1(new_n1097), .A2(new_n1100), .A3(new_n1104), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n258), .B1(new_n747), .B2(new_n205), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n769), .A2(new_n206), .B1(new_n786), .B2(new_n738), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(G77), .C2(new_n727), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n755), .A2(G116), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n739), .A2(new_n202), .B1(new_n742), .B2(new_n1051), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1116), .A2(KEYINPUT118), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n758), .A2(G87), .B1(KEYINPUT118), .B2(new_n1116), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1111), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1095), .B1(new_n1121), .B2(new_n721), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1093), .A2(new_n967), .B1(new_n1094), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1092), .A2(new_n1123), .ZN(G378));
  AND2_X1   g0924(.A1(new_n1091), .A2(new_n1082), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n916), .A2(new_n920), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1128), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n368), .A2(new_n369), .A3(new_n372), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n340), .A2(new_n847), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT119), .Z(new_n1134));
  XNOR2_X1  g0934(.A(new_n1132), .B(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n682), .A2(new_n883), .A3(new_n811), .A4(KEYINPUT40), .ZN(new_n1136));
  OAI21_X1  g0936(.A(G330), .B1(new_n1066), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n1137), .B2(new_n885), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n876), .A2(new_n884), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n835), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n834), .B1(new_n892), .B2(new_n893), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1134), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1132), .B(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1126), .A2(new_n1138), .A3(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1138), .A2(new_n1145), .B1(new_n916), .B2(new_n920), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT57), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n661), .B1(new_n1125), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1091), .A2(new_n1082), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1137), .A2(new_n1135), .A3(new_n885), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1144), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n921), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1126), .A2(new_n1138), .A3(new_n1145), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1149), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n967), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n254), .A2(G41), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n786), .B2(new_n742), .C1(new_n419), .C2(new_n747), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n971), .B(new_n1160), .C1(G77), .C2(new_n1012), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n769), .A2(new_n205), .B1(new_n284), .B2(new_n738), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G58), .B2(new_n767), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n206), .C2(new_n754), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT58), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G50), .B1(new_n251), .B2(new_n345), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1164), .A2(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1165), .B2(new_n1164), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n769), .A2(new_n800), .B1(new_n747), .B2(new_n1105), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n727), .A2(G150), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n734), .B2(new_n1106), .C1(new_n1098), .C2(new_n738), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G128), .C2(new_n755), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT59), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n973), .C2(G124), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n743), .B2(new_n739), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n721), .B1(new_n1169), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n707), .B1(new_n325), .B2(new_n783), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n1144), .C2(new_n719), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1158), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1157), .A2(new_n1184), .ZN(G375));
  AND2_X1   g0985(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n900), .A2(new_n637), .A3(new_n1081), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n947), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1089), .A3(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT120), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n759), .A2(new_n743), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G50), .A2(new_n727), .B1(new_n793), .B2(G150), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT121), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n766), .A2(G132), .B1(new_n973), .B2(G128), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n769), .B2(new_n1106), .C1(new_n754), .C2(new_n1105), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n254), .B1(new_n739), .B2(new_n201), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT122), .ZN(new_n1198));
  OR4_X1    g0998(.A1(new_n1192), .A2(new_n1194), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n769), .A2(new_n284), .B1(new_n1051), .B2(new_n738), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1024), .B(new_n1200), .C1(G77), .C2(new_n767), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n258), .B1(new_n742), .B2(new_n760), .C1(new_n206), .C2(new_n747), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n755), .B2(G283), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n205), .C2(new_n759), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n993), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n707), .B(new_n1205), .C1(new_n202), .C2(new_n783), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT123), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n719), .B2(new_n883), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1186), .B2(new_n966), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1191), .A2(new_n1209), .ZN(G381));
  OR2_X1    g1010(.A1(G393), .A2(G396), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(G384), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT124), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G381), .A2(G390), .A3(G378), .ZN(new_n1214));
  INV_X1    g1014(.A(G387), .ZN(new_n1215));
  INV_X1    g1015(.A(G375), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(G407));
  INV_X1    g1017(.A(G378), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n643), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G407), .B(G213), .C1(G375), .C2(new_n1219), .ZN(G409));
  NAND2_X1  g1020(.A1(new_n643), .A2(G213), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G378), .B(new_n1184), .C1(new_n1149), .C2(new_n1156), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n947), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT125), .B1(new_n1224), .B2(new_n1150), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(new_n1183), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1150), .A3(KEYINPUT125), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G378), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1221), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1209), .B1(new_n822), .B2(KEYINPUT126), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1188), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n661), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1231), .B1(new_n1188), .B2(new_n1089), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1230), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n822), .A2(KEYINPUT126), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1230), .B1(KEYINPUT126), .B2(new_n822), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n643), .A2(G213), .A3(G2897), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT61), .B1(new_n1229), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1222), .B1(new_n1244), .B2(G378), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1221), .A4(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1221), .B(new_n1247), .C1(new_n1223), .C2(new_n1228), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT62), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1243), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1211), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1059), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n964), .A2(new_n1058), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1211), .B(new_n1252), .C1(new_n1255), .C2(new_n1057), .ZN(new_n1256));
  AND4_X1   g1056(.A1(new_n968), .A2(new_n1254), .A3(new_n996), .A4(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1254), .A2(new_n1256), .B1(new_n968), .B2(new_n996), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1251), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1245), .A2(KEYINPUT63), .A3(new_n1221), .A4(new_n1247), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1249), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1259), .A2(new_n1243), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1261), .A2(new_n1265), .ZN(G405));
  INV_X1    g1066(.A(KEYINPUT127), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1247), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G375), .A2(new_n1218), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1222), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1222), .A3(new_n1268), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1260), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1270), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1259), .A3(new_n1271), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(G402));
endmodule


