//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1372, new_n1373, new_n1374;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  AND2_X1   g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n213), .A2(G20), .A3(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n211), .B(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT2), .B(G226), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XOR2_X1   g0033(.A(G107), .B(G116), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G351));
  AND2_X1   g0039(.A1(KEYINPUT3), .A2(G33), .ZN(new_n240));
  NOR2_X1   g0040(.A1(KEYINPUT3), .A2(G33), .ZN(new_n241));
  OAI211_X1 g0041(.A(G226), .B(G1698), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G1698), .ZN(new_n243));
  OAI211_X1 g0043(.A(G223), .B(new_n243), .C1(new_n240), .C2(new_n241), .ZN(new_n244));
  AND3_X1   g0044(.A1(KEYINPUT75), .A2(G33), .A3(G87), .ZN(new_n245));
  AOI21_X1  g0045(.A(KEYINPUT75), .B1(G33), .B2(G87), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n242), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(G33), .B2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G190), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n205), .A2(new_n255), .B1(new_n214), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(KEYINPUT64), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT64), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G45), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n260), .A3(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n257), .A2(G232), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n251), .A2(new_n252), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n261), .A2(new_n263), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n214), .A2(new_n256), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(new_n250), .B2(new_n248), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n265), .B1(new_n271), .B2(G200), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n249), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n240), .A2(new_n241), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT7), .B1(new_n276), .B2(new_n206), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G68), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G58), .ZN(new_n285));
  INV_X1    g0085(.A(G68), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G58), .A2(G68), .ZN(new_n288));
  OAI21_X1  g0088(.A(G20), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G159), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n289), .A2(KEYINPUT16), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n275), .B1(new_n284), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n280), .A2(new_n206), .A3(new_n281), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT7), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n286), .B1(new_n298), .B2(new_n282), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n289), .A2(new_n291), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT8), .B(G58), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n205), .B2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n305), .A2(new_n206), .A3(G1), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(new_n274), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n304), .A2(new_n307), .B1(new_n303), .B2(new_n306), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n272), .A2(new_n302), .A3(KEYINPUT77), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT17), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n308), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n293), .B2(new_n301), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n313), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n272), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n251), .A2(new_n316), .A3(new_n264), .ZN(new_n317));
  AOI21_X1  g0117(.A(G169), .B1(new_n251), .B2(new_n264), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n300), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n294), .B1(new_n284), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n289), .A2(KEYINPUT16), .A3(new_n291), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n274), .B1(new_n299), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n308), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT18), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT18), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n319), .A2(new_n324), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT18), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n315), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n305), .A2(G1), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT67), .B1(new_n335), .B2(G20), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AND4_X1   g0137(.A1(KEYINPUT67), .A2(new_n205), .A3(G13), .A4(G20), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT12), .B1(new_n340), .B2(G68), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT12), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n335), .A2(new_n342), .A3(G20), .A4(new_n286), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n286), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n279), .A2(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT66), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n206), .A2(G33), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT66), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n345), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n274), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n205), .A2(G20), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n340), .A2(G68), .A3(new_n275), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(KEYINPUT11), .A3(new_n274), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n344), .A2(new_n356), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n280), .A2(new_n281), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(G232), .A3(G1698), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(G226), .A3(new_n243), .ZN(new_n364));
  AND3_X1   g0164(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n250), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n257), .A2(G238), .B1(new_n261), .B2(new_n263), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n369), .B2(new_n370), .ZN(new_n373));
  OAI21_X1  g0173(.A(G200), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n369), .A2(new_n370), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(G190), .A3(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n361), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(G169), .B1(new_n372), .B2(new_n373), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(G179), .A3(new_n377), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT14), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(G169), .C1(new_n372), .C2(new_n373), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n379), .B1(new_n385), .B2(new_n360), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n334), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n362), .A2(G232), .A3(new_n243), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n362), .A2(G238), .A3(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n276), .A2(G107), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n250), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n257), .A2(G244), .B1(new_n261), .B2(new_n263), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G169), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n340), .A2(G77), .A3(new_n275), .A4(new_n357), .ZN(new_n397));
  INV_X1    g0197(.A(new_n290), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n303), .A2(new_n398), .B1(new_n206), .B2(new_n352), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT15), .B(G87), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n348), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n274), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n336), .A2(new_n338), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n352), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n392), .A2(new_n316), .A3(new_n393), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n396), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n394), .A2(new_n252), .ZN(new_n409));
  INV_X1    g0209(.A(G200), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n392), .B2(new_n393), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n405), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(KEYINPUT68), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT68), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n411), .B2(new_n405), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n408), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G226), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n267), .A2(new_n268), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n266), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n362), .A2(G222), .A3(new_n243), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n276), .A2(G77), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n362), .A2(G1698), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT65), .B(G223), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n420), .B(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n424), .B2(new_n250), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n316), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT8), .B(G58), .Z(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n350), .A3(new_n347), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n202), .A2(G20), .B1(G150), .B2(new_n290), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n275), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G50), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n205), .B2(G20), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n307), .A2(new_n432), .B1(new_n431), .B2(new_n306), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n426), .B1(G169), .B2(new_n425), .C1(new_n430), .C2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT69), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n434), .B2(new_n430), .ZN(new_n437));
  INV_X1    g0237(.A(G150), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n438), .A2(new_n398), .B1(new_n201), .B2(new_n206), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n347), .A2(new_n350), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n427), .ZN(new_n441));
  OAI211_X1 g0241(.A(KEYINPUT69), .B(new_n433), .C1(new_n441), .C2(new_n275), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(new_n442), .A3(KEYINPUT9), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT70), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n437), .A2(new_n442), .A3(KEYINPUT70), .A4(KEYINPUT9), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT71), .B1(new_n425), .B2(new_n410), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT10), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n425), .A2(KEYINPUT71), .A3(new_n410), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT9), .B1(new_n437), .B2(new_n442), .ZN(new_n453));
  INV_X1    g0253(.A(new_n425), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n252), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n447), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n425), .A2(new_n410), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n453), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n449), .B1(new_n459), .B2(new_n447), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n416), .B(new_n435), .C1(new_n457), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT72), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n447), .A2(new_n452), .A3(new_n456), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n459), .A2(new_n447), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(new_n449), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT72), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n435), .A4(new_n416), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n387), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n307), .B1(G1), .B2(new_n279), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n306), .A2(new_n471), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT25), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n206), .B(G87), .C1(new_n240), .C2(new_n241), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n362), .A2(new_n206), .A3(G87), .A4(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G116), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G20), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT23), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n206), .B2(G107), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n471), .A2(KEYINPUT23), .A3(G20), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT84), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT84), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n480), .A2(new_n481), .A3(new_n490), .A4(new_n487), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n489), .A2(KEYINPUT24), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(KEYINPUT84), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n274), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n492), .A2(KEYINPUT85), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n494), .A2(new_n274), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n489), .A2(KEYINPUT24), .A3(new_n491), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n475), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(G257), .B(G1698), .C1(new_n240), .C2(new_n241), .ZN(new_n502));
  OAI211_X1 g0302(.A(G250), .B(new_n243), .C1(new_n240), .C2(new_n241), .ZN(new_n503));
  INV_X1    g0303(.A(G294), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n502), .B(new_n503), .C1(new_n279), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n250), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n205), .A2(G45), .ZN(new_n507));
  OR2_X1    g0307(.A1(KEYINPUT5), .A2(G41), .ZN(new_n508));
  NAND2_X1  g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n250), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G264), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(G274), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G179), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n395), .B2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n501), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n505), .A2(new_n250), .B1(new_n511), .B2(G264), .ZN(new_n518));
  AOI21_X1  g0318(.A(G200), .B1(new_n518), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n506), .A2(new_n252), .A3(new_n512), .A4(new_n513), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n522), .B2(new_n519), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n475), .C1(new_n496), .C2(new_n500), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n254), .A2(G1), .ZN(new_n526));
  INV_X1    g0326(.A(new_n509), .ZN(new_n527));
  NOR2_X1   g0327(.A1(KEYINPUT5), .A2(G41), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G270), .A3(new_n267), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n530), .A2(new_n513), .ZN(new_n531));
  OAI211_X1 g0331(.A(G264), .B(G1698), .C1(new_n240), .C2(new_n241), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(new_n243), .C1(new_n240), .C2(new_n241), .ZN(new_n533));
  INV_X1    g0333(.A(G303), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n362), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n250), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n337), .A2(new_n339), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n205), .B2(G33), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n275), .B(new_n540), .C1(new_n336), .C2(new_n338), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n273), .A2(new_n249), .B1(G20), .B2(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  INV_X1    g0343(.A(G97), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n206), .C1(G33), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT20), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n542), .A2(KEYINPUT20), .A3(new_n545), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n539), .B(new_n541), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n537), .A2(new_n548), .A3(G169), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n548), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n531), .A2(new_n536), .A3(G190), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n530), .A2(new_n513), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n250), .B2(new_n535), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(new_n553), .C1(new_n555), .C2(new_n410), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(G179), .A3(new_n548), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n537), .A2(new_n548), .A3(KEYINPUT21), .A4(G169), .ZN(new_n558));
  AND4_X1   g0358(.A1(new_n551), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n400), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n340), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G87), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n470), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n346), .A2(G97), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n362), .A2(new_n206), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n286), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT19), .B1(new_n365), .B2(new_n366), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(new_n206), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  AOI211_X1 g0374(.A(new_n574), .B(new_n570), .C1(new_n571), .C2(new_n206), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n569), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n561), .B(new_n563), .C1(new_n576), .C2(new_n274), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT81), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n507), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n205), .A2(KEYINPUT81), .A3(G45), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n267), .A2(G250), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(G274), .B2(new_n526), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(G1698), .C1(new_n240), .C2(new_n241), .ZN(new_n584));
  OAI211_X1 g0384(.A(G238), .B(new_n243), .C1(new_n240), .C2(new_n241), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n482), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n250), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n583), .A2(new_n587), .A3(G190), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n410), .B1(new_n583), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n561), .ZN(new_n591));
  INV_X1    g0391(.A(new_n470), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n560), .ZN(new_n593));
  INV_X1    g0393(.A(new_n570), .ZN(new_n594));
  NAND2_X1  g0394(.A1(G33), .A2(G97), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT73), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n565), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n594), .B1(new_n599), .B2(G20), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n574), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n568), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n591), .B(new_n593), .C1(new_n603), .C2(new_n275), .ZN(new_n604));
  AOI21_X1  g0404(.A(G169), .B1(new_n583), .B2(new_n587), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n579), .A2(new_n580), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n267), .A2(G250), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n606), .A2(new_n607), .B1(new_n262), .B2(new_n507), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n250), .B2(new_n586), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n605), .B1(new_n316), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n577), .A2(new_n590), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n529), .A2(G257), .A3(new_n267), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n612), .A2(new_n513), .A3(KEYINPUT80), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT80), .B1(new_n612), .B2(new_n513), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G250), .B(G1698), .C1(new_n240), .C2(new_n241), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT79), .ZN(new_n617));
  OAI211_X1 g0417(.A(G244), .B(new_n243), .C1(new_n240), .C2(new_n241), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT4), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n362), .A2(KEYINPUT4), .A3(G244), .A4(new_n243), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n543), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n250), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n615), .A2(new_n623), .A3(new_n316), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n306), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n306), .A2(new_n544), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT78), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n625), .B(new_n628), .C1(new_n470), .C2(new_n544), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT6), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n631), .A2(new_n544), .A3(G107), .ZN(new_n632));
  XNOR2_X1  g0432(.A(G97), .B(G107), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  OAI22_X1  g0434(.A1(new_n634), .A2(new_n206), .B1(new_n352), .B2(new_n398), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n471), .B1(new_n298), .B2(new_n282), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n274), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n620), .A2(new_n621), .A3(new_n543), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT79), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n616), .B(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n267), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n612), .A2(new_n513), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT80), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n612), .A2(new_n513), .A3(KEYINPUT80), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n624), .B(new_n638), .C1(new_n648), .C2(G169), .ZN(new_n649));
  OAI21_X1  g0449(.A(G200), .B1(new_n642), .B2(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n633), .A2(new_n631), .ZN(new_n651));
  INV_X1    g0451(.A(new_n632), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n653), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n654));
  OAI21_X1  g0454(.A(G107), .B1(new_n277), .B2(new_n283), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n629), .B1(new_n656), .B2(new_n274), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n615), .A2(new_n623), .A3(G190), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n650), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n559), .A2(new_n611), .A3(new_n649), .A4(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n469), .A2(new_n525), .A3(new_n660), .ZN(G372));
  NOR2_X1   g0461(.A1(new_n329), .A2(new_n330), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n325), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n384), .A2(new_n382), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n376), .A2(new_n377), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n383), .B1(new_n665), .B2(G169), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n360), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n407), .B2(new_n379), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n663), .B1(new_n668), .B2(new_n315), .ZN(new_n669));
  INV_X1    g0469(.A(new_n465), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n435), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n558), .A2(new_n557), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n395), .B1(new_n531), .B2(new_n536), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT21), .B1(new_n673), .B2(new_n548), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n475), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT85), .B1(new_n492), .B2(new_n495), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n498), .A2(new_n497), .A3(new_n499), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n516), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n604), .A2(new_n610), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n561), .B1(new_n576), .B2(new_n274), .ZN(new_n683));
  INV_X1    g0483(.A(new_n563), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n590), .A3(new_n684), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n649), .A2(new_n659), .A3(new_n682), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n686), .A3(new_n524), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n682), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n649), .ZN(new_n690));
  INV_X1    g0490(.A(new_n649), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n611), .A2(new_n691), .A3(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n687), .A2(new_n693), .A3(new_n682), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n671), .B1(new_n468), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT87), .Z(G369));
  NOR2_X1   g0496(.A1(new_n679), .A2(new_n680), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n335), .A2(new_n206), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n703), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n679), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n525), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n705), .A2(new_n552), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n672), .B2(new_n674), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n556), .A2(new_n551), .A3(new_n557), .A4(new_n558), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT88), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT88), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n710), .B(new_n714), .C1(new_n711), .C2(new_n709), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n708), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n697), .A2(new_n705), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n675), .A2(new_n703), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n524), .B(new_n719), .C1(new_n679), .C2(new_n680), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n209), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n594), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n212), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n694), .A2(new_n729), .A3(new_n705), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n694), .B2(new_n705), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT90), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n705), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n506), .A2(new_n583), .A3(new_n587), .A4(new_n512), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n531), .A2(new_n536), .A3(G179), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n648), .A2(new_n739), .A3(KEYINPUT30), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n555), .A2(new_n609), .A3(G179), .A4(new_n518), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n615), .A2(new_n623), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n609), .A2(G179), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n744), .A2(new_n746), .A3(new_n514), .A4(new_n537), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT89), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n741), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT89), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n736), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n745), .A2(new_n740), .A3(new_n747), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n753), .B2(new_n703), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n733), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(KEYINPUT30), .B1(new_n648), .B2(new_n739), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n583), .A2(new_n587), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n514), .A2(new_n537), .A3(new_n316), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n648), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n749), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n740), .A3(new_n751), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n735), .ZN(new_n762));
  INV_X1    g0562(.A(new_n754), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(KEYINPUT90), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n649), .A2(new_n659), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n765), .A2(new_n689), .A3(new_n711), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n766), .A2(new_n524), .A3(new_n517), .A4(new_n705), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n755), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G330), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n732), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n728), .B1(new_n771), .B2(G1), .ZN(G364));
  INV_X1    g0572(.A(new_n716), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n305), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n205), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n723), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n713), .A2(new_n708), .A3(new_n715), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n209), .A2(new_n362), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(G116), .B2(new_n209), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n722), .A2(new_n362), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n258), .A2(new_n260), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n213), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n238), .A2(new_n254), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n249), .B1(G20), .B2(new_n395), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n777), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n206), .A2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n252), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n252), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n316), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n504), .B1(new_n805), .B2(new_n534), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n206), .A2(new_n316), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n252), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n800), .B(new_n806), .C1(G326), .C2(new_n809), .ZN(new_n810));
  AND3_X1   g0610(.A1(new_n807), .A2(KEYINPUT91), .A3(new_n801), .ZN(new_n811));
  AOI21_X1  g0611(.A(KEYINPUT91), .B1(new_n807), .B2(new_n801), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G322), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT92), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n808), .A2(G190), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(KEYINPUT92), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G190), .A2(G200), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n807), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n276), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n797), .A2(new_n821), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n824), .B1(G329), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n810), .A2(new_n815), .A3(new_n820), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n818), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n829), .A2(new_n286), .B1(new_n798), .B2(new_n471), .ZN(new_n830));
  INV_X1    g0630(.A(new_n809), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n826), .A2(G159), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n431), .B1(new_n832), .B2(KEYINPUT32), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n814), .A2(G58), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n362), .B1(new_n822), .B2(new_n352), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(KEYINPUT32), .B2(new_n832), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n805), .A2(new_n562), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G97), .B2(new_n803), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n828), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n796), .B1(new_n841), .B2(new_n793), .ZN(new_n842));
  INV_X1    g0642(.A(new_n792), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n712), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n780), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  OAI22_X1  g0646(.A1(new_n829), .A2(new_n799), .B1(new_n805), .B2(new_n471), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G303), .B2(new_n809), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n814), .A2(G294), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n276), .B1(new_n822), .B2(new_n538), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G311), .B2(new_n826), .ZN(new_n851));
  INV_X1    g0651(.A(new_n798), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(G87), .B1(new_n803), .B2(G97), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n848), .A2(new_n849), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n822), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n809), .A2(G137), .B1(new_n855), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G143), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n438), .B2(new_n829), .C1(new_n857), .C2(new_n813), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT34), .Z(new_n859));
  NOR2_X1   g0659(.A1(new_n804), .A2(new_n285), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n362), .B1(new_n825), .B2(new_n861), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n431), .A2(new_n805), .B1(new_n798), .B2(new_n286), .ZN(new_n863));
  OR3_X1    g0663(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n854), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n793), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n793), .A2(new_n790), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n778), .B1(new_n352), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n407), .A2(new_n703), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n405), .A2(new_n703), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n413), .B2(new_n415), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n873), .B2(new_n408), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n869), .B1(new_n790), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n416), .A2(new_n705), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n694), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n874), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n694), .B2(new_n705), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n769), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n777), .B1(new_n880), .B2(new_n769), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G384));
  OR2_X1    g0685(.A1(new_n653), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n653), .A2(KEYINPUT35), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n249), .A2(new_n206), .A3(new_n538), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT93), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(KEYINPUT36), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(KEYINPUT36), .ZN(new_n893));
  OAI21_X1  g0693(.A(G77), .B1(new_n285), .B2(new_n286), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n894), .A2(new_n212), .B1(G50), .B2(new_n286), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(G1), .A3(new_n305), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT94), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n892), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT95), .Z(new_n899));
  INV_X1    g0699(.A(new_n701), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n324), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n313), .A2(new_n272), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n329), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT97), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT37), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n903), .B2(KEYINPUT37), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n329), .A2(new_n901), .A3(new_n902), .A4(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT96), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n901), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n907), .A2(new_n911), .B1(new_n333), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n909), .A2(new_n910), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n905), .B2(new_n906), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n913), .A2(KEYINPUT98), .A3(KEYINPUT38), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n333), .A2(new_n912), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT97), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT37), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n911), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n917), .A2(KEYINPUT38), .A3(new_n915), .A4(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT98), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n915), .A3(new_n921), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n916), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n763), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n767), .ZN(new_n932));
  INV_X1    g0732(.A(new_n379), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n360), .A2(new_n703), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n667), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n360), .B(new_n703), .C1(new_n385), .C2(new_n379), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n874), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n928), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n311), .A2(new_n314), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n912), .B1(new_n663), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n918), .A2(KEYINPUT100), .A3(new_n909), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT100), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n903), .A2(new_n946), .A3(KEYINPUT37), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n922), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n932), .A2(KEYINPUT40), .A3(new_n937), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n942), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n468), .A2(new_n932), .ZN(new_n955));
  OAI21_X1  g0755(.A(G330), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n954), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n935), .A2(new_n936), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n694), .A2(new_n876), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(new_n871), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n928), .A2(new_n961), .B1(new_n663), .B2(new_n701), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n916), .A2(new_n924), .A3(KEYINPUT39), .A4(new_n927), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n385), .A2(new_n360), .A3(new_n705), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n951), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n468), .B1(new_n730), .B2(new_n731), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT101), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT101), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n468), .B(new_n972), .C1(new_n730), .C2(new_n731), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n671), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n969), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n957), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n957), .A2(new_n975), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT103), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n976), .B1(new_n205), .B2(new_n774), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n977), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(KEYINPUT103), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n899), .B1(new_n979), .B2(new_n981), .ZN(G367));
  OAI221_X1 g0782(.A(new_n794), .B1(new_n209), .B2(new_n400), .C1(new_n785), .C2(new_n231), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(new_n777), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n577), .A2(new_n705), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(new_n682), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n611), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n362), .B1(new_n822), .B2(new_n431), .ZN(new_n990));
  INV_X1    g0790(.A(G159), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n829), .A2(new_n991), .B1(new_n798), .B2(new_n352), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(G137), .C2(new_n826), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n831), .A2(new_n857), .B1(new_n804), .B2(new_n286), .ZN(new_n994));
  INV_X1    g0794(.A(new_n805), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(G58), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n993), .B(new_n996), .C1(new_n438), .C2(new_n813), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n852), .A2(G97), .B1(new_n803), .B2(G107), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT111), .B(G311), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n998), .B1(new_n829), .B2(new_n504), .C1(new_n831), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n276), .B1(new_n825), .B2(new_n1001), .C1(new_n799), .C2(new_n822), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT46), .B1(new_n995), .B2(G116), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n995), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n534), .C2(new_n813), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n997), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT47), .Z(new_n1008));
  INV_X1    g0808(.A(new_n793), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n984), .B1(new_n989), .B2(new_n843), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n723), .B(KEYINPUT41), .Z(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n720), .A2(new_n718), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT104), .B1(new_n649), .B2(new_n705), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n657), .B1(new_n395), .B2(new_n744), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT104), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n624), .A4(new_n703), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n649), .B(new_n659), .C1(new_n657), .C2(new_n705), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT44), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1013), .A2(new_n1020), .A3(KEYINPUT44), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(new_n718), .A3(new_n720), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1025), .A2(new_n720), .A3(KEYINPUT45), .A4(new_n718), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1023), .A2(new_n1024), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n717), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n720), .B1(new_n707), .B2(new_n719), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(new_n716), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1031), .A2(new_n1033), .A3(new_n732), .A4(new_n769), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT108), .B1(new_n707), .B2(new_n716), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n707), .A2(new_n716), .A3(KEYINPUT108), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1030), .A2(KEYINPUT107), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1029), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1013), .A2(new_n1020), .A3(KEYINPUT44), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT44), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1038), .A2(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT107), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT109), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1036), .A2(new_n1035), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT109), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1030), .A2(KEYINPUT107), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1034), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1012), .B1(new_n1051), .B2(new_n770), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT110), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT110), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n1012), .C1(new_n1051), .C2(new_n770), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n776), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT42), .B1(new_n1020), .B2(new_n720), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1013), .A2(new_n1058), .A3(new_n1025), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n649), .C2(new_n703), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT105), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1060), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n707), .A2(new_n716), .A3(new_n1025), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1067), .A2(new_n1068), .B1(KEYINPUT106), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(KEYINPUT106), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1010), .B1(new_n1056), .B2(new_n1072), .ZN(G387));
  OAI22_X1  g0873(.A1(new_n781), .A2(new_n725), .B1(G107), .B2(new_n209), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n228), .A2(new_n786), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n725), .ZN(new_n1076));
  AOI211_X1 g0876(.A(G45), .B(new_n1076), .C1(G68), .C2(G77), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n303), .A2(G50), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT50), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n785), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1074), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT112), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n794), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n777), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT113), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n276), .B1(new_n826), .B2(G150), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n352), .B2(new_n805), .C1(new_n544), .C2(new_n798), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT114), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n809), .A2(G159), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT115), .Z(new_n1091));
  AOI22_X1  g0891(.A1(new_n818), .A2(new_n427), .B1(new_n855), .B2(G68), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n400), .B2(new_n804), .C1(new_n813), .C2(new_n431), .ZN(new_n1093));
  OR3_X1    g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n362), .B1(new_n826), .B2(G326), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n804), .A2(new_n799), .B1(new_n805), .B2(new_n504), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT116), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n809), .A2(G322), .B1(new_n855), .B2(G303), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n829), .B2(new_n999), .C1(new_n1001), .C2(new_n813), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT48), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT49), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1095), .B1(new_n538), .B2(new_n798), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1094), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1086), .B1(new_n793), .B2(new_n1106), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n707), .A2(new_n843), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n776), .A2(new_n1033), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n771), .A2(new_n1033), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(KEYINPUT117), .A3(new_n723), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n771), .B2(new_n1033), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT117), .B1(new_n1110), .B2(new_n723), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(G393));
  XNOR2_X1  g0914(.A(new_n1030), .B(new_n717), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n775), .B1(new_n1115), .B2(KEYINPUT118), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(KEYINPUT118), .B2(new_n1115), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n814), .A2(G159), .B1(G150), .B2(new_n809), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT51), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n362), .B1(new_n825), .B2(new_n857), .C1(new_n303), .C2(new_n822), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n829), .A2(new_n431), .B1(new_n798), .B2(new_n562), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n804), .A2(new_n352), .B1(new_n805), .B2(new_n286), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n823), .A2(new_n813), .B1(new_n831), .B2(new_n1001), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT119), .B(KEYINPUT52), .Z(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n829), .A2(new_n534), .B1(new_n805), .B2(new_n799), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n804), .A2(new_n538), .B1(new_n798), .B2(new_n471), .ZN(new_n1130));
  INV_X1    g0930(.A(G322), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n276), .B1(new_n825), .B2(new_n1131), .C1(new_n504), .C2(new_n822), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1127), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n793), .B1(new_n1123), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n784), .A2(new_n235), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n795), .B1(G97), .B2(new_n722), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n778), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1135), .B(new_n1138), .C1(new_n1025), .C2(new_n843), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n723), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1117), .B(new_n1139), .C1(new_n1051), .C2(new_n1141), .ZN(G390));
  NAND2_X1  g0942(.A1(new_n951), .A2(new_n964), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT120), .B1(new_n935), .B2(new_n936), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT120), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n960), .A2(new_n871), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n963), .A2(new_n967), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n961), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n964), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1148), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n525), .A2(new_n660), .A3(new_n703), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n937), .B(G330), .C1(new_n1153), .C2(new_n930), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT121), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n768), .A2(G330), .A3(new_n878), .A4(new_n958), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT121), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1154), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n963), .A2(new_n967), .B1(new_n1150), .B2(new_n964), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1159), .C1(new_n1160), .C2(new_n1148), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n1157), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n775), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1149), .A2(new_n790), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n778), .B1(new_n303), .B2(new_n867), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n804), .A2(new_n352), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n831), .A2(new_n799), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G107), .C2(new_n818), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n276), .B1(new_n825), .B2(new_n504), .C1(new_n544), .C2(new_n822), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n838), .B(new_n1169), .C1(G68), .C2(new_n852), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n538), .C2(new_n813), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT123), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n276), .B1(new_n826), .B2(G125), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n822), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n814), .B2(G132), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n818), .A2(G137), .B1(new_n852), .B2(G50), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n804), .A2(new_n991), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G128), .B2(new_n809), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n805), .A2(new_n438), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT53), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1173), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1164), .B(new_n1165), .C1(new_n1009), .C2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1163), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n960), .A2(new_n871), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1146), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n1144), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G330), .B(new_n878), .C1(new_n1153), .C2(new_n930), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1156), .A2(new_n1190), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n754), .B1(new_n761), .B2(new_n735), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n767), .B1(new_n1196), .B2(KEYINPUT90), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n752), .A2(new_n733), .A3(new_n754), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G330), .B(new_n878), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1159), .B1(new_n1199), .B2(new_n959), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1195), .B1(new_n1200), .B2(new_n1190), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n468), .A2(G330), .A3(new_n932), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n974), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1203), .A2(new_n1155), .A3(new_n1157), .A4(new_n1161), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT122), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n723), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n974), .A2(new_n1202), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1201), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1162), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1205), .B1(new_n1204), .B2(new_n723), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1188), .B1(new_n1210), .B2(new_n1211), .ZN(G378));
  NAND2_X1  g1012(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n969), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n465), .A2(new_n435), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n437), .A2(new_n442), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n900), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n465), .A2(new_n435), .A3(new_n1218), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1221), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1220), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(G330), .B1(new_n952), .B2(new_n953), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n942), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n940), .B1(new_n928), .B2(new_n938), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1228), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1215), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n942), .A2(new_n1229), .A3(new_n1227), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1232), .B1(new_n1231), .B2(new_n1228), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n969), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1214), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT124), .B1(new_n1239), .B2(new_n1215), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1213), .B(KEYINPUT57), .C1(new_n1238), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n723), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(G33), .A2(G41), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G50), .B(new_n1246), .C1(new_n276), .C2(new_n253), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n804), .A2(new_n286), .B1(new_n805), .B2(new_n352), .ZN(new_n1248));
  AOI211_X1 g1048(.A(G41), .B(new_n362), .C1(new_n826), .C2(G283), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n400), .B2(new_n822), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(G107), .C2(new_n814), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G97), .A2(new_n818), .B1(new_n809), .B2(G116), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n285), .C2(new_n798), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT58), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1247), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1254), .B2(new_n1253), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n855), .A2(G137), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n829), .B2(new_n861), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n814), .B2(G128), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n809), .A2(G125), .B1(new_n803), .B2(G150), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(new_n805), .C2(new_n1175), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1261), .A2(KEYINPUT59), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(KEYINPUT59), .ZN(new_n1263));
  INV_X1    g1063(.A(G124), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1246), .B1(new_n825), .B2(new_n1264), .C1(new_n991), .C2(new_n798), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n793), .B1(new_n1256), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n778), .B1(new_n431), .B2(new_n867), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(new_n1232), .C2(new_n791), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1243), .B2(new_n776), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1245), .A2(new_n1271), .ZN(G375));
  INV_X1    g1072(.A(new_n1207), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1201), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1012), .A3(new_n1208), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1192), .A2(new_n790), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n829), .A2(new_n538), .B1(new_n805), .B2(new_n544), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G294), .B2(new_n809), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n814), .A2(G283), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n276), .B1(new_n822), .B2(new_n471), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G303), .B2(new_n826), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G77), .A2(new_n852), .B1(new_n803), .B2(new_n560), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1279), .A2(new_n1280), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n831), .A2(new_n861), .B1(new_n805), .B2(new_n991), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(G50), .B2(new_n803), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n814), .A2(G137), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n822), .A2(new_n438), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n276), .B(new_n1288), .C1(G128), .C2(new_n826), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1175), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n818), .A2(new_n1290), .B1(new_n852), .B2(G58), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1009), .B1(new_n1284), .B2(new_n1292), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n778), .B(new_n1293), .C1(new_n286), .C2(new_n867), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(KEYINPUT125), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1201), .A2(new_n776), .B1(new_n1277), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1276), .A2(new_n1296), .ZN(G381));
  OAI211_X1 g1097(.A(new_n845), .B(new_n1109), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1298));
  INV_X1    g1098(.A(G390), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n884), .ZN(new_n1300));
  OR4_X1    g1100(.A1(G387), .A2(G381), .A3(new_n1298), .A4(new_n1300), .ZN(new_n1301));
  OR3_X1    g1101(.A1(new_n1301), .A2(G375), .A3(G378), .ZN(G407));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n702), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G407), .B(G213), .C1(G375), .C2(new_n1304), .ZN(G409));
  NAND2_X1  g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1306), .A2(new_n1307), .A3(new_n1298), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1306), .B2(new_n1298), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1034), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1037), .A2(new_n1044), .A3(KEYINPUT109), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1048), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1311), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n771), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1054), .B1(new_n1315), .B2(new_n1012), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1055), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n775), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1072), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G390), .B1(new_n1320), .B2(new_n1010), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1010), .B(G390), .C1(new_n1056), .C2(new_n1072), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1310), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G387), .A2(new_n1299), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1326), .A3(new_n1322), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n702), .A2(G213), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G378), .B(new_n1271), .C1(new_n1242), .C2(new_n1244), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1213), .A2(new_n1012), .A3(new_n1243), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n776), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1269), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1334), .B(new_n1188), .C1(new_n1211), .C2(new_n1210), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1330), .B1(new_n1331), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1330), .A2(G2897), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1208), .A2(KEYINPUT60), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1275), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1273), .A2(KEYINPUT60), .A3(new_n1274), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n723), .A3(new_n1341), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1342), .A2(G384), .A3(new_n1296), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G384), .B1(new_n1342), .B2(new_n1296), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1338), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1296), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n884), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1342), .A2(G384), .A3(new_n1296), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1347), .A2(new_n1348), .A3(new_n1337), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1345), .A2(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1329), .B1(new_n1336), .B2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT62), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1352), .B1(new_n1336), .B2(new_n1353), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1351), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1336), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1328), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1328), .B(new_n1329), .C1(new_n1336), .C2(new_n1350), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT63), .B1(new_n1336), .B2(new_n1353), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1336), .A2(KEYINPUT63), .A3(new_n1353), .ZN(new_n1360));
  NOR3_X1   g1160(.A1(new_n1358), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(KEYINPUT127), .B1(new_n1357), .B2(new_n1361), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1360), .A2(new_n1359), .ZN(new_n1363));
  AND2_X1   g1163(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1351), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT127), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1356), .ZN(new_n1368));
  NOR3_X1   g1168(.A1(new_n1368), .A2(new_n1351), .A3(new_n1354), .ZN(new_n1369));
  OAI211_X1 g1169(.A(new_n1366), .B(new_n1367), .C1(new_n1369), .C2(new_n1328), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1362), .A2(new_n1370), .ZN(G405));
  NAND2_X1  g1171(.A1(G375), .A2(new_n1303), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1372), .A2(new_n1331), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1373), .B(new_n1353), .ZN(new_n1374));
  XNOR2_X1  g1174(.A(new_n1374), .B(new_n1364), .ZN(G402));
endmodule


