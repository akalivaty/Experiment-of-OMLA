//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n209), .A2(KEYINPUT0), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n215), .B1(KEYINPUT0), .B2(new_n209), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n217), .A2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n202), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n238), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n248), .B(KEYINPUT67), .Z(new_n249));
  NAND3_X1  g0049(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  AND3_X1   g0051(.A1(new_n250), .A2(new_n210), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n250), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n249), .A2(new_n252), .B1(new_n202), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n203), .A2(G20), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n211), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR4_X1   g0064(.A1(new_n256), .A2(new_n257), .A3(new_n260), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n251), .A2(new_n210), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n254), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n271), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G222), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(G1698), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  AND2_X1   g0083(.A1(G1), .A2(G13), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(new_n270), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G41), .A2(G45), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n290), .A2(new_n210), .B1(new_n291), .B2(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT65), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n271), .A2(new_n294), .A3(new_n286), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n289), .B1(new_n296), .B2(G226), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G190), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT68), .A2(KEYINPUT10), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n269), .A2(new_n298), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT68), .A2(KEYINPUT10), .ZN(new_n303));
  XOR2_X1   g0103(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n280), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G226), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G1698), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n273), .A2(new_n306), .A3(new_n275), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n271), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n292), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(G232), .B1(new_n285), .B2(new_n287), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT74), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n288), .B1(new_n228), .B2(new_n292), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n311), .ZN(new_n318));
  AOI21_X1  g0118(.A(G200), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n317), .A2(new_n311), .A3(G190), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT3), .B(G33), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT7), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n322), .A2(new_n323), .A3(G20), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT7), .B1(new_n276), .B2(new_n211), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT71), .ZN(new_n328));
  AND2_X1   g0128(.A1(G58), .A2(G68), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(G20), .C1(new_n329), .C2(new_n201), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n261), .A2(G159), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(G58), .B(G68), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n333), .B2(G20), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n327), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n329), .B2(new_n201), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT71), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(KEYINPUT72), .A3(new_n331), .A4(new_n330), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n326), .A2(new_n335), .A3(KEYINPUT16), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT16), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n274), .B2(G33), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n272), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n275), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n323), .A2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n323), .B1(new_n322), .B2(G20), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n240), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n337), .A2(new_n331), .A3(new_n330), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n340), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n339), .A2(new_n350), .A3(new_n266), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n258), .B1(new_n246), .B2(G20), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n252), .B1(new_n253), .B2(new_n258), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n321), .A2(KEYINPUT17), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n351), .B(new_n353), .C1(new_n319), .C2(new_n320), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT17), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n351), .A2(new_n353), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n317), .A2(new_n311), .A3(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n315), .A2(new_n318), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT18), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n359), .A2(KEYINPUT18), .A3(new_n363), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(KEYINPUT75), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(KEYINPUT18), .A3(new_n363), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n358), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n297), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n268), .C1(G169), .C2(new_n297), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n322), .A2(G232), .A3(new_n305), .ZN(new_n374));
  INV_X1    g0174(.A(G107), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n322), .A2(G1698), .ZN(new_n376));
  INV_X1    g0176(.A(G238), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n374), .B1(new_n375), .B2(new_n322), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n271), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n296), .A2(G244), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n288), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n362), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G20), .A2(G77), .ZN(new_n384));
  INV_X1    g0184(.A(G87), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT15), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT15), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G87), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n384), .B1(new_n258), .B2(new_n262), .C1(new_n390), .C2(new_n259), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n266), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n252), .A2(G77), .A3(new_n247), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(G77), .C2(new_n250), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n383), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n382), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n371), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n382), .A2(G200), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n394), .B1(new_n396), .B2(G190), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n304), .A2(new_n370), .A3(new_n373), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n228), .A2(G1698), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G226), .B2(G1698), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n404), .B1(new_n406), .B2(new_n276), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n379), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n377), .B1(new_n293), .B2(new_n295), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT69), .ZN(new_n410));
  INV_X1    g0210(.A(new_n288), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n271), .A2(new_n294), .A3(new_n286), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n294), .B1(new_n271), .B2(new_n286), .ZN(new_n414));
  OAI21_X1  g0214(.A(G238), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT69), .B1(new_n415), .B2(new_n288), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n408), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(KEYINPUT69), .A3(new_n288), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT13), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n408), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n418), .A2(KEYINPUT70), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n421), .A2(new_n425), .A3(new_n422), .A4(new_n408), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(G169), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n424), .A2(new_n429), .A3(new_n426), .A4(G169), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n418), .A2(G179), .A3(new_n423), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n253), .A2(new_n240), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT12), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n240), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n277), .B2(new_n259), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(KEYINPUT11), .A3(new_n266), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n252), .A2(G68), .A3(new_n247), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT11), .B1(new_n436), .B2(new_n266), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n432), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n424), .A2(G200), .A3(new_n426), .ZN(new_n443));
  INV_X1    g0243(.A(G190), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n417), .B2(KEYINPUT13), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n441), .B1(new_n445), .B2(new_n423), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n403), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT82), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n322), .A2(G264), .A3(G1698), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n322), .A2(G257), .A3(new_n305), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(new_n322), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n379), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT81), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT81), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n457), .A3(new_n379), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n246), .A2(G45), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT77), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G41), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n379), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n456), .A2(new_n458), .B1(G270), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n463), .A2(new_n285), .A3(new_n467), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  INV_X1    g0271(.A(G97), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n211), .C1(G33), .C2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(new_n266), .C1(new_n211), .C2(G116), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n250), .A2(G116), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n246), .A2(G33), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n250), .A2(new_n478), .A3(new_n210), .A4(new_n251), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n480), .B2(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n469), .A2(G179), .A3(new_n470), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n468), .A2(G270), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n454), .A2(new_n457), .A3(new_n379), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n457), .B1(new_n454), .B2(new_n379), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n470), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n362), .B1(new_n476), .B2(new_n481), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n483), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n469), .A2(G190), .A3(new_n470), .ZN(new_n493));
  INV_X1    g0293(.A(new_n482), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n487), .A2(G200), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n450), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n487), .A2(new_n494), .A3(new_n371), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n487), .A2(new_n489), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT21), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n273), .A2(new_n275), .A3(new_n211), .A4(G87), .ZN(new_n506));
  XOR2_X1   g0306(.A(KEYINPUT83), .B(KEYINPUT22), .Z(new_n507));
  XNOR2_X1  g0307(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(new_n375), .A3(G20), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT84), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n510), .A2(new_n512), .A3(new_n513), .A4(KEYINPUT84), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n508), .A2(new_n509), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n509), .B1(new_n508), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n266), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n253), .A2(new_n375), .ZN(new_n522));
  NOR2_X1   g0322(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n524), .A2(new_n526), .B1(new_n480), .B2(G107), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT77), .B1(new_n460), .B2(G41), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n461), .ZN(new_n530));
  INV_X1    g0330(.A(G45), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G1), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n466), .B2(KEYINPUT77), .ZN(new_n533));
  OAI211_X1 g0333(.A(G264), .B(new_n271), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n534), .A2(new_n470), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n273), .A2(new_n275), .A3(G257), .A4(G1698), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n273), .A2(new_n275), .A3(G250), .A4(new_n305), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G294), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n379), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n362), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n541), .A2(KEYINPUT86), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n535), .A2(new_n540), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n541), .A2(KEYINPUT86), .B1(new_n543), .B2(new_n371), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n528), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n535), .A2(G190), .A3(new_n540), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n543), .A2(G200), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n521), .A2(new_n527), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n530), .A2(new_n533), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n468), .A2(G257), .B1(new_n550), .B2(new_n285), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n273), .A2(new_n275), .A3(G250), .A4(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(new_n305), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n471), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n379), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  AND2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g0363(.A1(KEYINPUT6), .A2(G97), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(G107), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n375), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G20), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n261), .A2(G77), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n375), .B1(new_n346), .B2(new_n347), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n266), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n250), .A2(G97), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n480), .B2(G97), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n558), .A2(new_n371), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n551), .A2(new_n557), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n362), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n551), .A2(new_n557), .A3(new_n444), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n558), .B2(G200), .ZN(new_n579));
  INV_X1    g0379(.A(new_n574), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n346), .A2(new_n347), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n569), .B(new_n568), .C1(new_n581), .C2(new_n375), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n580), .B1(new_n582), .B2(new_n266), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n575), .A2(new_n577), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n273), .A2(new_n275), .A3(G238), .A4(new_n305), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n379), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n271), .A2(G274), .A3(new_n532), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n459), .B(G250), .C1(new_n290), .C2(new_n210), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT78), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT78), .B1(new_n591), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n590), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n362), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n591), .A2(new_n592), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT78), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n593), .B1(new_n379), .B2(new_n589), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n371), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n389), .A2(new_n250), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n211), .B1(new_n404), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n561), .A2(new_n385), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n273), .A2(new_n275), .A3(new_n211), .A4(G68), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n604), .B1(new_n259), .B2(new_n472), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n603), .B1(new_n610), .B2(new_n266), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n480), .A2(new_n389), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(KEYINPUT79), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT79), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n611), .B2(new_n612), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n597), .B(new_n602), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n601), .A2(G190), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n596), .A2(G200), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT80), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n252), .A2(new_n620), .A3(G87), .A4(new_n478), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT80), .B1(new_n479), .B2(new_n385), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n549), .A2(new_n585), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n449), .A2(new_n505), .A3(new_n627), .ZN(G372));
  NAND2_X1  g0428(.A1(new_n447), .A2(new_n399), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n358), .B1(new_n442), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n359), .A2(new_n363), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT18), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n367), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n304), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n373), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n596), .A2(new_n444), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n619), .A2(new_n624), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n619), .A2(KEYINPUT87), .A3(new_n624), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n613), .B(KEYINPUT79), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n602), .A2(new_n597), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n548), .A4(new_n584), .ZN(new_n647));
  INV_X1    g0447(.A(new_n578), .ZN(new_n648));
  AOI21_X1  g0448(.A(G200), .B1(new_n551), .B2(new_n557), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n583), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n572), .A2(new_n574), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n551), .A2(new_n557), .A3(new_n371), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n577), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n548), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n600), .A2(new_n593), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n299), .B1(new_n655), .B2(new_n590), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n611), .A2(new_n623), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n640), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n642), .A3(new_n618), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n617), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT88), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n545), .B(new_n483), .C1(new_n491), .C2(new_n490), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n647), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n626), .B2(new_n653), .ZN(new_n664));
  INV_X1    g0464(.A(new_n653), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n659), .A3(new_n666), .A4(new_n617), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n664), .A2(new_n617), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n449), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n637), .A2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n246), .A2(new_n211), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n545), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n528), .A2(new_n678), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n545), .A2(new_n548), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n494), .A2(new_n679), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n505), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT89), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n502), .A2(new_n686), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n685), .B1(new_n497), .B2(new_n504), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT89), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  AOI211_X1 g0493(.A(new_n672), .B(new_n684), .C1(new_n691), .C2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n502), .B2(new_n678), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n492), .A2(KEYINPUT90), .A3(new_n679), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n682), .B2(new_n680), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n545), .A2(new_n678), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n695), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n207), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT91), .B1(new_n703), .B2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n703), .A2(KEYINPUT91), .A3(G41), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n606), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n213), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n505), .A2(new_n627), .A3(new_n679), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n543), .A2(new_n371), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n576), .A2(new_n596), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n469), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n469), .A2(new_n714), .A3(new_n715), .A4(KEYINPUT30), .ZN(new_n719));
  AOI21_X1  g0519(.A(G179), .B1(new_n535), .B2(new_n540), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n487), .A2(new_n576), .A3(new_n596), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n722), .B2(new_n678), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n672), .B1(new_n713), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g0526(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n727));
  INV_X1    g0527(.A(new_n669), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(new_n678), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n660), .B(new_n654), .C1(new_n502), .C2(new_n545), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT26), .B1(new_n660), .B2(new_n653), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n665), .A2(new_n625), .A3(new_n617), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n617), .C1(KEYINPUT26), .C2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT29), .B(new_n679), .C1(new_n730), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n726), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n712), .B1(new_n735), .B2(G1), .ZN(G364));
  INV_X1    g0536(.A(G13), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n246), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n707), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n322), .A2(G355), .A3(new_n207), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n244), .A2(new_n531), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n703), .A2(new_n322), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G45), .B2(new_n213), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n743), .B1(G116), .B2(new_n207), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n210), .B1(G20), .B2(new_n362), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n742), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n211), .A2(new_n444), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n299), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n276), .B1(new_n756), .B2(new_n453), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n371), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n211), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G322), .A2(new_n760), .B1(new_n764), .B2(G329), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n761), .A2(new_n755), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n758), .A2(new_n761), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n765), .B1(new_n766), .B2(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n757), .B(new_n770), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n211), .B1(new_n762), .B2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(new_n444), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n776), .A2(G294), .B1(G326), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT95), .ZN(new_n779));
  INV_X1    g0579(.A(new_n769), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G58), .A2(new_n760), .B1(new_n780), .B2(G77), .ZN(new_n781));
  INV_X1    g0581(.A(new_n777), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n202), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n763), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n787));
  XNOR2_X1  g0587(.A(new_n786), .B(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n322), .B1(new_n767), .B2(new_n375), .C1(new_n385), .C2(new_n756), .ZN(new_n789));
  INV_X1    g0589(.A(new_n772), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n790), .A2(new_n240), .B1(new_n775), .B2(new_n472), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n774), .A2(new_n779), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n751), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n753), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n692), .A2(new_n689), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n750), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n672), .B1(new_n691), .B2(new_n693), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n741), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n691), .A2(new_n672), .A3(new_n693), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  NAND3_X1  g0602(.A1(new_n395), .A2(new_n397), .A3(new_n679), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n401), .A2(new_n400), .B1(new_n394), .B2(new_n678), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n399), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n678), .B(new_n805), .C1(new_n663), .C2(new_n668), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(KEYINPUT98), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n669), .B2(new_n679), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT99), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  INV_X1    g0611(.A(new_n726), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT100), .Z(new_n814));
  AOI21_X1  g0614(.A(new_n741), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n767), .A2(new_n240), .B1(new_n763), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n756), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n276), .B1(new_n819), .B2(G50), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n818), .B(new_n821), .C1(G58), .C2(new_n776), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G137), .A2(new_n777), .B1(new_n772), .B2(G150), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT97), .Z(new_n825));
  AOI22_X1  g0625(.A1(G143), .A2(new_n760), .B1(new_n780), .B2(G159), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n823), .B1(new_n828), .B2(KEYINPUT34), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n759), .A2(new_n832), .B1(new_n775), .B2(new_n472), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT96), .Z(new_n834));
  OAI221_X1 g0634(.A(new_n276), .B1(new_n756), .B2(new_n375), .C1(new_n453), .C2(new_n782), .ZN(new_n835));
  INV_X1    g0635(.A(new_n767), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G87), .A2(new_n836), .B1(new_n780), .B2(G116), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n768), .B2(new_n763), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n835), .B(new_n838), .C1(G283), .C2(new_n772), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n829), .A2(new_n831), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n794), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n751), .A2(new_n748), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n742), .B(new_n841), .C1(new_n277), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n805), .A2(new_n748), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n816), .A2(new_n845), .ZN(G384));
  NOR2_X1   g0646(.A1(new_n738), .A2(new_n246), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT40), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n713), .A2(new_n725), .ZN(new_n849));
  INV_X1    g0649(.A(new_n805), .ZN(new_n850));
  INV_X1    g0650(.A(new_n447), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n441), .B(new_n678), .C1(new_n432), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n441), .A2(new_n678), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n855), .B(new_n851), .C1(new_n432), .C2(new_n441), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n849), .B(new_n850), .C1(new_n853), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  INV_X1    g0658(.A(new_n676), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n359), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n631), .A2(new_n860), .A3(new_n861), .A4(new_n355), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n326), .A2(new_n335), .A3(new_n338), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n340), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n339), .A2(new_n266), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n353), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n363), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n859), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n355), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n863), .B1(KEYINPUT37), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n359), .A2(KEYINPUT75), .A3(new_n363), .A4(KEYINPUT18), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n369), .A2(new_n872), .A3(new_n633), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n355), .B(KEYINPUT17), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n858), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n353), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n339), .A2(new_n266), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n864), .A2(new_n340), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n355), .B1(new_n880), .B2(new_n676), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n867), .A2(new_n363), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n862), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(KEYINPUT38), .C1(new_n370), .C2(new_n869), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n876), .A2(new_n885), .A3(KEYINPUT102), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT102), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n858), .C1(new_n871), .C2(new_n875), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n848), .B1(new_n857), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n848), .C1(new_n857), .C2(new_n889), .ZN(new_n893));
  INV_X1    g0693(.A(new_n857), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n631), .A2(new_n860), .A3(new_n355), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n896), .A2(new_n862), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n860), .B1(new_n874), .B2(new_n634), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n858), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n848), .B1(new_n885), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n891), .A2(new_n893), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n449), .A2(new_n849), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT104), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n672), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n885), .A2(new_n899), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n432), .A2(new_n441), .A3(new_n679), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT101), .ZN(new_n913));
  INV_X1    g0713(.A(new_n803), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n806), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n669), .A2(new_n850), .A3(new_n679), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(KEYINPUT101), .A3(new_n803), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n889), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n442), .A2(new_n447), .A3(new_n854), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n852), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n635), .A2(new_n676), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n912), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n449), .A2(new_n729), .A3(new_n734), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n637), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n847), .B1(new_n905), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n905), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(G116), .A3(new_n212), .A4(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT36), .ZN(new_n933));
  INV_X1    g0733(.A(G58), .ZN(new_n934));
  OAI21_X1  g0734(.A(G77), .B1(new_n934), .B2(new_n240), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n239), .B1(new_n935), .B2(new_n213), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n737), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n929), .A2(new_n933), .A3(new_n937), .ZN(G367));
  OAI21_X1  g0738(.A(new_n584), .B1(new_n583), .B2(new_n679), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n665), .A2(new_n678), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n699), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n653), .B1(new_n939), .B2(new_n545), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n679), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT105), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n943), .A2(new_n947), .A3(new_n945), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT42), .B2(new_n942), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT43), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n624), .A2(new_n679), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n660), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n643), .A2(new_n644), .A3(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n949), .A2(new_n952), .A3(new_n953), .A4(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n941), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n695), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n953), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(new_n948), .C2(new_n951), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n959), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n961), .B1(new_n959), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n707), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(KEYINPUT108), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n684), .A2(new_n697), .A3(new_n698), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n697), .A2(new_n698), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n683), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n691), .A2(new_n693), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n969), .B(new_n973), .C1(new_n974), .C2(new_n672), .ZN(new_n975));
  INV_X1    g0775(.A(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n798), .B2(KEYINPUT108), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n977), .A3(new_n735), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT109), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n980));
  OAI211_X1 g0780(.A(new_n960), .B(new_n980), .C1(new_n699), .C2(new_n700), .ZN(new_n981));
  INV_X1    g0781(.A(new_n980), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n701), .B2(new_n941), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT45), .B1(new_n701), .B2(new_n941), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  NOR4_X1   g0785(.A1(new_n699), .A2(new_n985), .A3(new_n960), .A4(new_n700), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n981), .B(new_n983), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT107), .B1(new_n987), .B2(new_n694), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n694), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n975), .A2(new_n977), .A3(new_n991), .A4(new_n735), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n987), .A2(KEYINPUT107), .A3(new_n694), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n979), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n968), .B1(new_n994), .B2(new_n735), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n967), .B1(new_n995), .B2(new_n740), .ZN(new_n996));
  INV_X1    g0796(.A(new_n745), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n752), .B1(new_n207), .B2(new_n390), .C1(new_n234), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n741), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT110), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n322), .B1(new_n769), .B2(new_n202), .C1(new_n790), .C2(new_n785), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n836), .A2(G77), .ZN(new_n1002));
  INV_X1    g0802(.A(G137), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n934), .B2(new_n756), .C1(new_n1003), .C2(new_n763), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1001), .B(new_n1004), .C1(G143), .C2(new_n777), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n776), .A2(G68), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n263), .B2(new_n759), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT111), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n819), .A2(G116), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n769), .A2(new_n766), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n767), .A2(new_n472), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G317), .C2(new_n764), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n776), .A2(G107), .B1(G311), .B2(new_n777), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n276), .B1(new_n759), .B2(new_n453), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G294), .B2(new_n772), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT47), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n794), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1009), .A2(KEYINPUT47), .A3(new_n1018), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1000), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n750), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n957), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n996), .A2(new_n1024), .ZN(G387));
  AND2_X1   g0825(.A1(new_n978), .A2(new_n707), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n975), .A2(new_n977), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n735), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n684), .A2(new_n750), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n322), .A2(new_n207), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1031), .A2(new_n709), .B1(G107), .B2(new_n207), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n231), .A2(new_n531), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n709), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n1034), .C1(G68), .C2(G77), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n258), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n997), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1032), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n752), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n741), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n276), .B(new_n1013), .C1(G159), .C2(new_n777), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G68), .A2(new_n780), .B1(new_n764), .B2(G150), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G50), .A2(new_n760), .B1(new_n819), .B2(G77), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n258), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n389), .A2(new_n776), .B1(new_n1046), .B2(new_n772), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n819), .A2(G294), .B1(new_n776), .B2(G283), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G317), .A2(new_n760), .B1(new_n780), .B2(G303), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n777), .A2(G322), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n768), .C2(new_n790), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT113), .Z(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(KEYINPUT49), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n322), .B1(new_n764), .B2(G326), .ZN(new_n1058));
  INV_X1    g0858(.A(G116), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1058), .C1(new_n1059), .C2(new_n767), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT49), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1048), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1042), .B1(new_n1062), .B2(new_n751), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1028), .A2(new_n740), .B1(new_n1030), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1029), .A2(new_n1064), .ZN(G393));
  XNOR2_X1  g0865(.A(new_n987), .B(new_n694), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n708), .B1(new_n1066), .B2(new_n978), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n994), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n760), .A2(G159), .B1(G150), .B2(new_n777), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n764), .A2(G143), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n240), .B2(new_n756), .C1(new_n258), .C2(new_n769), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n775), .A2(new_n277), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n322), .B1(new_n767), .B2(new_n385), .C1(new_n790), .C2(new_n202), .ZN(new_n1074));
  OR4_X1    g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n760), .A2(G311), .B1(G317), .B2(new_n777), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n756), .A2(new_n766), .B1(new_n769), .B2(new_n832), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G322), .B2(new_n764), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n276), .B1(new_n775), .B2(new_n1059), .C1(new_n375), .C2(new_n767), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G303), .B2(new_n772), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n794), .B1(new_n1075), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n238), .A2(new_n997), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1041), .B(new_n1085), .C1(G97), .C2(new_n703), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n742), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n941), .B2(new_n1023), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1066), .B2(new_n739), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1068), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(new_n842), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n741), .B1(new_n1046), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n769), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n767), .A2(new_n202), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G125), .C2(new_n764), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n322), .B1(new_n759), .B2(new_n817), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G137), .B2(new_n772), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n776), .A2(G159), .B1(G128), .B2(new_n777), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n756), .A2(new_n263), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n276), .B1(new_n756), .B2(new_n385), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n240), .A2(new_n767), .B1(new_n769), .B2(new_n472), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n759), .A2(new_n1059), .B1(new_n763), .B2(new_n832), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1105), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1073), .B1(new_n772), .B2(G107), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n766), .B2(new_n782), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1103), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1093), .B1(new_n1113), .B2(new_n751), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n909), .B2(new_n749), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n911), .B1(new_n899), .B2(new_n885), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n679), .B1(new_n730), .B2(new_n733), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n399), .A2(new_n804), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n914), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n921), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n911), .B1(new_n918), .B2(new_n921), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n909), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n805), .B1(new_n920), .B2(new_n852), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n726), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1122), .B(new_n1126), .C1(new_n1123), .C2(new_n909), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1115), .B1(new_n1130), .B2(new_n739), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n449), .A2(new_n726), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n637), .A2(new_n925), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1121), .B1(new_n812), .B2(new_n805), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1126), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n918), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n726), .A2(new_n807), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1120), .B(new_n1126), .C1(new_n1137), .C2(new_n921), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n708), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1128), .A2(new_n1129), .A3(new_n1139), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1131), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(G378));
  XNOR2_X1  g0944(.A(new_n1133), .B(KEYINPUT119), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n672), .B1(new_n894), .B2(new_n900), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n893), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1125), .A2(new_n849), .A3(new_n888), .A4(new_n886), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n892), .B1(new_n1149), .B2(new_n848), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1147), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n912), .A2(new_n922), .A3(new_n923), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n304), .A2(new_n373), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n268), .A2(new_n859), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT118), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n891), .A2(new_n893), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n924), .A3(new_n1147), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1153), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1160), .B1(new_n1153), .B2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1146), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1146), .B(KEYINPUT57), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n707), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n740), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1158), .A2(new_n748), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n322), .A2(G41), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G50), .B(new_n1172), .C1(new_n272), .C2(new_n464), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT116), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n767), .A2(new_n934), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n389), .B2(new_n780), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n375), .B2(new_n759), .C1(new_n766), .C2(new_n763), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1006), .B(new_n1172), .C1(new_n277), .C2(new_n756), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n790), .A2(new_n472), .B1(new_n782), .B2(new_n1059), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1174), .B1(new_n1180), .B2(KEYINPUT58), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n756), .A2(new_n1094), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1183), .A2(KEYINPUT117), .B1(new_n777), .B2(G125), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n776), .A2(G150), .B1(G132), .B2(new_n772), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(KEYINPUT117), .ZN(new_n1187));
  INV_X1    g0987(.A(G128), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n759), .A2(new_n1188), .B1(new_n769), .B2(new_n1003), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n272), .B(new_n464), .C1(new_n767), .C2(new_n785), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G124), .B2(new_n764), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT59), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1181), .B1(KEYINPUT58), .B2(new_n1180), .C1(new_n1192), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n751), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n842), .A2(new_n202), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1171), .A2(new_n741), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1170), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1169), .A2(new_n1201), .ZN(G375));
  AND2_X1   g1002(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(new_n739), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1121), .A2(new_n748), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n741), .B1(G68), .B2(new_n1092), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1002), .B(new_n276), .C1(new_n390), .C2(new_n775), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n759), .A2(new_n766), .B1(new_n769), .B2(new_n375), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n756), .A2(new_n472), .B1(new_n763), .B2(new_n453), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n790), .A2(new_n1059), .B1(new_n782), .B2(new_n832), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT120), .Z(new_n1212));
  NAND2_X1  g1012(.A1(new_n777), .A2(G132), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n759), .B2(new_n1003), .C1(new_n790), .C2(new_n1094), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT121), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n276), .B(new_n1175), .C1(G50), .C2(new_n776), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n769), .A2(new_n263), .B1(new_n763), .B2(new_n1188), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G159), .B2(new_n819), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1212), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1206), .B1(new_n1222), .B2(new_n751), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1204), .B1(new_n1205), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n968), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1140), .A2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1203), .A2(new_n1133), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1224), .B1(new_n1226), .B2(new_n1227), .ZN(G381));
  NAND3_X1  g1028(.A1(new_n996), .A2(new_n1090), .A3(new_n1024), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1029), .A2(new_n801), .A3(new_n1064), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1229), .A2(G381), .A3(G384), .A4(new_n1230), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT122), .Z(new_n1232));
  NAND2_X1  g1032(.A1(new_n1170), .A2(new_n1200), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n924), .B1(new_n1161), .B2(new_n1147), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1159), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1153), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1236), .A2(new_n1237), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n708), .B1(new_n1238), .B2(KEYINPUT57), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1233), .B1(new_n1239), .B2(new_n1167), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1143), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1232), .A2(new_n1241), .ZN(G407));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(G343), .C2(new_n1241), .ZN(G409));
  NAND2_X1  g1043(.A1(G387), .A2(G390), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1229), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT125), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1230), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1244), .A2(new_n1252), .A3(new_n1229), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1246), .A2(KEYINPUT125), .A3(new_n1249), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G375), .A2(G378), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1238), .A2(new_n1225), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1201), .A2(new_n1143), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n677), .A2(G213), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1227), .B1(new_n1140), .B2(KEYINPUT60), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1203), .A2(KEYINPUT60), .A3(new_n1133), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n707), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1224), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n816), .A2(new_n845), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G384), .B(new_n1224), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1266), .A2(new_n1267), .A3(KEYINPUT62), .ZN(new_n1268));
  AND4_X1   g1068(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .A4(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1143), .B1(new_n1169), .B2(new_n1201), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1201), .A2(new_n1143), .A3(new_n1258), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(KEYINPUT123), .B(new_n1259), .C1(new_n1240), .C2(new_n1143), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .A4(new_n1260), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1269), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n677), .A2(G213), .A3(G2897), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1274), .B(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1280), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1256), .B1(new_n1279), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1274), .A2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1289), .A2(new_n1257), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1255), .A2(new_n1287), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1277), .A2(new_n1288), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1273), .A2(new_n1276), .A3(new_n1260), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1282), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1286), .A2(new_n1295), .ZN(G405));
  AND2_X1   g1096(.A1(new_n1257), .A2(new_n1241), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1297), .A2(new_n1274), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1274), .ZN(new_n1299));
  OR3_X1    g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1255), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1255), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


