

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757;

  NAND2_X1 U363 ( .A1(n345), .A2(n356), .ZN(n546) );
  XNOR2_X1 U364 ( .A(n537), .B(n422), .ZN(n421) );
  AND2_X1 U365 ( .A1(n409), .A2(KEYINPUT44), .ZN(n377) );
  XNOR2_X1 U366 ( .A(n373), .B(n568), .ZN(n619) );
  OR2_X1 U367 ( .A1(n671), .A2(n670), .ZN(n665) );
  INV_X1 U368 ( .A(G953), .ZN(n751) );
  AND2_X1 U369 ( .A1(n558), .A2(n557), .ZN(n653) );
  NOR2_X1 U370 ( .A1(n558), .A2(n557), .ZN(n656) );
  NOR2_X1 U371 ( .A1(n382), .A2(n361), .ZN(n646) );
  XNOR2_X2 U372 ( .A(n601), .B(n526), .ZN(n589) );
  NAND2_X2 U373 ( .A1(n417), .A2(n606), .ZN(n601) );
  XNOR2_X2 U374 ( .A(n418), .B(G119), .ZN(n489) );
  XNOR2_X2 U375 ( .A(n378), .B(n490), .ZN(n739) );
  NAND2_X1 U376 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U377 ( .A1(n564), .A2(n563), .ZN(n565) );
  INV_X1 U378 ( .A(n549), .ZN(n668) );
  AND2_X1 U379 ( .A1(n432), .A2(n427), .ZN(n426) );
  INV_X1 U380 ( .A(n619), .ZN(n351) );
  NOR2_X1 U381 ( .A1(n646), .A2(n546), .ZN(n548) );
  XNOR2_X1 U382 ( .A(n572), .B(n571), .ZN(n701) );
  INV_X1 U383 ( .A(n700), .ZN(n339) );
  XNOR2_X1 U384 ( .A(n560), .B(n559), .ZN(n681) );
  XNOR2_X1 U385 ( .A(n416), .B(G472), .ZN(n549) );
  XNOR2_X1 U386 ( .A(n634), .B(n633), .ZN(n635) );
  XOR2_X1 U387 ( .A(n717), .B(KEYINPUT59), .Z(n718) );
  XNOR2_X1 U388 ( .A(n506), .B(n400), .ZN(n717) );
  XNOR2_X1 U389 ( .A(n402), .B(n401), .ZN(n400) );
  XNOR2_X1 U390 ( .A(n505), .B(n501), .ZN(n401) );
  XNOR2_X1 U391 ( .A(n459), .B(G140), .ZN(n746) );
  XNOR2_X1 U392 ( .A(n488), .B(G104), .ZN(n501) );
  XOR2_X1 U393 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n568) );
  XNOR2_X2 U394 ( .A(n570), .B(n569), .ZN(n682) );
  XNOR2_X2 U395 ( .A(n363), .B(n411), .ZN(n365) );
  XNOR2_X2 U396 ( .A(n500), .B(KEYINPUT39), .ZN(n580) );
  XNOR2_X2 U397 ( .A(n410), .B(n437), .ZN(n745) );
  XNOR2_X2 U398 ( .A(n516), .B(KEYINPUT4), .ZN(n410) );
  INV_X1 U399 ( .A(G237), .ZN(n444) );
  XNOR2_X1 U400 ( .A(G902), .B(KEYINPUT15), .ZN(n615) );
  XNOR2_X1 U401 ( .A(G122), .B(G107), .ZN(n514) );
  INV_X1 U402 ( .A(KEYINPUT34), .ZN(n369) );
  XNOR2_X1 U403 ( .A(G119), .B(G128), .ZN(n455) );
  XOR2_X1 U404 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n456) );
  INV_X1 U405 ( .A(KEYINPUT102), .ZN(n559) );
  NOR2_X1 U406 ( .A1(n393), .A2(n392), .ZN(n588) );
  OR2_X1 U407 ( .A1(n650), .A2(n397), .ZN(n392) );
  NOR2_X1 U408 ( .A1(n756), .A2(KEYINPUT44), .ZN(n406) );
  NOR2_X1 U409 ( .A1(G237), .A2(G953), .ZN(n438) );
  XNOR2_X1 U410 ( .A(n405), .B(KEYINPUT95), .ZN(n404) );
  INV_X1 U411 ( .A(KEYINPUT12), .ZN(n405) );
  XNOR2_X1 U412 ( .A(G134), .B(G131), .ZN(n436) );
  XNOR2_X1 U413 ( .A(KEYINPUT68), .B(G101), .ZN(n478) );
  XNOR2_X1 U414 ( .A(n494), .B(n492), .ZN(n381) );
  XOR2_X1 U415 ( .A(G125), .B(G146), .Z(n494) );
  XNOR2_X1 U416 ( .A(n491), .B(n493), .ZN(n380) );
  XNOR2_X1 U417 ( .A(KEYINPUT74), .B(KEYINPUT86), .ZN(n493) );
  INV_X1 U418 ( .A(KEYINPUT48), .ZN(n411) );
  XNOR2_X1 U419 ( .A(n366), .B(KEYINPUT38), .ZN(n684) );
  XNOR2_X1 U420 ( .A(n499), .B(n498), .ZN(n524) );
  XNOR2_X1 U421 ( .A(n510), .B(n509), .ZN(n542) );
  NOR2_X1 U422 ( .A1(n717), .A2(G902), .ZN(n510) );
  NAND2_X1 U423 ( .A1(n365), .A2(n614), .ZN(n616) );
  XNOR2_X1 U424 ( .A(n489), .B(n501), .ZN(n378) );
  XNOR2_X1 U425 ( .A(n461), .B(KEYINPUT24), .ZN(n462) );
  XOR2_X1 U426 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n466) );
  XNOR2_X1 U427 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U428 ( .A(G146), .ZN(n457) );
  XNOR2_X1 U429 ( .A(KEYINPUT10), .B(G125), .ZN(n458) );
  XNOR2_X1 U430 ( .A(n745), .B(G146), .ZN(n355) );
  INV_X1 U431 ( .A(G140), .ZN(n479) );
  NAND2_X1 U432 ( .A1(n339), .A2(n540), .ZN(n354) );
  NOR2_X1 U433 ( .A1(n556), .A2(n369), .ZN(n368) );
  NOR2_X1 U434 ( .A1(n536), .A2(n348), .ZN(n357) );
  NAND2_X1 U435 ( .A1(n564), .A2(n348), .ZN(n360) );
  AND2_X1 U436 ( .A1(n388), .A2(n486), .ZN(n586) );
  NOR2_X1 U437 ( .A1(n487), .A2(n389), .ZN(n388) );
  INV_X1 U438 ( .A(n577), .ZN(n389) );
  BUF_X1 U439 ( .A(n524), .Z(n366) );
  OR2_X1 U440 ( .A1(n544), .A2(n384), .ZN(n383) );
  NOR2_X1 U441 ( .A1(n399), .A2(KEYINPUT47), .ZN(n397) );
  NAND2_X1 U442 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U443 ( .A1(n396), .A2(KEYINPUT79), .ZN(n395) );
  INV_X1 U444 ( .A(n615), .ZN(n431) );
  NOR2_X1 U445 ( .A1(n757), .A2(n631), .ZN(n413) );
  NOR2_X1 U446 ( .A1(n415), .A2(n596), .ZN(n414) );
  NAND2_X1 U447 ( .A1(n343), .A2(n661), .ZN(n415) );
  INV_X1 U448 ( .A(n478), .ZN(n477) );
  NOR2_X1 U449 ( .A1(n616), .A2(n349), .ZN(n419) );
  NAND2_X1 U450 ( .A1(n429), .A2(n428), .ZN(n427) );
  NAND2_X1 U451 ( .A1(n615), .A2(KEYINPUT66), .ZN(n428) );
  NAND2_X1 U452 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U453 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n430) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n446) );
  AND2_X1 U455 ( .A1(n614), .A2(KEYINPUT2), .ZN(n364) );
  OR2_X1 U456 ( .A1(n624), .A2(G902), .ZN(n416) );
  XNOR2_X1 U457 ( .A(n531), .B(n435), .ZN(n539) );
  BUF_X1 U458 ( .A(n619), .Z(n732) );
  XNOR2_X1 U459 ( .A(G116), .B(KEYINPUT9), .ZN(n513) );
  XOR2_X1 U460 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n505) );
  XNOR2_X1 U461 ( .A(n503), .B(n403), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n504), .B(n404), .ZN(n403) );
  XNOR2_X1 U463 ( .A(G143), .B(G122), .ZN(n504) );
  XNOR2_X1 U464 ( .A(n386), .B(n496), .ZN(n632) );
  XNOR2_X1 U465 ( .A(n739), .B(n379), .ZN(n386) );
  XNOR2_X1 U466 ( .A(n381), .B(n380), .ZN(n379) );
  INV_X1 U467 ( .A(n616), .ZN(n617) );
  XNOR2_X1 U468 ( .A(n616), .B(n750), .ZN(n752) );
  XNOR2_X1 U469 ( .A(n462), .B(n464), .ZN(n390) );
  XNOR2_X1 U470 ( .A(G107), .B(G104), .ZN(n483) );
  XNOR2_X1 U471 ( .A(n495), .B(n481), .ZN(n482) );
  AND2_X1 U472 ( .A1(n627), .A2(G953), .ZN(n731) );
  INV_X1 U473 ( .A(n366), .ZN(n610) );
  NAND2_X1 U474 ( .A1(n352), .A2(n543), .ZN(n370) );
  NAND2_X1 U475 ( .A1(n353), .A2(n367), .ZN(n352) );
  NAND2_X1 U476 ( .A1(n358), .A2(n357), .ZN(n356) );
  NOR2_X1 U477 ( .A1(n366), .A2(n584), .ZN(n585) );
  NAND2_X1 U478 ( .A1(n362), .A2(n347), .ZN(n361) );
  XOR2_X1 U479 ( .A(n473), .B(n472), .Z(n340) );
  NOR2_X1 U480 ( .A1(n556), .A2(n555), .ZN(n341) );
  INV_X1 U481 ( .A(n670), .ZN(n385) );
  OR2_X1 U482 ( .A1(n728), .A2(G902), .ZN(n342) );
  XOR2_X1 U483 ( .A(n588), .B(n587), .Z(n343) );
  AND2_X1 U484 ( .A1(n668), .A2(n671), .ZN(n344) );
  AND2_X1 U485 ( .A1(n360), .A2(n359), .ZN(n345) );
  NAND2_X1 U486 ( .A1(n544), .A2(n384), .ZN(n346) );
  AND2_X1 U487 ( .A1(n383), .A2(n344), .ZN(n347) );
  XOR2_X1 U488 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n348) );
  INV_X1 U489 ( .A(KEYINPUT79), .ZN(n399) );
  INV_X1 U490 ( .A(KEYINPUT104), .ZN(n384) );
  INV_X1 U491 ( .A(KEYINPUT66), .ZN(n434) );
  OR2_X1 U492 ( .A1(n615), .A2(n434), .ZN(n349) );
  XNOR2_X1 U493 ( .A(n355), .B(n484), .ZN(n711) );
  AND2_X1 U494 ( .A1(n434), .A2(n424), .ZN(n350) );
  INV_X1 U495 ( .A(KEYINPUT2), .ZN(n424) );
  NAND2_X1 U496 ( .A1(n351), .A2(n419), .ZN(n432) );
  NAND2_X1 U497 ( .A1(n351), .A2(n617), .ZN(n425) );
  NAND2_X1 U498 ( .A1(n354), .A2(n369), .ZN(n353) );
  XNOR2_X1 U499 ( .A(n355), .B(n443), .ZN(n624) );
  INV_X1 U500 ( .A(n564), .ZN(n358) );
  NAND2_X1 U501 ( .A1(n536), .A2(n348), .ZN(n359) );
  NAND2_X1 U502 ( .A1(n564), .A2(KEYINPUT104), .ZN(n362) );
  XNOR2_X2 U503 ( .A(n387), .B(KEYINPUT22), .ZN(n564) );
  NAND2_X1 U504 ( .A1(n406), .A2(n407), .ZN(n374) );
  NAND2_X1 U505 ( .A1(n567), .A2(n408), .ZN(n376) );
  XNOR2_X1 U506 ( .A(n463), .B(n390), .ZN(n469) );
  XNOR2_X1 U507 ( .A(n413), .B(KEYINPUT46), .ZN(n412) );
  NAND2_X1 U508 ( .A1(n412), .A2(n414), .ZN(n363) );
  XNOR2_X1 U509 ( .A(n579), .B(KEYINPUT42), .ZN(n757) );
  NAND2_X1 U510 ( .A1(n365), .A2(n364), .ZN(n618) );
  NAND2_X1 U511 ( .A1(n368), .A2(n339), .ZN(n367) );
  XNOR2_X2 U512 ( .A(n370), .B(KEYINPUT35), .ZN(n756) );
  NOR2_X2 U513 ( .A1(n666), .A2(n371), .ZN(n537) );
  NAND2_X1 U514 ( .A1(n545), .A2(n385), .ZN(n371) );
  XNOR2_X2 U515 ( .A(n342), .B(n340), .ZN(n545) );
  XNOR2_X2 U516 ( .A(n553), .B(KEYINPUT1), .ZN(n666) );
  XNOR2_X2 U517 ( .A(n372), .B(n710), .ZN(n553) );
  NAND2_X1 U518 ( .A1(n711), .A2(n485), .ZN(n372) );
  NOR2_X2 U519 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U520 ( .A1(n564), .A2(n346), .ZN(n382) );
  NAND2_X1 U521 ( .A1(n539), .A2(n534), .ZN(n387) );
  NAND2_X1 U522 ( .A1(n589), .A2(n530), .ZN(n531) );
  NAND2_X1 U523 ( .A1(n425), .A2(n350), .ZN(n423) );
  NAND2_X1 U524 ( .A1(n426), .A2(n423), .ZN(n433) );
  XNOR2_X2 U525 ( .A(n391), .B(n538), .ZN(n700) );
  NAND2_X1 U526 ( .A1(n421), .A2(n599), .ZN(n391) );
  NAND2_X1 U527 ( .A1(n681), .A2(n398), .ZN(n394) );
  INV_X1 U528 ( .A(n681), .ZN(n396) );
  AND2_X1 U529 ( .A1(n399), .A2(KEYINPUT47), .ZN(n398) );
  INV_X1 U530 ( .A(n409), .ZN(n407) );
  XNOR2_X1 U531 ( .A(n548), .B(n547), .ZN(n409) );
  NAND2_X1 U532 ( .A1(n756), .A2(KEYINPUT44), .ZN(n408) );
  XNOR2_X1 U533 ( .A(n410), .B(n495), .ZN(n496) );
  NAND2_X1 U534 ( .A1(n632), .A2(n615), .ZN(n499) );
  INV_X1 U535 ( .A(n524), .ZN(n417) );
  XNOR2_X2 U536 ( .A(G116), .B(KEYINPUT3), .ZN(n418) );
  AND2_X1 U537 ( .A1(n425), .A2(n424), .ZN(n663) );
  INV_X1 U538 ( .A(n709), .ZN(n716) );
  NOR2_X2 U539 ( .A1(n637), .A2(n731), .ZN(n638) );
  XNOR2_X2 U540 ( .A(n420), .B(G143), .ZN(n516) );
  XNOR2_X2 U541 ( .A(G128), .B(KEYINPUT65), .ZN(n420) );
  NAND2_X1 U542 ( .A1(n421), .A2(n549), .ZN(n550) );
  INV_X1 U543 ( .A(KEYINPUT71), .ZN(n422) );
  NAND2_X1 U544 ( .A1(n433), .A2(n662), .ZN(n709) );
  BUF_X1 U545 ( .A(n709), .Z(n722) );
  BUF_X1 U546 ( .A(n632), .Z(n634) );
  XOR2_X1 U547 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n435) );
  INV_X1 U548 ( .A(KEYINPUT78), .ZN(n587) );
  INV_X1 U549 ( .A(KEYINPUT82), .ZN(n547) );
  XNOR2_X1 U550 ( .A(n480), .B(n479), .ZN(n481) );
  INV_X1 U551 ( .A(KEYINPUT110), .ZN(n569) );
  XNOR2_X1 U552 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n571) );
  INV_X1 U553 ( .A(n604), .ZN(n544) );
  XNOR2_X1 U554 ( .A(n436), .B(G137), .ZN(n437) );
  XNOR2_X1 U555 ( .A(n489), .B(n477), .ZN(n442) );
  XNOR2_X1 U556 ( .A(KEYINPUT72), .B(n438), .ZN(n502) );
  NAND2_X1 U557 ( .A1(n502), .A2(G210), .ZN(n440) );
  XNOR2_X1 U558 ( .A(G113), .B(KEYINPUT5), .ZN(n439) );
  XNOR2_X1 U559 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U560 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U561 ( .A(G472), .ZN(n622) );
  INV_X1 U562 ( .A(G902), .ZN(n485) );
  NAND2_X1 U563 ( .A1(n485), .A2(n444), .ZN(n497) );
  NAND2_X1 U564 ( .A1(n497), .A2(G214), .ZN(n606) );
  NAND2_X1 U565 ( .A1(n549), .A2(n606), .ZN(n445) );
  XNOR2_X1 U566 ( .A(n445), .B(KEYINPUT30), .ZN(n487) );
  XNOR2_X1 U567 ( .A(n446), .B(KEYINPUT14), .ZN(n451) );
  NAND2_X1 U568 ( .A1(n451), .A2(G902), .ZN(n447) );
  XNOR2_X1 U569 ( .A(n447), .B(KEYINPUT88), .ZN(n527) );
  OR2_X1 U570 ( .A1(n751), .A2(n527), .ZN(n448) );
  XOR2_X1 U571 ( .A(KEYINPUT105), .B(n448), .Z(n449) );
  NOR2_X1 U572 ( .A1(G900), .A2(n449), .ZN(n450) );
  XNOR2_X1 U573 ( .A(n450), .B(KEYINPUT106), .ZN(n453) );
  NAND2_X1 U574 ( .A1(G952), .A2(n451), .ZN(n699) );
  OR2_X1 U575 ( .A1(n699), .A2(G953), .ZN(n528) );
  INV_X1 U576 ( .A(n528), .ZN(n452) );
  NOR2_X1 U577 ( .A1(n453), .A2(n452), .ZN(n454) );
  XOR2_X1 U578 ( .A(KEYINPUT77), .B(n454), .Z(n573) );
  XNOR2_X1 U579 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U580 ( .A(n460), .B(n746), .ZN(n463) );
  XOR2_X1 U581 ( .A(KEYINPUT70), .B(KEYINPUT90), .Z(n461) );
  XOR2_X1 U582 ( .A(G137), .B(G110), .Z(n464) );
  NAND2_X1 U583 ( .A1(G234), .A2(n751), .ZN(n465) );
  XNOR2_X1 U584 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U585 ( .A(KEYINPUT80), .B(n467), .Z(n519) );
  AND2_X1 U586 ( .A1(G221), .A2(n519), .ZN(n468) );
  XNOR2_X1 U587 ( .A(n469), .B(n468), .ZN(n728) );
  XOR2_X1 U588 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n473) );
  XOR2_X1 U589 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n471) );
  NAND2_X1 U590 ( .A1(G234), .A2(n615), .ZN(n470) );
  XNOR2_X1 U591 ( .A(n471), .B(n470), .ZN(n474) );
  NAND2_X1 U592 ( .A1(n474), .A2(G217), .ZN(n472) );
  NAND2_X1 U593 ( .A1(n474), .A2(G221), .ZN(n476) );
  XNOR2_X1 U594 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n475) );
  XNOR2_X1 U595 ( .A(n476), .B(n475), .ZN(n670) );
  NOR2_X1 U596 ( .A1(n573), .A2(n665), .ZN(n486) );
  XNOR2_X1 U597 ( .A(G110), .B(n478), .ZN(n495) );
  NAND2_X1 U598 ( .A1(G227), .A2(n751), .ZN(n480) );
  XNOR2_X1 U599 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U600 ( .A(G469), .ZN(n710) );
  INV_X1 U601 ( .A(n553), .ZN(n577) );
  INV_X1 U602 ( .A(G113), .ZN(n488) );
  XNOR2_X1 U603 ( .A(n514), .B(KEYINPUT16), .ZN(n490) );
  XNOR2_X1 U604 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n492) );
  NAND2_X1 U605 ( .A1(n751), .A2(G224), .ZN(n491) );
  NAND2_X1 U606 ( .A1(n497), .A2(G210), .ZN(n498) );
  NAND2_X1 U607 ( .A1(n586), .A2(n684), .ZN(n500) );
  XNOR2_X1 U608 ( .A(G131), .B(n746), .ZN(n506) );
  NAND2_X1 U609 ( .A1(G214), .A2(n502), .ZN(n503) );
  XOR2_X1 U610 ( .A(KEYINPUT96), .B(KEYINPUT13), .Z(n508) );
  XNOR2_X1 U611 ( .A(KEYINPUT97), .B(G475), .ZN(n507) );
  XNOR2_X1 U612 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n542), .B(KEYINPUT98), .ZN(n558) );
  XOR2_X1 U614 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n512) );
  XNOR2_X1 U615 ( .A(G134), .B(KEYINPUT7), .ZN(n511) );
  XNOR2_X1 U616 ( .A(n512), .B(n511), .ZN(n518) );
  XNOR2_X1 U617 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U619 ( .A(n518), .B(n517), .Z(n521) );
  NAND2_X1 U620 ( .A1(G217), .A2(n519), .ZN(n520) );
  XNOR2_X1 U621 ( .A(n521), .B(n520), .ZN(n723) );
  NOR2_X1 U622 ( .A1(G902), .A2(n723), .ZN(n523) );
  XNOR2_X1 U623 ( .A(KEYINPUT101), .B(G478), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n523), .B(n522), .ZN(n541) );
  INV_X1 U625 ( .A(n541), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n580), .A2(n656), .ZN(n613) );
  XNOR2_X1 U627 ( .A(n613), .B(G134), .ZN(G36) );
  INV_X1 U628 ( .A(n606), .ZN(n685) );
  INV_X1 U629 ( .A(KEYINPUT67), .ZN(n525) );
  XNOR2_X1 U630 ( .A(n525), .B(KEYINPUT19), .ZN(n526) );
  XNOR2_X1 U631 ( .A(G898), .B(KEYINPUT87), .ZN(n735) );
  NAND2_X1 U632 ( .A1(G953), .A2(n735), .ZN(n740) );
  OR2_X1 U633 ( .A1(n527), .A2(n740), .ZN(n529) );
  NAND2_X1 U634 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U635 ( .A1(n542), .A2(n541), .ZN(n533) );
  INV_X1 U636 ( .A(KEYINPUT103), .ZN(n532) );
  XNOR2_X1 U637 ( .A(n533), .B(n532), .ZN(n688) );
  AND2_X1 U638 ( .A1(n688), .A2(n385), .ZN(n534) );
  INV_X1 U639 ( .A(n666), .ZN(n604) );
  XNOR2_X1 U640 ( .A(n668), .B(KEYINPUT6), .ZN(n599) );
  NOR2_X1 U641 ( .A1(n545), .A2(n599), .ZN(n535) );
  NAND2_X1 U642 ( .A1(n604), .A2(n535), .ZN(n536) );
  XOR2_X1 U643 ( .A(n546), .B(G119), .Z(G21) );
  INV_X1 U644 ( .A(KEYINPUT63), .ZN(n630) );
  INV_X1 U645 ( .A(KEYINPUT33), .ZN(n538) );
  BUF_X1 U646 ( .A(n539), .Z(n540) );
  INV_X1 U647 ( .A(n540), .ZN(n556) );
  NAND2_X1 U648 ( .A1(n542), .A2(n541), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT75), .B(n584), .ZN(n543) );
  INV_X1 U650 ( .A(n545), .ZN(n671) );
  XNOR2_X1 U651 ( .A(n550), .B(KEYINPUT93), .ZN(n678) );
  NAND2_X1 U652 ( .A1(n678), .A2(n540), .ZN(n551) );
  XNOR2_X1 U653 ( .A(n551), .B(KEYINPUT31), .ZN(n657) );
  INV_X1 U654 ( .A(n665), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n668), .A2(n552), .ZN(n554) );
  OR2_X1 U656 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U657 ( .A1(n657), .A2(n341), .ZN(n561) );
  OR2_X1 U658 ( .A1(n656), .A2(n653), .ZN(n560) );
  NOR2_X1 U659 ( .A1(n561), .A2(n681), .ZN(n566) );
  NOR2_X1 U660 ( .A1(n599), .A2(n671), .ZN(n562) );
  NAND2_X1 U661 ( .A1(n562), .A2(n666), .ZN(n563) );
  NOR2_X1 U662 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U663 ( .A1(n684), .A2(n606), .ZN(n570) );
  NAND2_X1 U664 ( .A1(n682), .A2(n688), .ZN(n572) );
  NOR2_X1 U665 ( .A1(n573), .A2(n670), .ZN(n574) );
  NAND2_X1 U666 ( .A1(n671), .A2(n574), .ZN(n597) );
  OR2_X1 U667 ( .A1(n668), .A2(n597), .ZN(n576) );
  INV_X1 U668 ( .A(KEYINPUT28), .ZN(n575) );
  XNOR2_X1 U669 ( .A(n576), .B(n575), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n591) );
  NOR2_X1 U671 ( .A1(n701), .A2(n591), .ZN(n579) );
  NAND2_X1 U672 ( .A1(n580), .A2(n653), .ZN(n583) );
  XNOR2_X1 U673 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n581) );
  XNOR2_X1 U674 ( .A(n581), .B(KEYINPUT108), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n583), .B(n582), .ZN(n631) );
  AND2_X1 U676 ( .A1(n586), .A2(n585), .ZN(n650) );
  NOR2_X1 U677 ( .A1(n681), .A2(KEYINPUT47), .ZN(n592) );
  INV_X1 U678 ( .A(n589), .ZN(n590) );
  OR2_X1 U679 ( .A1(n591), .A2(n590), .ZN(n593) );
  NOR2_X1 U680 ( .A1(n592), .A2(n593), .ZN(n595) );
  INV_X1 U681 ( .A(n593), .ZN(n651) );
  NOR2_X1 U682 ( .A1(n651), .A2(KEYINPUT47), .ZN(n594) );
  NOR2_X1 U683 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U684 ( .A(n597), .ZN(n598) );
  AND2_X1 U685 ( .A1(n653), .A2(n598), .ZN(n600) );
  NAND2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n608) );
  NOR2_X1 U687 ( .A1(n608), .A2(n601), .ZN(n603) );
  XOR2_X1 U688 ( .A(KEYINPUT83), .B(KEYINPUT36), .Z(n602) );
  XNOR2_X1 U689 ( .A(n603), .B(n602), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n605), .A2(n604), .ZN(n661) );
  NAND2_X1 U691 ( .A1(n666), .A2(n606), .ZN(n607) );
  NOR2_X1 U692 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n609), .B(KEYINPUT43), .ZN(n611) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U695 ( .A(n612), .B(KEYINPUT107), .ZN(n755) );
  AND2_X1 U696 ( .A1(n755), .A2(n613), .ZN(n614) );
  XNOR2_X1 U697 ( .A(n618), .B(KEYINPUT81), .ZN(n621) );
  INV_X1 U698 ( .A(n732), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n662) );
  NOR2_X1 U700 ( .A1(n709), .A2(n622), .ZN(n626) );
  XNOR2_X1 U701 ( .A(KEYINPUT85), .B(KEYINPUT62), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(n628) );
  INV_X1 U704 ( .A(G952), .ZN(n627) );
  NOR2_X1 U705 ( .A1(n628), .A2(n731), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(G57) );
  XOR2_X1 U707 ( .A(G131), .B(n631), .Z(G33) );
  NAND2_X1 U708 ( .A1(n716), .A2(G210), .ZN(n636) );
  XNOR2_X1 U709 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U712 ( .A(G101), .B(n565), .Z(G3) );
  NAND2_X1 U713 ( .A1(n341), .A2(n653), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n639), .B(KEYINPUT112), .ZN(n640) );
  XNOR2_X1 U715 ( .A(G104), .B(n640), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n642) );
  XNOR2_X1 U717 ( .A(G107), .B(KEYINPUT26), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(n641), .ZN(n643) );
  XOR2_X1 U719 ( .A(KEYINPUT113), .B(n643), .Z(n645) );
  NAND2_X1 U720 ( .A1(n341), .A2(n656), .ZN(n644) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U722 ( .A(n646), .B(G110), .Z(G12) );
  XOR2_X1 U723 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n648) );
  NAND2_X1 U724 ( .A1(n651), .A2(n656), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U726 ( .A(G128), .B(n649), .Z(G30) );
  XOR2_X1 U727 ( .A(G143), .B(n650), .Z(G45) );
  NAND2_X1 U728 ( .A1(n651), .A2(n653), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n652), .B(G146), .ZN(G48) );
  NAND2_X1 U730 ( .A1(n657), .A2(n653), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(KEYINPUT116), .ZN(n655) );
  XNOR2_X1 U732 ( .A(G113), .B(n655), .ZN(G15) );
  XOR2_X1 U733 ( .A(G116), .B(KEYINPUT117), .Z(n659) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(G18) );
  XOR2_X1 U736 ( .A(G125), .B(KEYINPUT37), .Z(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(G27) );
  INV_X1 U738 ( .A(n662), .ZN(n664) );
  NOR2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n707) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n667), .B(KEYINPUT50), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n676) );
  XOR2_X1 U743 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n673) );
  NAND2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U745 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT118), .ZN(n675) );
  NOR2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U749 ( .A(KEYINPUT51), .B(n679), .Z(n680) );
  NOR2_X1 U750 ( .A1(n701), .A2(n680), .ZN(n696) );
  NAND2_X1 U751 ( .A1(n396), .A2(n682), .ZN(n683) );
  XNOR2_X1 U752 ( .A(KEYINPUT121), .B(n683), .ZN(n691) );
  INV_X1 U753 ( .A(n684), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U756 ( .A(KEYINPUT120), .B(n689), .Z(n690) );
  NOR2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U758 ( .A(n692), .B(KEYINPUT122), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n700), .A2(n693), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT123), .B(n694), .Z(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U762 ( .A(n697), .B(KEYINPUT52), .ZN(n698) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n704), .B(KEYINPUT124), .ZN(n705) );
  NAND2_X1 U767 ( .A1(n705), .A2(n751), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U769 ( .A(KEYINPUT53), .B(n708), .ZN(G75) );
  NOR2_X1 U770 ( .A1(n722), .A2(n710), .ZN(n714) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  XNOR2_X1 U772 ( .A(n711), .B(n712), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n731), .A2(n715), .ZN(G54) );
  NAND2_X1 U775 ( .A1(n716), .A2(G475), .ZN(n719) );
  XNOR2_X1 U776 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X2 U777 ( .A1(n720), .A2(n731), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U779 ( .A(n722), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n727), .A2(G478), .ZN(n725) );
  XOR2_X1 U781 ( .A(n723), .B(KEYINPUT125), .Z(n724) );
  XNOR2_X1 U782 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U783 ( .A1(n731), .A2(n726), .ZN(G63) );
  NAND2_X1 U784 ( .A1(n727), .A2(G217), .ZN(n729) );
  XNOR2_X1 U785 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n731), .A2(n730), .ZN(G66) );
  NOR2_X1 U787 ( .A1(n732), .A2(G953), .ZN(n737) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n733) );
  XOR2_X1 U789 ( .A(KEYINPUT61), .B(n733), .Z(n734) );
  NOR2_X1 U790 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n737), .A2(n736), .ZN(n743) );
  XNOR2_X1 U792 ( .A(G101), .B(G110), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n741) );
  NAND2_X1 U794 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U795 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U796 ( .A(KEYINPUT126), .B(n744), .ZN(G69) );
  XNOR2_X1 U797 ( .A(n745), .B(n746), .ZN(n749) );
  XOR2_X1 U798 ( .A(G227), .B(n749), .Z(n747) );
  NAND2_X1 U799 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(G953), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n749), .B(KEYINPUT127), .ZN(n750) );
  NAND2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U803 ( .A1(n754), .A2(n753), .ZN(G72) );
  XNOR2_X1 U804 ( .A(G140), .B(n755), .ZN(G42) );
  XOR2_X1 U805 ( .A(n756), .B(G122), .Z(G24) );
  XOR2_X1 U806 ( .A(G137), .B(n757), .Z(G39) );
endmodule

