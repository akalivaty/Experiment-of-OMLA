

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  AND2_X1 U323 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U324 ( .A(KEYINPUT96), .B(KEYINPUT27), .ZN(n367) );
  XNOR2_X1 U325 ( .A(n551), .B(n367), .ZN(n390) );
  XNOR2_X1 U326 ( .A(n447), .B(n291), .ZN(n363) );
  XNOR2_X1 U327 ( .A(n364), .B(n363), .ZN(n365) );
  INV_X1 U328 ( .A(G43GAT), .ZN(n460) );
  XNOR2_X1 U329 ( .A(n460), .B(KEYINPUT40), .ZN(n461) );
  XNOR2_X1 U330 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  XOR2_X1 U331 ( .A(G43GAT), .B(G134GAT), .Z(n316) );
  XOR2_X1 U332 ( .A(KEYINPUT0), .B(G127GAT), .Z(n335) );
  XNOR2_X1 U333 ( .A(n316), .B(n335), .ZN(n293) );
  XNOR2_X1 U334 ( .A(G99GAT), .B(G120GAT), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n292), .B(G71GAT), .ZN(n449) );
  XNOR2_X1 U336 ( .A(n293), .B(n449), .ZN(n294) );
  XOR2_X1 U337 ( .A(n294), .B(KEYINPUT20), .Z(n296) );
  XOR2_X1 U338 ( .A(G113GAT), .B(G15GAT), .Z(n436) );
  XNOR2_X1 U339 ( .A(n436), .B(KEYINPUT81), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n298) );
  NAND2_X1 U342 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(n300), .B(n299), .Z(n307) );
  XOR2_X1 U345 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(G176GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U348 ( .A(n303), .B(G183GAT), .Z(n305) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n366) );
  XNOR2_X1 U351 ( .A(n366), .B(KEYINPUT84), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n519) );
  XOR2_X1 U353 ( .A(G106GAT), .B(G218GAT), .Z(n309) );
  XNOR2_X1 U354 ( .A(G190GAT), .B(KEYINPUT76), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n311) );
  INV_X1 U356 ( .A(G92GAT), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U358 ( .A(G85GAT), .B(KEYINPUT74), .Z(n453) );
  XOR2_X1 U359 ( .A(G36GAT), .B(n453), .Z(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U361 ( .A(G50GAT), .B(G162GAT), .Z(n375) );
  XNOR2_X1 U362 ( .A(n314), .B(n375), .ZN(n318) );
  XNOR2_X1 U363 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n315), .B(KEYINPUT8), .ZN(n430) );
  XNOR2_X1 U365 ( .A(n430), .B(n316), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n320) );
  NAND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XOR2_X1 U369 ( .A(n320), .B(n319), .Z(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT77), .B(KEYINPUT66), .Z(n324) );
  XNOR2_X1 U372 ( .A(KEYINPUT65), .B(KEYINPUT9), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(G99GAT), .B(n325), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n548) );
  XNOR2_X1 U376 ( .A(n548), .B(KEYINPUT108), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n328), .B(KEYINPUT36), .ZN(n589) );
  XOR2_X1 U378 ( .A(KEYINPUT6), .B(G148GAT), .Z(n330) );
  XNOR2_X1 U379 ( .A(G1GAT), .B(G113GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U381 ( .A(G85GAT), .B(G162GAT), .Z(n332) );
  XNOR2_X1 U382 ( .A(G120GAT), .B(KEYINPUT76), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n353) );
  XOR2_X1 U385 ( .A(n335), .B(KEYINPUT1), .Z(n337) );
  NAND2_X1 U386 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U387 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U388 ( .A(KEYINPUT88), .B(KEYINPUT2), .Z(n339) );
  XNOR2_X1 U389 ( .A(KEYINPUT89), .B(G155GAT), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U391 ( .A(KEYINPUT3), .B(n340), .Z(n380) );
  XOR2_X1 U392 ( .A(n341), .B(n380), .Z(n343) );
  XNOR2_X1 U393 ( .A(G29GAT), .B(G134GAT), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n351) );
  XOR2_X1 U395 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n345) );
  XNOR2_X1 U396 ( .A(G141GAT), .B(KEYINPUT92), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U398 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n347) );
  XNOR2_X1 U399 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U401 ( .A(n349), .B(n348), .Z(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n553) );
  INV_X1 U404 ( .A(KEYINPUT87), .ZN(n354) );
  NAND2_X1 U405 ( .A1(KEYINPUT21), .A2(n354), .ZN(n357) );
  INV_X1 U406 ( .A(KEYINPUT21), .ZN(n355) );
  NAND2_X1 U407 ( .A1(n355), .A2(KEYINPUT87), .ZN(n356) );
  NAND2_X1 U408 ( .A1(n357), .A2(n356), .ZN(n359) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(G218GAT), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n360), .B(G211GAT), .ZN(n385) );
  XNOR2_X1 U412 ( .A(KEYINPUT95), .B(n385), .ZN(n362) );
  XOR2_X1 U413 ( .A(G36GAT), .B(G8GAT), .Z(n433) );
  XNOR2_X1 U414 ( .A(n433), .B(G204GAT), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U416 ( .A(G92GAT), .B(G64GAT), .Z(n447) );
  XOR2_X1 U417 ( .A(n366), .B(n365), .Z(n551) );
  NOR2_X1 U418 ( .A1(n553), .A2(n390), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n368), .B(KEYINPUT97), .ZN(n518) );
  XNOR2_X1 U420 ( .A(G78GAT), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n369), .B(KEYINPUT72), .ZN(n370) );
  XOR2_X1 U422 ( .A(n370), .B(KEYINPUT73), .Z(n372) );
  XNOR2_X1 U423 ( .A(G148GAT), .B(G106GAT), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n446) );
  XOR2_X1 U425 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n374) );
  XNOR2_X1 U426 ( .A(KEYINPUT86), .B(KEYINPUT24), .ZN(n373) );
  XNOR2_X1 U427 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U428 ( .A(n375), .B(KEYINPUT22), .Z(n377) );
  NAND2_X1 U429 ( .A1(G228GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U431 ( .A(n379), .B(n378), .Z(n382) );
  XOR2_X1 U432 ( .A(G141GAT), .B(G22GAT), .Z(n435) );
  XNOR2_X1 U433 ( .A(n435), .B(n380), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U435 ( .A(n446), .B(n383), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n556) );
  XNOR2_X1 U437 ( .A(KEYINPUT28), .B(n556), .ZN(n522) );
  NOR2_X1 U438 ( .A1(n518), .A2(n522), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n386), .B(KEYINPUT98), .ZN(n388) );
  XOR2_X1 U440 ( .A(n519), .B(KEYINPUT85), .Z(n387) );
  NAND2_X1 U441 ( .A1(n388), .A2(n387), .ZN(n401) );
  NAND2_X1 U442 ( .A1(n556), .A2(n519), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n389), .B(KEYINPUT26), .ZN(n575) );
  NOR2_X1 U444 ( .A1(n390), .A2(n575), .ZN(n396) );
  XNOR2_X1 U445 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n391), .B(KEYINPUT100), .ZN(n394) );
  NOR2_X1 U447 ( .A1(n519), .A2(n551), .ZN(n392) );
  NOR2_X1 U448 ( .A1(n556), .A2(n392), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  NOR2_X1 U450 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n397), .B(KEYINPUT101), .ZN(n398) );
  NAND2_X1 U452 ( .A1(n398), .A2(n553), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n399), .B(KEYINPUT102), .ZN(n400) );
  NAND2_X1 U454 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n402), .B(KEYINPUT103), .ZN(n465) );
  NOR2_X1 U456 ( .A1(n589), .A2(n465), .ZN(n422) );
  XOR2_X1 U457 ( .A(G211GAT), .B(KEYINPUT14), .Z(n404) );
  XNOR2_X1 U458 ( .A(G22GAT), .B(KEYINPUT79), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U460 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n406) );
  XNOR2_X1 U461 ( .A(G183GAT), .B(KEYINPUT80), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n421) );
  XOR2_X1 U464 ( .A(G155GAT), .B(G71GAT), .Z(n410) );
  XNOR2_X1 U465 ( .A(G1GAT), .B(G127GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n419) );
  XNOR2_X1 U467 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n411), .B(KEYINPUT13), .ZN(n448) );
  XOR2_X1 U469 ( .A(n448), .B(KEYINPUT15), .Z(n413) );
  NAND2_X1 U470 ( .A1(G231GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U472 ( .A(G64GAT), .B(G78GAT), .Z(n415) );
  XNOR2_X1 U473 ( .A(G8GAT), .B(G15GAT), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U475 ( .A(n417), .B(n416), .Z(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n545) );
  NAND2_X1 U478 ( .A1(n422), .A2(n545), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n423), .B(KEYINPUT37), .ZN(n497) );
  XOR2_X1 U480 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n425) );
  XNOR2_X1 U481 ( .A(G169GAT), .B(G1GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U483 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n427) );
  XNOR2_X1 U484 ( .A(KEYINPUT68), .B(G197GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n442) );
  XOR2_X1 U487 ( .A(n430), .B(KEYINPUT70), .Z(n432) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n440) );
  XOR2_X1 U491 ( .A(G50GAT), .B(G43GAT), .Z(n438) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n577) );
  INV_X1 U496 ( .A(n577), .ZN(n536) );
  XOR2_X1 U497 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n444) );
  XNOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n457) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n455) );
  XOR2_X1 U502 ( .A(n449), .B(KEYINPUT32), .Z(n451) );
  NAND2_X1 U503 ( .A1(G230GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n457), .B(n456), .ZN(n484) );
  INV_X1 U508 ( .A(n484), .ZN(n582) );
  NOR2_X1 U509 ( .A1(n536), .A2(n582), .ZN(n466) );
  AND2_X1 U510 ( .A1(n497), .A2(n466), .ZN(n459) );
  INV_X1 U511 ( .A(KEYINPUT38), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n482) );
  NOR2_X1 U513 ( .A1(n519), .A2(n482), .ZN(n462) );
  INV_X1 U514 ( .A(n548), .ZN(n568) );
  NOR2_X1 U515 ( .A1(n568), .A2(n545), .ZN(n463) );
  XOR2_X1 U516 ( .A(KEYINPUT16), .B(n463), .Z(n464) );
  NOR2_X1 U517 ( .A1(n465), .A2(n464), .ZN(n485) );
  NAND2_X1 U518 ( .A1(n466), .A2(n485), .ZN(n475) );
  NOR2_X1 U519 ( .A1(n553), .A2(n475), .ZN(n467) );
  XOR2_X1 U520 ( .A(KEYINPUT34), .B(n467), .Z(n468) );
  XNOR2_X1 U521 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NOR2_X1 U522 ( .A1(n551), .A2(n475), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT104), .B(n469), .Z(n470) );
  XNOR2_X1 U524 ( .A(G8GAT), .B(n470), .ZN(G1325GAT) );
  NOR2_X1 U525 ( .A1(n475), .A2(n519), .ZN(n474) );
  XOR2_X1 U526 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n472) );
  XNOR2_X1 U527 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  INV_X1 U530 ( .A(n522), .ZN(n502) );
  NOR2_X1 U531 ( .A1(n502), .A2(n475), .ZN(n477) );
  XNOR2_X1 U532 ( .A(G22GAT), .B(KEYINPUT107), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n477), .B(n476), .ZN(G1327GAT) );
  NOR2_X1 U534 ( .A1(n482), .A2(n553), .ZN(n479) );
  XNOR2_X1 U535 ( .A(KEYINPUT109), .B(KEYINPUT39), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U537 ( .A(G29GAT), .B(n480), .Z(G1328GAT) );
  NOR2_X1 U538 ( .A1(n551), .A2(n482), .ZN(n481) );
  XOR2_X1 U539 ( .A(G36GAT), .B(n481), .Z(G1329GAT) );
  NOR2_X1 U540 ( .A1(n482), .A2(n502), .ZN(n483) );
  XOR2_X1 U541 ( .A(G50GAT), .B(n483), .Z(G1331GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT41), .B(n484), .Z(n539) );
  NOR2_X1 U543 ( .A1(n577), .A2(n539), .ZN(n496) );
  NAND2_X1 U544 ( .A1(n496), .A2(n485), .ZN(n492) );
  NOR2_X1 U545 ( .A1(n553), .A2(n492), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U548 ( .A(G57GAT), .B(n488), .Z(G1332GAT) );
  NOR2_X1 U549 ( .A1(n551), .A2(n492), .ZN(n489) );
  XOR2_X1 U550 ( .A(G64GAT), .B(n489), .Z(G1333GAT) );
  NOR2_X1 U551 ( .A1(n519), .A2(n492), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1334GAT) );
  NOR2_X1 U554 ( .A1(n502), .A2(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G78GAT), .B(n495), .ZN(G1335GAT) );
  NAND2_X1 U558 ( .A1(n497), .A2(n496), .ZN(n501) );
  NOR2_X1 U559 ( .A1(n553), .A2(n501), .ZN(n498) );
  XOR2_X1 U560 ( .A(G85GAT), .B(n498), .Z(G1336GAT) );
  NOR2_X1 U561 ( .A1(n551), .A2(n501), .ZN(n499) );
  XOR2_X1 U562 ( .A(G92GAT), .B(n499), .Z(G1337GAT) );
  NOR2_X1 U563 ( .A1(n519), .A2(n501), .ZN(n500) );
  XOR2_X1 U564 ( .A(G99GAT), .B(n500), .Z(G1338GAT) );
  NOR2_X1 U565 ( .A1(n502), .A2(n501), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT113), .B(KEYINPUT44), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G106GAT), .B(n505), .ZN(G1339GAT) );
  NOR2_X1 U569 ( .A1(n589), .A2(n545), .ZN(n506) );
  XNOR2_X1 U570 ( .A(KEYINPUT45), .B(n506), .ZN(n508) );
  NOR2_X1 U571 ( .A1(n577), .A2(n582), .ZN(n507) );
  AND2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT115), .ZN(n516) );
  XOR2_X1 U574 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n511) );
  INV_X1 U575 ( .A(n539), .ZN(n563) );
  NAND2_X1 U576 ( .A1(n577), .A2(n563), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(n513) );
  NAND2_X1 U578 ( .A1(n548), .A2(n545), .ZN(n512) );
  NOR2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(KEYINPUT47), .B(n514), .ZN(n515) );
  AND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT48), .ZN(n550) );
  NOR2_X1 U583 ( .A1(n550), .A2(n518), .ZN(n535) );
  INV_X1 U584 ( .A(n519), .ZN(n569) );
  NAND2_X1 U585 ( .A1(n535), .A2(n569), .ZN(n520) );
  XNOR2_X1 U586 ( .A(KEYINPUT116), .B(n520), .ZN(n521) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n577), .A2(n530), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G113GAT), .B(n523), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .Z(n525) );
  NAND2_X1 U591 ( .A1(n530), .A2(n563), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n527) );
  INV_X1 U595 ( .A(n545), .ZN(n585) );
  NAND2_X1 U596 ( .A1(n530), .A2(n585), .ZN(n526) );
  XNOR2_X1 U597 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n532) );
  NAND2_X1 U600 ( .A1(n530), .A2(n568), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U602 ( .A(G134GAT), .B(n533), .Z(G1343GAT) );
  INV_X1 U603 ( .A(n575), .ZN(n534) );
  NAND2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n536), .A2(n547), .ZN(n537) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n537), .Z(n538) );
  XNOR2_X1 U607 ( .A(KEYINPUT120), .B(n538), .ZN(G1344GAT) );
  NOR2_X1 U608 ( .A1(n539), .A2(n547), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n541) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U612 ( .A(KEYINPUT121), .B(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n545), .A2(n547), .ZN(n546) );
  XOR2_X1 U615 ( .A(G155GAT), .B(n546), .Z(G1346GAT) );
  NOR2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(G162GAT), .B(n549), .Z(G1347GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT54), .B(n552), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT64), .ZN(n576) );
  NOR2_X1 U622 ( .A1(n576), .A2(n556), .ZN(n557) );
  XOR2_X1 U623 ( .A(n557), .B(KEYINPUT55), .Z(n570) );
  AND2_X1 U624 ( .A1(n569), .A2(n570), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n577), .A2(n566), .ZN(n559) );
  XOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n561) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n562), .Z(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n563), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n566), .A2(n585), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n573) );
  AND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G190GAT), .B(n574), .Z(G1351GAT) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT127), .Z(n579) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n587), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n587), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U652 ( .A(n587), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(n590), .B(KEYINPUT62), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

