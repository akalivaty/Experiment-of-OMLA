

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745;

  OR2_X1 U370 ( .A1(n745), .A2(n527), .ZN(n528) );
  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n499) );
  NOR2_X1 U372 ( .A1(n617), .A2(n471), .ZN(n473) );
  XNOR2_X1 U373 ( .A(n435), .B(n434), .ZN(n524) );
  NOR2_X2 U374 ( .A1(n534), .A2(n533), .ZN(n577) );
  XNOR2_X2 U375 ( .A(n473), .B(n472), .ZN(n564) );
  INV_X1 U376 ( .A(n635), .ZN(n348) );
  NAND2_X2 U377 ( .A1(n371), .A2(n369), .ZN(n713) );
  NAND2_X1 U378 ( .A1(n368), .A2(n613), .ZN(n371) );
  NAND2_X1 U379 ( .A1(n373), .A2(n366), .ZN(n368) );
  AND2_X1 U380 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U381 ( .A1(n362), .A2(n562), .ZN(n598) );
  NOR2_X1 U382 ( .A1(n605), .A2(n602), .ZN(n581) );
  XNOR2_X1 U383 ( .A(n397), .B(KEYINPUT41), .ZN(n697) );
  XNOR2_X1 U384 ( .A(n475), .B(n404), .ZN(n556) );
  XNOR2_X1 U385 ( .A(n511), .B(n361), .ZN(n532) );
  XNOR2_X1 U386 ( .A(n458), .B(n457), .ZN(n671) );
  OR2_X1 U387 ( .A1(n636), .A2(G902), .ZN(n435) );
  XNOR2_X1 U388 ( .A(n468), .B(n406), .ZN(n494) );
  XNOR2_X1 U389 ( .A(n469), .B(KEYINPUT10), .ZN(n730) );
  XNOR2_X1 U390 ( .A(G143), .B(KEYINPUT12), .ZN(n502) );
  XOR2_X1 U391 ( .A(G113), .B(G104), .Z(n507) );
  XNOR2_X1 U392 ( .A(KEYINPUT24), .B(G110), .ZN(n418) );
  XNOR2_X1 U393 ( .A(KEYINPUT88), .B(G119), .ZN(n419) );
  XNOR2_X1 U394 ( .A(G146), .B(G125), .ZN(n469) );
  XNOR2_X1 U395 ( .A(G140), .B(G137), .ZN(n420) );
  INV_X1 U396 ( .A(n528), .ZN(n381) );
  XOR2_X1 U397 ( .A(n564), .B(n588), .Z(n681) );
  INV_X1 U398 ( .A(KEYINPUT2), .ZN(n367) );
  NAND2_X1 U399 ( .A1(n365), .A2(n363), .ZN(n373) );
  NAND2_X1 U400 ( .A1(n359), .A2(n610), .ZN(n365) );
  NAND2_X1 U401 ( .A1(n364), .A2(n355), .ZN(n363) );
  XOR2_X1 U402 ( .A(G110), .B(KEYINPUT67), .Z(n467) );
  NAND2_X1 U403 ( .A1(n713), .A2(G475), .ZN(n403) );
  AND2_X1 U404 ( .A1(n584), .A2(n563), .ZN(n362) );
  NOR2_X1 U405 ( .A1(n650), .A2(n658), .ZN(n584) );
  NAND2_X1 U406 ( .A1(n348), .A2(n383), .ZN(n382) );
  NOR2_X1 U407 ( .A1(n528), .A2(n385), .ZN(n383) );
  XNOR2_X1 U408 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n416) );
  INV_X1 U409 ( .A(n610), .ZN(n364) );
  XNOR2_X1 U410 ( .A(n494), .B(n407), .ZN(n733) );
  XNOR2_X1 U411 ( .A(KEYINPUT4), .B(G131), .ZN(n407) );
  NAND2_X1 U412 ( .A1(n681), .A2(n680), .ZN(n686) );
  XNOR2_X1 U413 ( .A(n512), .B(G475), .ZN(n361) );
  XOR2_X1 U414 ( .A(G122), .B(G107), .Z(n485) );
  XNOR2_X1 U415 ( .A(n452), .B(n451), .ZN(n464) );
  XNOR2_X1 U416 ( .A(G119), .B(KEYINPUT3), .ZN(n451) );
  XNOR2_X1 U417 ( .A(G101), .B(G116), .ZN(n450) );
  XNOR2_X1 U418 ( .A(G101), .B(G107), .ZN(n408) );
  XOR2_X1 U419 ( .A(KEYINPUT74), .B(G104), .Z(n409) );
  XNOR2_X1 U420 ( .A(n733), .B(G146), .ZN(n455) );
  XNOR2_X1 U421 ( .A(n393), .B(n391), .ZN(n390) );
  XNOR2_X1 U422 ( .A(n468), .B(n392), .ZN(n391) );
  XNOR2_X1 U423 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X1 U424 ( .A(n593), .B(n592), .ZN(n601) );
  INV_X1 U425 ( .A(KEYINPUT39), .ZN(n592) );
  AND2_X1 U426 ( .A1(n389), .A2(n350), .ZN(n378) );
  NAND2_X1 U427 ( .A1(n388), .A2(n349), .ZN(n377) );
  XNOR2_X1 U428 ( .A(n498), .B(n497), .ZN(n534) );
  NAND2_X1 U429 ( .A1(n354), .A2(n373), .ZN(n369) );
  XOR2_X1 U430 ( .A(G131), .B(KEYINPUT94), .Z(n501) );
  XOR2_X1 U431 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n503) );
  INV_X1 U432 ( .A(KEYINPUT105), .ZN(n443) );
  XNOR2_X1 U433 ( .A(n470), .B(n352), .ZN(n394) );
  XOR2_X1 U434 ( .A(KEYINPUT4), .B(KEYINPUT17), .Z(n470) );
  XNOR2_X1 U435 ( .A(n466), .B(n467), .ZN(n395) );
  XNOR2_X1 U436 ( .A(n469), .B(KEYINPUT18), .ZN(n392) );
  NAND2_X1 U437 ( .A1(G234), .A2(G237), .ZN(n476) );
  XNOR2_X1 U438 ( .A(G137), .B(G113), .ZN(n447) );
  AND2_X1 U439 ( .A1(n471), .A2(KEYINPUT64), .ZN(n370) );
  AND2_X1 U440 ( .A1(n372), .A2(n471), .ZN(n366) );
  XNOR2_X1 U441 ( .A(n599), .B(KEYINPUT48), .ZN(n609) );
  INV_X1 U442 ( .A(KEYINPUT1), .ZN(n374) );
  INV_X1 U443 ( .A(n686), .ZN(n398) );
  INV_X1 U444 ( .A(n684), .ZN(n399) );
  XNOR2_X1 U445 ( .A(n654), .B(n360), .ZN(n600) );
  INV_X1 U446 ( .A(KEYINPUT102), .ZN(n360) );
  XNOR2_X1 U447 ( .A(n568), .B(n567), .ZN(n573) );
  XNOR2_X1 U448 ( .A(n555), .B(n554), .ZN(n585) );
  XNOR2_X1 U449 ( .A(n553), .B(KEYINPUT28), .ZN(n554) );
  XNOR2_X1 U450 ( .A(n396), .B(n465), .ZN(n718) );
  XNOR2_X1 U451 ( .A(n490), .B(n351), .ZN(n491) );
  XNOR2_X1 U452 ( .A(n455), .B(n414), .ZN(n709) );
  NAND2_X1 U453 ( .A1(n378), .A2(n377), .ZN(n376) );
  AND2_X1 U454 ( .A1(n533), .A2(n534), .ZN(n654) );
  INV_X1 U455 ( .A(KEYINPUT60), .ZN(n400) );
  INV_X1 U456 ( .A(n379), .ZN(n519) );
  AND2_X1 U457 ( .A1(n517), .A2(KEYINPUT34), .ZN(n349) );
  OR2_X1 U458 ( .A1(n517), .A2(KEYINPUT34), .ZN(n350) );
  XOR2_X1 U459 ( .A(n489), .B(n488), .Z(n351) );
  AND2_X1 U460 ( .A1(G224), .A2(n737), .ZN(n352) );
  OR2_X1 U461 ( .A1(n560), .A2(n542), .ZN(n353) );
  AND2_X1 U462 ( .A1(n372), .A2(n370), .ZN(n354) );
  OR2_X1 U463 ( .A1(KEYINPUT71), .A2(KEYINPUT2), .ZN(n355) );
  XOR2_X1 U464 ( .A(n633), .B(n632), .Z(n356) );
  XNOR2_X2 U465 ( .A(n357), .B(n513), .ZN(n635) );
  NAND2_X1 U466 ( .A1(n376), .A2(n574), .ZN(n357) );
  NAND2_X1 U467 ( .A1(n358), .A2(n355), .ZN(n359) );
  INV_X1 U468 ( .A(n611), .ZN(n358) );
  INV_X1 U469 ( .A(KEYINPUT44), .ZN(n385) );
  XNOR2_X1 U470 ( .A(n403), .B(n356), .ZN(n402) );
  NAND2_X1 U471 ( .A1(n709), .A2(n495), .ZN(n375) );
  INV_X1 U472 ( .A(n611), .ZN(n721) );
  NAND2_X1 U473 ( .A1(n611), .A2(n367), .ZN(n372) );
  XNOR2_X2 U474 ( .A(n386), .B(n546), .ZN(n611) );
  NAND2_X1 U475 ( .A1(n440), .A2(n379), .ZN(n442) );
  XNOR2_X2 U476 ( .A(n538), .B(n374), .ZN(n379) );
  NAND2_X1 U477 ( .A1(n402), .A2(n634), .ZN(n401) );
  XNOR2_X2 U478 ( .A(n375), .B(n415), .ZN(n538) );
  NAND2_X1 U479 ( .A1(n380), .A2(n385), .ZN(n384) );
  NAND2_X1 U480 ( .A1(n348), .A2(n381), .ZN(n380) );
  NAND2_X1 U481 ( .A1(n384), .A2(n382), .ZN(n387) );
  NAND2_X1 U482 ( .A1(n387), .A2(n545), .ZN(n386) );
  XNOR2_X2 U483 ( .A(n463), .B(n462), .ZN(n691) );
  INV_X1 U484 ( .A(n691), .ZN(n388) );
  NAND2_X1 U485 ( .A1(n691), .A2(n484), .ZN(n389) );
  XNOR2_X1 U486 ( .A(n718), .B(n390), .ZN(n617) );
  XNOR2_X1 U487 ( .A(n464), .B(KEYINPUT16), .ZN(n396) );
  NAND2_X1 U488 ( .A1(n589), .A2(n697), .ZN(n590) );
  NAND2_X1 U489 ( .A1(n399), .A2(n398), .ZN(n397) );
  XNOR2_X1 U490 ( .A(n401), .B(n400), .ZN(G60) );
  XNOR2_X1 U491 ( .A(KEYINPUT72), .B(KEYINPUT19), .ZN(n404) );
  NOR2_X1 U492 ( .A1(n692), .A2(n699), .ZN(n405) );
  INV_X1 U493 ( .A(KEYINPUT5), .ZN(n446) );
  XNOR2_X1 U494 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U495 ( .A(n449), .B(n448), .ZN(n453) );
  BUF_X1 U496 ( .A(n691), .Z(n699) );
  INV_X1 U497 ( .A(n665), .ZN(n515) );
  XNOR2_X1 U498 ( .A(n566), .B(KEYINPUT107), .ZN(n567) );
  INV_X1 U499 ( .A(KEYINPUT109), .ZN(n553) );
  XNOR2_X1 U500 ( .A(n492), .B(n491), .ZN(n493) );
  AND2_X1 U501 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X2 U502 ( .A(G128), .B(G143), .ZN(n468) );
  INV_X1 U503 ( .A(G134), .ZN(n406) );
  XNOR2_X1 U504 ( .A(n420), .B(KEYINPUT86), .ZN(n729) );
  XNOR2_X1 U505 ( .A(n467), .B(n729), .ZN(n413) );
  XNOR2_X1 U506 ( .A(n409), .B(n408), .ZN(n411) );
  INV_X2 U507 ( .A(G953), .ZN(n737) );
  NAND2_X1 U508 ( .A1(n737), .A2(G227), .ZN(n410) );
  XNOR2_X1 U509 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U510 ( .A(n413), .B(n412), .ZN(n414) );
  INV_X1 U511 ( .A(G902), .ZN(n495) );
  INV_X1 U512 ( .A(G469), .ZN(n415) );
  NAND2_X1 U513 ( .A1(n737), .A2(G234), .ZN(n417) );
  XNOR2_X1 U514 ( .A(n417), .B(n416), .ZN(n487) );
  NAND2_X1 U515 ( .A1(n487), .A2(G221), .ZN(n423) );
  XNOR2_X1 U516 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U517 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U518 ( .A(n423), .B(n422), .ZN(n428) );
  XNOR2_X1 U519 ( .A(G128), .B(KEYINPUT87), .ZN(n425) );
  XNOR2_X1 U520 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U521 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U522 ( .A(n730), .B(n426), .ZN(n427) );
  XNOR2_X1 U523 ( .A(n428), .B(n427), .ZN(n636) );
  INV_X1 U524 ( .A(KEYINPUT15), .ZN(n429) );
  XNOR2_X1 U525 ( .A(n429), .B(G902), .ZN(n471) );
  INV_X1 U526 ( .A(n471), .ZN(n612) );
  NAND2_X1 U527 ( .A1(G234), .A2(n612), .ZN(n430) );
  XNOR2_X1 U528 ( .A(KEYINPUT20), .B(n430), .ZN(n436) );
  NAND2_X1 U529 ( .A1(n436), .A2(G217), .ZN(n433) );
  INV_X1 U530 ( .A(KEYINPUT73), .ZN(n431) );
  XNOR2_X1 U531 ( .A(n431), .B(KEYINPUT25), .ZN(n432) );
  XNOR2_X1 U532 ( .A(n433), .B(n432), .ZN(n434) );
  INV_X1 U533 ( .A(n524), .ZN(n666) );
  NAND2_X1 U534 ( .A1(n436), .A2(G221), .ZN(n439) );
  INV_X1 U535 ( .A(KEYINPUT90), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n437), .B(KEYINPUT21), .ZN(n438) );
  XNOR2_X1 U537 ( .A(n439), .B(n438), .ZN(n665) );
  NAND2_X1 U538 ( .A1(n666), .A2(n665), .ZN(n669) );
  INV_X1 U539 ( .A(n669), .ZN(n440) );
  INV_X1 U540 ( .A(KEYINPUT70), .ZN(n441) );
  XNOR2_X2 U541 ( .A(n442), .B(n441), .ZN(n535) );
  XNOR2_X1 U542 ( .A(n535), .B(n443), .ZN(n461) );
  XOR2_X1 U543 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n445) );
  NAND2_X1 U544 ( .A1(n499), .A2(G210), .ZN(n444) );
  XNOR2_X1 U545 ( .A(n445), .B(n444), .ZN(n449) );
  INV_X1 U546 ( .A(n450), .ZN(n452) );
  XNOR2_X1 U547 ( .A(n453), .B(n464), .ZN(n454) );
  XNOR2_X1 U548 ( .A(n455), .B(n454), .ZN(n626) );
  NAND2_X1 U549 ( .A1(n626), .A2(n495), .ZN(n458) );
  XNOR2_X1 U550 ( .A(KEYINPUT68), .B(KEYINPUT93), .ZN(n456) );
  XNOR2_X1 U551 ( .A(n456), .B(G472), .ZN(n457) );
  INV_X1 U552 ( .A(KEYINPUT6), .ZN(n459) );
  XNOR2_X1 U553 ( .A(n671), .B(n459), .ZN(n579) );
  INV_X1 U554 ( .A(n579), .ZN(n460) );
  NAND2_X1 U555 ( .A1(n461), .A2(n460), .ZN(n463) );
  XNOR2_X1 U556 ( .A(KEYINPUT81), .B(KEYINPUT33), .ZN(n462) );
  XOR2_X1 U557 ( .A(n507), .B(n485), .Z(n465) );
  XOR2_X1 U558 ( .A(KEYINPUT75), .B(KEYINPUT84), .Z(n466) );
  OR2_X1 U559 ( .A1(G237), .A2(G902), .ZN(n474) );
  NAND2_X1 U560 ( .A1(G210), .A2(n474), .ZN(n472) );
  NAND2_X1 U561 ( .A1(G214), .A2(n474), .ZN(n680) );
  NAND2_X1 U562 ( .A1(n564), .A2(n680), .ZN(n475) );
  XNOR2_X1 U563 ( .A(n476), .B(KEYINPUT14), .ZN(n478) );
  NAND2_X1 U564 ( .A1(G902), .A2(n478), .ZN(n547) );
  INV_X1 U565 ( .A(n547), .ZN(n477) );
  NOR2_X1 U566 ( .A1(G898), .A2(n737), .ZN(n720) );
  NAND2_X1 U567 ( .A1(n477), .A2(n720), .ZN(n480) );
  NAND2_X1 U568 ( .A1(G952), .A2(n478), .ZN(n696) );
  NOR2_X1 U569 ( .A1(n696), .A2(G953), .ZN(n479) );
  XNOR2_X1 U570 ( .A(n479), .B(KEYINPUT85), .ZN(n550) );
  NAND2_X1 U571 ( .A1(n480), .A2(n550), .ZN(n481) );
  NAND2_X1 U572 ( .A1(n556), .A2(n481), .ZN(n483) );
  XNOR2_X1 U573 ( .A(KEYINPUT80), .B(KEYINPUT0), .ZN(n482) );
  XNOR2_X1 U574 ( .A(n483), .B(n482), .ZN(n537) );
  INV_X1 U575 ( .A(KEYINPUT34), .ZN(n484) );
  XNOR2_X1 U576 ( .A(G116), .B(n485), .ZN(n486) );
  XNOR2_X1 U577 ( .A(n486), .B(KEYINPUT98), .ZN(n492) );
  NAND2_X1 U578 ( .A1(G217), .A2(n487), .ZN(n490) );
  XOR2_X1 U579 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n489) );
  XNOR2_X1 U580 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n488) );
  XNOR2_X1 U581 ( .A(n494), .B(n493), .ZN(n715) );
  NAND2_X1 U582 ( .A1(n715), .A2(n495), .ZN(n498) );
  INV_X1 U583 ( .A(KEYINPUT101), .ZN(n496) );
  XNOR2_X1 U584 ( .A(n496), .B(G478), .ZN(n497) );
  XNOR2_X1 U585 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n512) );
  NAND2_X1 U586 ( .A1(G214), .A2(n499), .ZN(n500) );
  XNOR2_X1 U587 ( .A(n501), .B(n500), .ZN(n505) );
  XNOR2_X1 U588 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U589 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U590 ( .A(n506), .B(n730), .ZN(n510) );
  XNOR2_X1 U591 ( .A(G122), .B(n507), .ZN(n508) );
  XOR2_X1 U592 ( .A(n508), .B(G140), .Z(n509) );
  XNOR2_X1 U593 ( .A(n510), .B(n509), .ZN(n633) );
  NOR2_X1 U594 ( .A1(n633), .A2(G902), .ZN(n511) );
  AND2_X1 U595 ( .A1(n534), .A2(n532), .ZN(n574) );
  XNOR2_X1 U596 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n513) );
  INV_X1 U597 ( .A(n537), .ZN(n517) );
  NOR2_X1 U598 ( .A1(n532), .A2(n534), .ZN(n514) );
  XNOR2_X1 U599 ( .A(n514), .B(KEYINPUT103), .ZN(n684) );
  NOR2_X1 U600 ( .A1(n684), .A2(n515), .ZN(n516) );
  NAND2_X1 U601 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U602 ( .A(KEYINPUT22), .B(n518), .ZN(n523) );
  XNOR2_X1 U603 ( .A(n519), .B(KEYINPUT82), .ZN(n582) );
  NAND2_X1 U604 ( .A1(n579), .A2(n524), .ZN(n520) );
  OR2_X1 U605 ( .A1(n582), .A2(n520), .ZN(n521) );
  NOR2_X1 U606 ( .A1(n523), .A2(n521), .ZN(n522) );
  XNOR2_X1 U607 ( .A(n522), .B(KEYINPUT32), .ZN(n745) );
  INV_X1 U608 ( .A(n523), .ZN(n531) );
  AND2_X1 U609 ( .A1(n671), .A2(n524), .ZN(n525) );
  AND2_X1 U610 ( .A1(n519), .A2(n525), .ZN(n526) );
  NAND2_X1 U611 ( .A1(n531), .A2(n526), .ZN(n647) );
  INV_X1 U612 ( .A(n647), .ZN(n527) );
  AND2_X1 U613 ( .A1(n519), .A2(n666), .ZN(n529) );
  AND2_X1 U614 ( .A1(n529), .A2(n579), .ZN(n530) );
  NAND2_X1 U615 ( .A1(n531), .A2(n530), .ZN(n639) );
  XNOR2_X1 U616 ( .A(KEYINPUT97), .B(n532), .ZN(n533) );
  INV_X1 U617 ( .A(n577), .ZN(n594) );
  NAND2_X1 U618 ( .A1(n600), .A2(n594), .ZN(n685) );
  XOR2_X1 U619 ( .A(KEYINPUT76), .B(n685), .Z(n560) );
  INV_X1 U620 ( .A(n671), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n535), .A2(n565), .ZN(n664) );
  OR2_X1 U622 ( .A1(n537), .A2(n664), .ZN(n536) );
  XNOR2_X1 U623 ( .A(n536), .B(KEYINPUT31), .ZN(n655) );
  BUF_X1 U624 ( .A(n538), .Z(n539) );
  NOR2_X1 U625 ( .A1(n539), .A2(n669), .ZN(n540) );
  NAND2_X1 U626 ( .A1(n517), .A2(n540), .ZN(n541) );
  NOR2_X1 U627 ( .A1(n565), .A2(n541), .ZN(n642) );
  NOR2_X1 U628 ( .A1(n655), .A2(n642), .ZN(n542) );
  NAND2_X1 U629 ( .A1(n639), .A2(n353), .ZN(n544) );
  INV_X1 U630 ( .A(KEYINPUT104), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n544), .B(n543), .ZN(n545) );
  INV_X1 U632 ( .A(KEYINPUT45), .ZN(n546) );
  NOR2_X1 U633 ( .A1(G900), .A2(n547), .ZN(n548) );
  NAND2_X1 U634 ( .A1(G953), .A2(n548), .ZN(n549) );
  NAND2_X1 U635 ( .A1(n550), .A2(n549), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n665), .A2(n569), .ZN(n551) );
  NOR2_X1 U637 ( .A1(n666), .A2(n551), .ZN(n552) );
  XNOR2_X1 U638 ( .A(n552), .B(KEYINPUT66), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n576), .A2(n565), .ZN(n555) );
  INV_X1 U640 ( .A(n539), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n556), .A2(n586), .ZN(n557) );
  NOR2_X1 U642 ( .A1(n585), .A2(n557), .ZN(n651) );
  NAND2_X1 U643 ( .A1(n685), .A2(n651), .ZN(n558) );
  NAND2_X1 U644 ( .A1(n558), .A2(KEYINPUT47), .ZN(n563) );
  XOR2_X1 U645 ( .A(KEYINPUT65), .B(KEYINPUT47), .Z(n559) );
  NOR2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U647 ( .A1(n561), .A2(n651), .ZN(n562) );
  INV_X1 U648 ( .A(n564), .ZN(n605) );
  NAND2_X1 U649 ( .A1(n565), .A2(n680), .ZN(n568) );
  XOR2_X1 U650 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n566) );
  INV_X1 U651 ( .A(n569), .ZN(n570) );
  NOR2_X1 U652 ( .A1(n669), .A2(n570), .ZN(n571) );
  NAND2_X1 U653 ( .A1(n586), .A2(n571), .ZN(n572) );
  NOR2_X1 U654 ( .A1(n573), .A2(n572), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n591), .A2(n574), .ZN(n575) );
  NOR2_X1 U656 ( .A1(n605), .A2(n575), .ZN(n650) );
  NAND2_X1 U657 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U659 ( .A1(n580), .A2(n680), .ZN(n602) );
  XOR2_X1 U660 ( .A(KEYINPUT36), .B(n581), .Z(n583) );
  NOR2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n658) );
  INV_X1 U662 ( .A(n585), .ZN(n587) );
  XOR2_X1 U663 ( .A(KEYINPUT69), .B(KEYINPUT38), .Z(n588) );
  XOR2_X1 U664 ( .A(KEYINPUT42), .B(n590), .Z(n744) );
  NAND2_X1 U665 ( .A1(n591), .A2(n681), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n601), .ZN(n595) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT40), .ZN(n743) );
  NOR2_X1 U668 ( .A1(n744), .A2(n743), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n596), .B(KEYINPUT46), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n660) );
  NOR2_X1 U671 ( .A1(n602), .A2(n379), .ZN(n604) );
  XOR2_X1 U672 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n603) );
  XNOR2_X1 U673 ( .A(n604), .B(n603), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n661) );
  INV_X1 U675 ( .A(n661), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n660), .A2(n607), .ZN(n608) );
  AND2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n610) );
  INV_X1 U678 ( .A(KEYINPUT64), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n713), .A2(G210), .ZN(n619) );
  XOR2_X1 U680 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n615) );
  XNOR2_X1 U681 ( .A(KEYINPUT79), .B(KEYINPUT55), .ZN(n614) );
  XNOR2_X1 U682 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U683 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U684 ( .A(n619), .B(n618), .ZN(n623) );
  INV_X1 U685 ( .A(G952), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n620), .A2(G953), .ZN(n622) );
  INV_X1 U687 ( .A(KEYINPUT83), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n622), .B(n621), .ZN(n634) );
  NAND2_X1 U689 ( .A1(n623), .A2(n634), .ZN(n625) );
  INV_X1 U690 ( .A(KEYINPUT56), .ZN(n624) );
  XNOR2_X1 U691 ( .A(n625), .B(n624), .ZN(G51) );
  NAND2_X1 U692 ( .A1(n713), .A2(G472), .ZN(n629) );
  XNOR2_X1 U693 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n627) );
  XNOR2_X1 U694 ( .A(n626), .B(n627), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U696 ( .A1(n630), .A2(n634), .ZN(n631) );
  XNOR2_X1 U697 ( .A(n631), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U698 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n632) );
  INV_X1 U699 ( .A(n634), .ZN(n717) );
  XOR2_X1 U700 ( .A(n635), .B(G122), .Z(G24) );
  NAND2_X1 U701 ( .A1(n713), .A2(G217), .ZN(n637) );
  XNOR2_X1 U702 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U703 ( .A1(n638), .A2(n717), .ZN(G66) );
  XOR2_X1 U704 ( .A(G101), .B(n639), .Z(n640) );
  XNOR2_X1 U705 ( .A(n640), .B(KEYINPUT111), .ZN(G3) );
  NAND2_X1 U706 ( .A1(n642), .A2(n577), .ZN(n641) );
  XNOR2_X1 U707 ( .A(n641), .B(G104), .ZN(G6) );
  XNOR2_X1 U708 ( .A(G107), .B(KEYINPUT26), .ZN(n646) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n644) );
  NAND2_X1 U710 ( .A1(n642), .A2(n654), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U712 ( .A(n646), .B(n645), .ZN(G9) );
  XNOR2_X1 U713 ( .A(n647), .B(G110), .ZN(G12) );
  XOR2_X1 U714 ( .A(G128), .B(KEYINPUT29), .Z(n649) );
  NAND2_X1 U715 ( .A1(n651), .A2(n654), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n650), .Z(G45) );
  NAND2_X1 U718 ( .A1(n651), .A2(n577), .ZN(n652) );
  XNOR2_X1 U719 ( .A(n652), .B(G146), .ZN(G48) );
  NAND2_X1 U720 ( .A1(n655), .A2(n577), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n653), .B(G113), .ZN(G15) );
  XOR2_X1 U722 ( .A(G116), .B(KEYINPUT113), .Z(n657) );
  NAND2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n657), .B(n656), .ZN(G18) );
  XNOR2_X1 U725 ( .A(G125), .B(n658), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n659), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U727 ( .A(G134), .B(n660), .Z(G36) );
  XNOR2_X1 U728 ( .A(G140), .B(KEYINPUT114), .ZN(n662) );
  XNOR2_X1 U729 ( .A(n662), .B(n661), .ZN(G42) );
  NAND2_X1 U730 ( .A1(n721), .A2(n610), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(KEYINPUT2), .ZN(n703) );
  INV_X1 U732 ( .A(n664), .ZN(n676) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n668) );
  XNOR2_X1 U734 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n674) );
  NAND2_X1 U736 ( .A1(n519), .A2(n669), .ZN(n670) );
  XNOR2_X1 U737 ( .A(KEYINPUT50), .B(n670), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U741 ( .A(KEYINPUT51), .B(n677), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n678), .A2(n697), .ZN(n679) );
  XOR2_X1 U743 ( .A(KEYINPUT116), .B(n679), .Z(n693) );
  NOR2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT117), .B(n682), .Z(n683) );
  NOR2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n690) );
  INV_X1 U747 ( .A(n685), .ZN(n687) );
  NOR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT118), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n405), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n694), .B(KEYINPUT52), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n701) );
  INV_X1 U754 ( .A(n697), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n699), .A2(n698), .ZN(n700) );
  OR2_X1 U756 ( .A1(n701), .A2(n700), .ZN(n702) );
  OR2_X2 U757 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U758 ( .A(KEYINPUT119), .B(n704), .Z(n705) );
  NOR2_X2 U759 ( .A1(G953), .A2(n705), .ZN(n706) );
  XNOR2_X1 U760 ( .A(KEYINPUT53), .B(n706), .ZN(G75) );
  NAND2_X1 U761 ( .A1(n713), .A2(G469), .ZN(n711) );
  XOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n707) );
  XNOR2_X1 U763 ( .A(n707), .B(KEYINPUT121), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n717), .A2(n712), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n713), .A2(G478), .ZN(n714) );
  XOR2_X1 U768 ( .A(n715), .B(n714), .Z(n716) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(G63) );
  XNOR2_X1 U770 ( .A(n718), .B(G110), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n728) );
  NAND2_X1 U772 ( .A1(n721), .A2(n737), .ZN(n726) );
  XOR2_X1 U773 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n723) );
  NAND2_X1 U774 ( .A1(G224), .A2(G953), .ZN(n722) );
  XNOR2_X1 U775 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(G69) );
  XNOR2_X1 U779 ( .A(n729), .B(KEYINPUT124), .ZN(n731) );
  XNOR2_X1 U780 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(n736) );
  XOR2_X1 U782 ( .A(G227), .B(n736), .Z(n734) );
  NOR2_X1 U783 ( .A1(n737), .A2(n734), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(G900), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n610), .B(n736), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n741), .ZN(G72) );
  XOR2_X1 U789 ( .A(G131), .B(KEYINPUT126), .Z(n742) );
  XNOR2_X1 U790 ( .A(n743), .B(n742), .ZN(G33) );
  XOR2_X1 U791 ( .A(n744), .B(G137), .Z(G39) );
  XOR2_X1 U792 ( .A(G119), .B(n745), .Z(G21) );
endmodule

