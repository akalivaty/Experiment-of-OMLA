

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755;

  XNOR2_X1 U365 ( .A(n554), .B(n553), .ZN(n561) );
  XNOR2_X1 U366 ( .A(n461), .B(KEYINPUT41), .ZN(n703) );
  OR2_X1 U367 ( .A1(n641), .A2(n452), .ZN(n456) );
  XNOR2_X1 U368 ( .A(n343), .B(n439), .ZN(n727) );
  XNOR2_X1 U369 ( .A(n462), .B(n347), .ZN(n463) );
  XNOR2_X1 U370 ( .A(n472), .B(n437), .ZN(n343) );
  XNOR2_X2 U371 ( .A(n344), .B(n613), .ZN(n706) );
  NOR2_X2 U372 ( .A1(n707), .A2(n612), .ZN(n344) );
  NOR2_X2 U373 ( .A1(n621), .A2(n725), .ZN(n623) );
  NOR2_X2 U374 ( .A1(n629), .A2(n725), .ZN(n630) );
  AND2_X2 U375 ( .A1(n345), .A2(n552), .ZN(n554) );
  XNOR2_X1 U376 ( .A(n384), .B(KEYINPUT46), .ZN(n345) );
  NAND2_X1 U377 ( .A1(n703), .A2(n530), .ZN(n510) );
  INV_X2 U378 ( .A(G953), .ZN(n744) );
  AND2_X1 U379 ( .A1(n755), .A2(n587), .ZN(n346) );
  XNOR2_X2 U380 ( .A(n441), .B(n418), .ZN(n464) );
  OR2_X2 U381 ( .A1(n617), .A2(G902), .ZN(n401) );
  XNOR2_X2 U382 ( .A(n507), .B(n506), .ZN(n624) );
  AND2_X1 U383 ( .A1(n718), .A2(G472), .ZN(n635) );
  AND2_X1 U384 ( .A1(n718), .A2(G210), .ZN(n643) );
  INV_X1 U385 ( .A(n702), .ZN(n392) );
  INV_X1 U386 ( .A(n517), .ZN(n670) );
  INV_X1 U387 ( .A(G125), .ZN(n396) );
  INV_X2 U388 ( .A(G143), .ZN(n417) );
  NAND2_X1 U389 ( .A1(n365), .A2(n361), .ZN(n755) );
  NAND2_X1 U390 ( .A1(n364), .A2(n362), .ZN(n361) );
  NAND2_X1 U391 ( .A1(n379), .A2(n377), .ZN(n590) );
  AND2_X1 U392 ( .A1(n381), .A2(n349), .ZN(n379) );
  NAND2_X1 U393 ( .A1(n378), .A2(KEYINPUT108), .ZN(n377) );
  OR2_X1 U394 ( .A1(n599), .A2(n572), .ZN(n393) );
  XNOR2_X1 U395 ( .A(n382), .B(n351), .ZN(n568) );
  AND2_X1 U396 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U397 ( .A(n396), .B(G146), .ZN(n442) );
  XNOR2_X1 U398 ( .A(n435), .B(n434), .ZN(n472) );
  XNOR2_X1 U399 ( .A(KEYINPUT69), .B(G107), .ZN(n503) );
  XNOR2_X1 U400 ( .A(KEYINPUT3), .B(G116), .ZN(n434) );
  XNOR2_X1 U401 ( .A(G113), .B(G101), .ZN(n435) );
  NOR2_X1 U402 ( .A1(n593), .A2(n602), .ZN(n564) );
  NOR2_X1 U403 ( .A1(n754), .A2(n753), .ZN(n384) );
  NAND2_X1 U404 ( .A1(n624), .A2(n390), .ZN(n376) );
  XNOR2_X1 U405 ( .A(n571), .B(n570), .ZN(n576) );
  INV_X1 U406 ( .A(KEYINPUT44), .ZN(n358) );
  INV_X1 U407 ( .A(n631), .ZN(n354) );
  NOR2_X1 U408 ( .A1(n631), .A2(n358), .ZN(n356) );
  XNOR2_X1 U409 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n436) );
  INV_X1 U410 ( .A(G134), .ZN(n418) );
  INV_X1 U411 ( .A(KEYINPUT11), .ZN(n413) );
  XOR2_X1 U412 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n404) );
  NAND2_X2 U413 ( .A1(n374), .A2(n371), .ZN(n516) );
  OR2_X1 U414 ( .A1(n624), .A2(n372), .ZN(n371) );
  NAND2_X1 U415 ( .A1(G469), .A2(n373), .ZN(n372) );
  XNOR2_X1 U416 ( .A(n395), .B(n412), .ZN(n740) );
  XNOR2_X1 U417 ( .A(n442), .B(G140), .ZN(n395) );
  XNOR2_X1 U418 ( .A(n387), .B(n386), .ZN(n555) );
  INV_X1 U419 ( .A(KEYINPUT39), .ZN(n386) );
  NAND2_X1 U420 ( .A1(n388), .A2(n537), .ZN(n387) );
  AND2_X1 U421 ( .A1(n512), .A2(n536), .ZN(n388) );
  NOR2_X1 U422 ( .A1(n522), .A2(n687), .ZN(n557) );
  NAND2_X1 U423 ( .A1(n370), .A2(n348), .ZN(n368) );
  AND2_X1 U424 ( .A1(n363), .A2(n575), .ZN(n362) );
  NAND2_X1 U425 ( .A1(n392), .A2(n391), .ZN(n363) );
  INV_X1 U426 ( .A(KEYINPUT107), .ZN(n581) );
  XNOR2_X1 U427 ( .A(n416), .B(n400), .ZN(n399) );
  INV_X1 U428 ( .A(G475), .ZN(n400) );
  INV_X1 U429 ( .A(KEYINPUT22), .ZN(n397) );
  XOR2_X1 U430 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n406) );
  XNOR2_X1 U431 ( .A(G131), .B(G113), .ZN(n405) );
  NAND2_X1 U432 ( .A1(n390), .A2(G902), .ZN(n375) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n468) );
  NAND2_X1 U434 ( .A1(n346), .A2(n356), .ZN(n355) );
  INV_X1 U435 ( .A(n572), .ZN(n391) );
  XNOR2_X1 U436 ( .A(n511), .B(KEYINPUT30), .ZN(n537) );
  NOR2_X1 U437 ( .A1(G902), .A2(G237), .ZN(n454) );
  XNOR2_X1 U438 ( .A(n433), .B(n432), .ZN(n690) );
  XNOR2_X1 U439 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n483) );
  XNOR2_X1 U440 ( .A(G128), .B(G137), .ZN(n486) );
  XNOR2_X1 U441 ( .A(n414), .B(n415), .ZN(n617) );
  INV_X1 U442 ( .A(G146), .ZN(n465) );
  XNOR2_X1 U443 ( .A(G101), .B(G110), .ZN(n500) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n477) );
  OR2_X1 U445 ( .A1(n517), .A2(n589), .ZN(n380) );
  AND2_X1 U446 ( .A1(n620), .A2(G953), .ZN(n725) );
  XNOR2_X1 U447 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U448 ( .A(n515), .B(n385), .ZN(n753) );
  XNOR2_X1 U449 ( .A(KEYINPUT36), .B(KEYINPUT112), .ZN(n523) );
  AND2_X1 U450 ( .A1(n367), .A2(n366), .ZN(n365) );
  INV_X1 U451 ( .A(n368), .ZN(n364) );
  XNOR2_X1 U452 ( .A(n586), .B(n585), .ZN(n752) );
  XNOR2_X1 U453 ( .A(n531), .B(KEYINPUT104), .ZN(n653) );
  XOR2_X1 U454 ( .A(KEYINPUT4), .B(G137), .Z(n347) );
  AND2_X1 U455 ( .A1(n393), .A2(n574), .ZN(n348) );
  INV_X1 U456 ( .A(G469), .ZN(n390) );
  AND2_X1 U457 ( .A1(n380), .A2(n592), .ZN(n349) );
  AND2_X1 U458 ( .A1(n517), .A2(n589), .ZN(n350) );
  XOR2_X1 U459 ( .A(n529), .B(n528), .Z(n351) );
  INV_X1 U460 ( .A(G902), .ZN(n373) );
  AND2_X1 U461 ( .A1(n391), .A2(n369), .ZN(n352) );
  INV_X1 U462 ( .A(KEYINPUT108), .ZN(n589) );
  AND2_X1 U463 ( .A1(n583), .A2(n602), .ZN(n398) );
  NAND2_X1 U464 ( .A1(n353), .A2(n358), .ZN(n357) );
  NAND2_X1 U465 ( .A1(n346), .A2(n354), .ZN(n353) );
  NAND2_X1 U466 ( .A1(n357), .A2(n355), .ZN(n360) );
  XNOR2_X2 U467 ( .A(n359), .B(n607), .ZN(n707) );
  NAND2_X1 U468 ( .A1(n360), .A2(n606), .ZN(n359) );
  NAND2_X1 U469 ( .A1(n392), .A2(n352), .ZN(n366) );
  NAND2_X1 U470 ( .A1(n368), .A2(n369), .ZN(n367) );
  INV_X1 U471 ( .A(n575), .ZN(n369) );
  NAND2_X1 U472 ( .A1(n394), .A2(n702), .ZN(n370) );
  XNOR2_X2 U473 ( .A(n564), .B(n563), .ZN(n702) );
  XNOR2_X2 U474 ( .A(n516), .B(KEYINPUT1), .ZN(n517) );
  AND2_X2 U475 ( .A1(n615), .A2(n706), .ZN(n718) );
  NAND2_X1 U476 ( .A1(n588), .A2(n517), .ZN(n604) );
  INV_X1 U477 ( .A(n588), .ZN(n378) );
  NAND2_X1 U478 ( .A1(n588), .A2(n350), .ZN(n381) );
  XNOR2_X2 U479 ( .A(n578), .B(n397), .ZN(n588) );
  NAND2_X1 U480 ( .A1(n568), .A2(n402), .ZN(n571) );
  NAND2_X1 U481 ( .A1(n527), .A2(n526), .ZN(n382) );
  XNOR2_X1 U482 ( .A(n590), .B(KEYINPUT64), .ZN(n591) );
  XNOR2_X2 U483 ( .A(G119), .B(G110), .ZN(n485) );
  INV_X1 U484 ( .A(KEYINPUT40), .ZN(n385) );
  NAND2_X1 U485 ( .A1(n669), .A2(n389), .ZN(n597) );
  INV_X1 U486 ( .A(n516), .ZN(n389) );
  XNOR2_X2 U487 ( .A(n741), .B(n465), .ZN(n507) );
  AND2_X1 U488 ( .A1(n599), .A2(n572), .ZN(n394) );
  NAND2_X1 U489 ( .A1(n398), .A2(n588), .ZN(n586) );
  XNOR2_X2 U490 ( .A(n401), .B(n399), .ZN(n540) );
  AND2_X1 U491 ( .A1(n567), .A2(n698), .ZN(n402) );
  INV_X1 U492 ( .A(KEYINPUT47), .ZN(n533) );
  XNOR2_X1 U493 ( .A(n534), .B(n533), .ZN(n547) );
  INV_X1 U494 ( .A(KEYINPUT73), .ZN(n548) );
  INV_X1 U495 ( .A(KEYINPUT45), .ZN(n607) );
  AND2_X1 U496 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U497 ( .A(KEYINPUT48), .ZN(n553) );
  INV_X1 U498 ( .A(KEYINPUT78), .ZN(n613) );
  INV_X1 U499 ( .A(n573), .ZN(n574) );
  BUF_X1 U500 ( .A(n709), .Z(n743) );
  BUF_X1 U501 ( .A(n576), .Z(n599) );
  XNOR2_X1 U502 ( .A(n510), .B(n509), .ZN(n754) );
  XNOR2_X1 U503 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n416) );
  NAND2_X1 U504 ( .A1(G214), .A2(n468), .ZN(n403) );
  XNOR2_X1 U505 ( .A(n404), .B(n403), .ZN(n408) );
  XNOR2_X1 U506 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U507 ( .A(n408), .B(n407), .ZN(n411) );
  INV_X1 U508 ( .A(G122), .ZN(n409) );
  XNOR2_X1 U509 ( .A(n409), .B(G104), .ZN(n438) );
  XNOR2_X1 U510 ( .A(n438), .B(G143), .ZN(n410) );
  XNOR2_X1 U511 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U512 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n412) );
  XNOR2_X1 U513 ( .A(n740), .B(n413), .ZN(n414) );
  XNOR2_X1 U514 ( .A(KEYINPUT103), .B(G478), .ZN(n430) );
  XNOR2_X2 U515 ( .A(n417), .B(G128), .ZN(n441) );
  INV_X1 U516 ( .A(n464), .ZN(n422) );
  XOR2_X1 U517 ( .A(KEYINPUT102), .B(G107), .Z(n420) );
  XNOR2_X1 U518 ( .A(G116), .B(G122), .ZN(n419) );
  XNOR2_X1 U519 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U520 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U521 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n426) );
  XOR2_X1 U522 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n424) );
  NAND2_X1 U523 ( .A1(G234), .A2(n744), .ZN(n423) );
  XNOR2_X1 U524 ( .A(n424), .B(n423), .ZN(n489) );
  NAND2_X1 U525 ( .A1(G217), .A2(n489), .ZN(n425) );
  XNOR2_X1 U526 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U527 ( .A(n428), .B(n427), .ZN(n719) );
  NOR2_X1 U528 ( .A1(G902), .A2(n719), .ZN(n429) );
  XNOR2_X1 U529 ( .A(n430), .B(n429), .ZN(n542) );
  INV_X1 U530 ( .A(n542), .ZN(n431) );
  NAND2_X1 U531 ( .A1(n540), .A2(n431), .ZN(n433) );
  INV_X1 U532 ( .A(KEYINPUT106), .ZN(n432) );
  XNOR2_X1 U533 ( .A(n436), .B(KEYINPUT16), .ZN(n437) );
  XNOR2_X1 U534 ( .A(n438), .B(n485), .ZN(n439) );
  XNOR2_X1 U535 ( .A(n442), .B(n441), .ZN(n445) );
  XNOR2_X1 U536 ( .A(KEYINPUT4), .B(KEYINPUT90), .ZN(n443) );
  XNOR2_X1 U537 ( .A(n503), .B(n443), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n445), .B(n444), .ZN(n450) );
  XOR2_X1 U539 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n448) );
  NAND2_X1 U540 ( .A1(G224), .A2(n744), .ZN(n446) );
  XNOR2_X1 U541 ( .A(n446), .B(KEYINPUT88), .ZN(n447) );
  XNOR2_X1 U542 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U543 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U544 ( .A(n727), .B(n451), .ZN(n641) );
  XNOR2_X1 U545 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  INV_X1 U546 ( .A(n610), .ZN(n452) );
  INV_X1 U547 ( .A(KEYINPUT75), .ZN(n453) );
  XNOR2_X1 U548 ( .A(n454), .B(n453), .ZN(n458) );
  INV_X1 U549 ( .A(G210), .ZN(n639) );
  NOR2_X1 U550 ( .A1(n458), .A2(n639), .ZN(n455) );
  XNOR2_X2 U551 ( .A(n456), .B(n455), .ZN(n527) );
  XNOR2_X1 U552 ( .A(n527), .B(KEYINPUT38), .ZN(n688) );
  INV_X1 U553 ( .A(G214), .ZN(n457) );
  OR2_X1 U554 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U555 ( .A(n459), .B(KEYINPUT91), .ZN(n687) );
  NOR2_X1 U556 ( .A1(n688), .A2(n687), .ZN(n460) );
  XNOR2_X1 U557 ( .A(n460), .B(KEYINPUT110), .ZN(n684) );
  NAND2_X1 U558 ( .A1(n690), .A2(n684), .ZN(n461) );
  XOR2_X1 U559 ( .A(KEYINPUT67), .B(G131), .Z(n462) );
  XNOR2_X2 U560 ( .A(n464), .B(n463), .ZN(n741) );
  XOR2_X1 U561 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n467) );
  XNOR2_X1 U562 ( .A(G119), .B(KEYINPUT96), .ZN(n466) );
  XNOR2_X1 U563 ( .A(n467), .B(n466), .ZN(n470) );
  NAND2_X1 U564 ( .A1(n468), .A2(G210), .ZN(n469) );
  XNOR2_X1 U565 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U566 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U567 ( .A(n507), .B(n473), .ZN(n633) );
  NAND2_X1 U568 ( .A1(n633), .A2(n373), .ZN(n474) );
  INV_X1 U569 ( .A(G472), .ZN(n632) );
  XNOR2_X2 U570 ( .A(n474), .B(n632), .ZN(n592) );
  INV_X1 U571 ( .A(n592), .ZN(n677) );
  NOR2_X1 U572 ( .A1(G900), .A2(n744), .ZN(n475) );
  NAND2_X1 U573 ( .A1(n475), .A2(G902), .ZN(n476) );
  NAND2_X1 U574 ( .A1(G952), .A2(n744), .ZN(n565) );
  NAND2_X1 U575 ( .A1(n476), .A2(n565), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n477), .B(KEYINPUT14), .ZN(n698) );
  NAND2_X1 U577 ( .A1(n478), .A2(n698), .ZN(n535) );
  NAND2_X1 U578 ( .A1(G234), .A2(n610), .ZN(n479) );
  XNOR2_X1 U579 ( .A(KEYINPUT20), .B(n479), .ZN(n493) );
  AND2_X1 U580 ( .A1(n493), .A2(G221), .ZN(n482) );
  INV_X1 U581 ( .A(KEYINPUT95), .ZN(n480) );
  XNOR2_X1 U582 ( .A(n480), .B(KEYINPUT21), .ZN(n481) );
  XNOR2_X1 U583 ( .A(n482), .B(n481), .ZN(n673) );
  XOR2_X1 U584 ( .A(KEYINPUT24), .B(KEYINPUT68), .Z(n484) );
  XNOR2_X1 U585 ( .A(n484), .B(n483), .ZN(n488) );
  XNOR2_X1 U586 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U587 ( .A(n488), .B(n487), .ZN(n491) );
  NAND2_X1 U588 ( .A1(n489), .A2(G221), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U590 ( .A(n740), .B(n492), .ZN(n722) );
  NOR2_X1 U591 ( .A1(n722), .A2(G902), .ZN(n497) );
  XOR2_X1 U592 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n495) );
  NAND2_X1 U593 ( .A1(G217), .A2(n493), .ZN(n494) );
  XNOR2_X1 U594 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U595 ( .A(n497), .B(n496), .ZN(n579) );
  NAND2_X1 U596 ( .A1(n673), .A2(n579), .ZN(n498) );
  NOR2_X1 U597 ( .A1(n535), .A2(n498), .ZN(n519) );
  NAND2_X1 U598 ( .A1(n677), .A2(n519), .ZN(n499) );
  XNOR2_X1 U599 ( .A(KEYINPUT28), .B(n499), .ZN(n508) );
  XOR2_X1 U600 ( .A(G140), .B(G104), .Z(n501) );
  XNOR2_X1 U601 ( .A(n501), .B(n500), .ZN(n505) );
  NAND2_X1 U602 ( .A1(G227), .A2(n744), .ZN(n502) );
  XOR2_X1 U603 ( .A(n503), .B(n502), .Z(n504) );
  XNOR2_X1 U604 ( .A(n505), .B(n504), .ZN(n506) );
  NOR2_X1 U605 ( .A1(n508), .A2(n516), .ZN(n530) );
  NOR2_X1 U606 ( .A1(n687), .A2(n592), .ZN(n511) );
  NOR2_X1 U607 ( .A1(n688), .A2(n535), .ZN(n512) );
  INV_X1 U608 ( .A(n673), .ZN(n513) );
  NOR2_X1 U609 ( .A1(n513), .A2(n579), .ZN(n669) );
  INV_X1 U610 ( .A(n555), .ZN(n514) );
  NOR2_X2 U611 ( .A1(n542), .A2(n540), .ZN(n660) );
  NAND2_X1 U612 ( .A1(n514), .A2(n660), .ZN(n515) );
  XOR2_X1 U613 ( .A(KEYINPUT89), .B(n517), .Z(n580) );
  INV_X1 U614 ( .A(KEYINPUT6), .ZN(n518) );
  XNOR2_X1 U615 ( .A(n592), .B(n518), .ZN(n602) );
  NAND2_X1 U616 ( .A1(n660), .A2(n519), .ZN(n520) );
  NOR2_X1 U617 ( .A1(n602), .A2(n520), .ZN(n521) );
  XNOR2_X1 U618 ( .A(n521), .B(KEYINPUT109), .ZN(n522) );
  NAND2_X1 U619 ( .A1(n557), .A2(n527), .ZN(n524) );
  XNOR2_X1 U620 ( .A(n524), .B(n523), .ZN(n525) );
  NOR2_X1 U621 ( .A1(n580), .A2(n525), .ZN(n665) );
  INV_X1 U622 ( .A(n665), .ZN(n551) );
  INV_X1 U623 ( .A(n687), .ZN(n526) );
  XNOR2_X1 U624 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n529) );
  INV_X1 U625 ( .A(KEYINPUT65), .ZN(n528) );
  NAND2_X1 U626 ( .A1(n530), .A2(n568), .ZN(n658) );
  INV_X1 U627 ( .A(n660), .ZN(n657) );
  NAND2_X1 U628 ( .A1(n540), .A2(n542), .ZN(n531) );
  NAND2_X1 U629 ( .A1(n657), .A2(n653), .ZN(n685) );
  INV_X1 U630 ( .A(n685), .ZN(n532) );
  NOR2_X1 U631 ( .A1(n658), .A2(n532), .ZN(n534) );
  INV_X1 U632 ( .A(n535), .ZN(n539) );
  INV_X1 U633 ( .A(n597), .ZN(n536) );
  AND2_X1 U634 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U635 ( .A1(n539), .A2(n538), .ZN(n545) );
  INV_X1 U636 ( .A(n527), .ZN(n543) );
  INV_X1 U637 ( .A(n540), .ZN(n541) );
  NAND2_X1 U638 ( .A1(n542), .A2(n541), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n543), .A2(n573), .ZN(n544) );
  AND2_X1 U640 ( .A1(n545), .A2(n544), .ZN(n656) );
  XOR2_X1 U641 ( .A(KEYINPUT81), .B(n656), .Z(n546) );
  NOR2_X1 U642 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X1 U643 ( .A(n549), .B(n548), .ZN(n550) );
  NOR2_X1 U644 ( .A1(n555), .A2(n653), .ZN(n556) );
  XNOR2_X1 U645 ( .A(n556), .B(KEYINPUT113), .ZN(n751) );
  NAND2_X1 U646 ( .A1(n517), .A2(n557), .ZN(n558) );
  XOR2_X1 U647 ( .A(KEYINPUT43), .B(n558), .Z(n559) );
  OR2_X1 U648 ( .A1(n559), .A2(n527), .ZN(n667) );
  NAND2_X1 U649 ( .A1(n751), .A2(n667), .ZN(n560) );
  NOR2_X2 U650 ( .A1(n561), .A2(n560), .ZN(n709) );
  XNOR2_X1 U651 ( .A(n709), .B(KEYINPUT77), .ZN(n608) );
  NAND2_X1 U652 ( .A1(n669), .A2(n670), .ZN(n562) );
  XNOR2_X1 U653 ( .A(n562), .B(KEYINPUT74), .ZN(n593) );
  XNOR2_X1 U654 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n563) );
  XNOR2_X1 U655 ( .A(G898), .B(KEYINPUT92), .ZN(n733) );
  NOR2_X1 U656 ( .A1(n744), .A2(n733), .ZN(n728) );
  NAND2_X1 U657 ( .A1(n728), .A2(G902), .ZN(n566) );
  NAND2_X1 U658 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U659 ( .A(KEYINPUT86), .ZN(n569) );
  XNOR2_X1 U660 ( .A(n569), .B(KEYINPUT0), .ZN(n570) );
  XOR2_X1 U661 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n572) );
  XNOR2_X1 U662 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n575) );
  AND2_X1 U663 ( .A1(n690), .A2(n673), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n578) );
  INV_X1 U665 ( .A(n579), .ZN(n674) );
  NOR2_X1 U666 ( .A1(n674), .A2(n580), .ZN(n582) );
  XNOR2_X1 U667 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U668 ( .A(KEYINPUT80), .ZN(n584) );
  XNOR2_X1 U669 ( .A(n584), .B(KEYINPUT32), .ZN(n585) );
  INV_X1 U670 ( .A(n752), .ZN(n587) );
  NOR2_X2 U671 ( .A1(n591), .A2(n674), .ZN(n631) );
  OR2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n680) );
  INV_X1 U673 ( .A(n599), .ZN(n594) );
  NOR2_X1 U674 ( .A1(n680), .A2(n594), .ZN(n596) );
  XNOR2_X1 U675 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n595) );
  XNOR2_X1 U676 ( .A(n596), .B(n595), .ZN(n662) );
  NOR2_X1 U677 ( .A1(n677), .A2(n597), .ZN(n598) );
  AND2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n649) );
  OR2_X1 U679 ( .A1(n662), .A2(n649), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n600), .A2(n685), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT105), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n602), .A2(n674), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n647) );
  NOR2_X1 U684 ( .A1(n605), .A2(n647), .ZN(n606) );
  NOR2_X1 U685 ( .A1(n608), .A2(n707), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n609), .A2(KEYINPUT2), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n709), .A2(KEYINPUT2), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n718), .A2(G475), .ZN(n619) );
  XNOR2_X1 U690 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n619), .B(n618), .ZN(n621) );
  INV_X1 U693 ( .A(G952), .ZN(n620) );
  XNOR2_X1 U694 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(G60) );
  NAND2_X1 U696 ( .A1(n718), .A2(G469), .ZN(n628) );
  XNOR2_X1 U697 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(KEYINPUT58), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n624), .B(n626), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(KEYINPUT120), .ZN(G54) );
  XOR2_X1 U702 ( .A(n631), .B(G110), .Z(G12) );
  XNOR2_X1 U703 ( .A(n633), .B(KEYINPUT62), .ZN(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X1 U705 ( .A1(n636), .A2(n725), .ZN(n638) );
  XNOR2_X1 U706 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n638), .B(n637), .ZN(G57) );
  XNOR2_X1 U708 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U710 ( .A(n643), .B(n642), .ZN(n644) );
  NOR2_X1 U711 ( .A1(n644), .A2(n725), .ZN(n646) );
  XNOR2_X1 U712 ( .A(KEYINPUT118), .B(KEYINPUT56), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n646), .B(n645), .ZN(G51) );
  XOR2_X1 U714 ( .A(G101), .B(n647), .Z(G3) );
  NAND2_X1 U715 ( .A1(n649), .A2(n660), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n648), .B(G104), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n651) );
  INV_X1 U718 ( .A(n653), .ZN(n663) );
  NAND2_X1 U719 ( .A1(n649), .A2(n663), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(G107), .B(n652), .ZN(G9) );
  NOR2_X1 U722 ( .A1(n653), .A2(n658), .ZN(n655) );
  XNOR2_X1 U723 ( .A(G128), .B(KEYINPUT29), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(G30) );
  XOR2_X1 U725 ( .A(G143), .B(n656), .Z(G45) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(G146), .B(n659), .Z(G48) );
  NAND2_X1 U728 ( .A1(n662), .A2(n660), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(G113), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n664), .B(G116), .ZN(G18) );
  XNOR2_X1 U732 ( .A(G125), .B(n665), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U734 ( .A(n667), .B(G140), .ZN(n668) );
  XNOR2_X1 U735 ( .A(KEYINPUT114), .B(n668), .ZN(G42) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT115), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT50), .ZN(n679) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U744 ( .A(KEYINPUT51), .B(n682), .Z(n683) );
  NAND2_X1 U745 ( .A1(n703), .A2(n683), .ZN(n696) );
  NAND2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U747 ( .A(KEYINPUT117), .B(n686), .Z(n693) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U749 ( .A(n689), .B(KEYINPUT116), .ZN(n691) );
  NAND2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n702), .A2(n694), .ZN(n695) );
  NAND2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U754 ( .A(KEYINPUT52), .B(n697), .Z(n700) );
  NAND2_X1 U755 ( .A1(G952), .A2(n698), .ZN(n699) );
  NOR2_X1 U756 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U757 ( .A1(G953), .A2(n701), .ZN(n705) );
  NAND2_X1 U758 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U759 ( .A1(n705), .A2(n704), .ZN(n716) );
  INV_X1 U760 ( .A(n706), .ZN(n714) );
  INV_X1 U761 ( .A(KEYINPUT2), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n707), .A2(n708), .ZN(n712) );
  NOR2_X1 U763 ( .A1(n743), .A2(KEYINPUT2), .ZN(n710) );
  XNOR2_X1 U764 ( .A(KEYINPUT83), .B(n710), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U768 ( .A(KEYINPUT53), .B(n717), .ZN(G75) );
  NAND2_X1 U769 ( .A1(n718), .A2(G478), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n725), .A2(n721), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n718), .A2(G217), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U774 ( .A1(n725), .A2(n724), .ZN(G66) );
  XOR2_X1 U775 ( .A(G107), .B(KEYINPUT125), .Z(n726) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n729) );
  NOR2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n738) );
  INV_X1 U778 ( .A(n707), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n730), .A2(n744), .ZN(n736) );
  XOR2_X1 U780 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n732) );
  NAND2_X1 U781 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U785 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U786 ( .A(KEYINPUT124), .B(n739), .ZN(G69) );
  XOR2_X1 U787 ( .A(n741), .B(n740), .Z(n742) );
  XOR2_X1 U788 ( .A(KEYINPUT126), .B(n742), .Z(n746) );
  XOR2_X1 U789 ( .A(n746), .B(n743), .Z(n745) );
  NAND2_X1 U790 ( .A1(n745), .A2(n744), .ZN(n750) );
  XNOR2_X1 U791 ( .A(G227), .B(n746), .ZN(n747) );
  NAND2_X1 U792 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U793 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U794 ( .A1(n750), .A2(n749), .ZN(G72) );
  XNOR2_X1 U795 ( .A(G134), .B(n751), .ZN(G36) );
  XOR2_X1 U796 ( .A(n752), .B(G119), .Z(G21) );
  XOR2_X1 U797 ( .A(G131), .B(n753), .Z(G33) );
  XOR2_X1 U798 ( .A(G137), .B(n754), .Z(G39) );
  XNOR2_X1 U799 ( .A(G122), .B(n755), .ZN(G24) );
endmodule

