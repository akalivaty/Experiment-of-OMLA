//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G78gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT95), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(KEYINPUT95), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n206), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT21), .ZN(new_n214));
  AND2_X1   g013(.A1(G231gat), .A2(G233gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G127gat), .ZN(new_n219));
  INV_X1    g018(.A(G127gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n220), .A3(new_n217), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT16), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G1gat), .B2(new_n223), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(G8gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(G8gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(KEYINPUT21), .B2(new_n213), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n231), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n219), .A2(new_n233), .A3(new_n221), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n236));
  INV_X1    g035(.A(G155gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G183gat), .B(G211gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(new_n234), .A3(new_n240), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT41), .ZN(new_n247));
  XNOR2_X1  g046(.A(G134gat), .B(G162gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT14), .ZN(new_n251));
  INV_X1    g050(.A(G29gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n254));
  AOI21_X1  g053(.A(G36gat), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G36gat), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n251), .A2(new_n256), .A3(G29gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT15), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  INV_X1    g058(.A(new_n254), .ZN(new_n260));
  NOR2_X1   g059(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n256), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT15), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G43gat), .B(G50gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n267), .B(KEYINPUT15), .C1(new_n255), .C2(new_n257), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT17), .ZN(new_n270));
  NAND2_X1  g069(.A1(G85gat), .A2(G92gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT7), .ZN(new_n272));
  OR2_X1    g071(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n273));
  INV_X1    g072(.A(G92gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G99gat), .ZN(new_n277));
  INV_X1    g076(.A(G106gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT8), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n272), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G99gat), .B(G106gat), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n283), .A2(new_n272), .A3(new_n276), .A4(new_n279), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n287), .A2(new_n269), .B1(KEYINPUT41), .B2(new_n246), .ZN(new_n288));
  XNOR2_X1  g087(.A(G190gat), .B(G218gat), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n286), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n250), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT98), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT98), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n294), .B(new_n250), .C1(new_n290), .C2(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n286), .A2(new_n288), .ZN(new_n297));
  INV_X1    g096(.A(new_n289), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(new_n249), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT97), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT97), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n299), .A2(new_n300), .A3(new_n303), .A4(new_n249), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n245), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT103), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n211), .A2(new_n212), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n285), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n213), .A2(new_n284), .A3(new_n282), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT99), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n310), .A2(new_n316), .A3(new_n311), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n287), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n314), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT101), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT101), .ZN(new_n322));
  AOI211_X1 g121(.A(new_n322), .B(new_n314), .C1(new_n317), .C2(new_n318), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n315), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT102), .ZN(new_n325));
  XNOR2_X1  g124(.A(G120gat), .B(G148gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G176gat), .B(G204gat), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n326), .B(new_n327), .Z(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(new_n320), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n331), .A2(KEYINPUT100), .A3(new_n328), .A4(new_n315), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT100), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n328), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n325), .B1(new_n324), .B2(new_n329), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n308), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n329), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT102), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n342), .A2(KEYINPUT103), .A3(new_n337), .A4(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n307), .A2(new_n345), .A3(KEYINPUT104), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n296), .A2(new_n305), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n347), .A2(new_n244), .A3(new_n340), .A4(new_n343), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT104), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT94), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT69), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT69), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G113gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n356), .A3(G120gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT70), .ZN(new_n358));
  INV_X1    g157(.A(G120gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G113gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G134gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G127gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n220), .A2(G134gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT1), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n358), .B1(new_n357), .B2(new_n360), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n353), .A2(G120gat), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT1), .B1(new_n360), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT68), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT68), .ZN(new_n374));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n365), .B(new_n374), .C1(new_n375), .C2(KEYINPUT1), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT71), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n360), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT70), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n361), .A3(new_n366), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT71), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n373), .A2(new_n376), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n386));
  NOR2_X1   g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT24), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT24), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n387), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G169gat), .ZN(new_n393));
  INV_X1    g192(.A(G176gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT23), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT23), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(G169gat), .B2(G176gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(G169gat), .A2(G176gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n386), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT64), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT64), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(new_n386), .C1(new_n392), .C2(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT67), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n389), .A2(new_n391), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n407));
  INV_X1    g206(.A(G183gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G190gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT66), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT66), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n409), .A2(new_n414), .A3(new_n410), .A4(new_n411), .ZN(new_n415));
  AOI211_X1 g214(.A(new_n405), .B(new_n406), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n399), .A2(new_n386), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n406), .ZN(new_n420));
  AND2_X1   g219(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n423), .B2(new_n410), .ZN(new_n424));
  INV_X1    g223(.A(new_n415), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n420), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n419), .B1(new_n426), .B2(new_n405), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n404), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT27), .B(G183gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(KEYINPUT28), .A3(new_n410), .ZN(new_n430));
  NOR2_X1   g229(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n411), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(KEYINPUT27), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(G190gat), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n430), .B1(new_n434), .B2(KEYINPUT28), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n393), .A2(new_n394), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT26), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n388), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT26), .B1(new_n393), .B2(new_n394), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n398), .B2(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n385), .B1(new_n428), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n406), .B1(new_n413), .B2(new_n415), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n418), .B1(new_n443), .B2(KEYINPUT67), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n401), .B(new_n403), .C1(new_n444), .C2(new_n416), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n435), .A2(new_n440), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n445), .A2(new_n378), .A3(new_n384), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT73), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT34), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT72), .B(G71gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(new_n277), .ZN(new_n456));
  XOR2_X1   g255(.A(G15gat), .B(G43gat), .Z(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n448), .B1(new_n442), .B2(new_n447), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(KEYINPUT33), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n447), .ZN(new_n464));
  INV_X1    g263(.A(new_n448), .ZN(new_n465));
  AOI221_X4 g264(.A(new_n461), .B1(KEYINPUT33), .B2(new_n458), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n454), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n454), .B(KEYINPUT75), .C1(new_n463), .C2(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n464), .A2(new_n465), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT32), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n474), .A3(new_n458), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n449), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT34), .B1(new_n449), .B2(KEYINPUT73), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n462), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT74), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT74), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n475), .A2(new_n478), .A3(new_n482), .A4(new_n479), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n469), .A2(new_n470), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT77), .ZN(new_n485));
  NAND2_X1  g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n428), .B2(new_n441), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT29), .B1(new_n445), .B2(new_n446), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n487), .ZN(new_n490));
  XNOR2_X1  g289(.A(G197gat), .B(G204gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT22), .ZN(new_n492));
  INV_X1    g291(.A(G211gat), .ZN(new_n493));
  INV_X1    g292(.A(G218gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G211gat), .B(G218gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n488), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n486), .B1(new_n445), .B2(new_n446), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n428), .B2(new_n441), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n504), .B2(new_n486), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n501), .B1(new_n505), .B2(new_n500), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n499), .B1(new_n506), .B2(new_n498), .ZN(new_n507));
  XNOR2_X1  g306(.A(G8gat), .B(G36gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G64gat), .B(G92gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  OAI21_X1  g309(.A(new_n485), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n498), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n502), .A2(KEYINPUT76), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n490), .B2(KEYINPUT76), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n515), .B2(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(new_n510), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT77), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n507), .A2(new_n519), .A3(new_n510), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n513), .B(new_n510), .C1(new_n515), .C2(new_n512), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT30), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n511), .A2(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT78), .ZN(new_n524));
  INV_X1    g323(.A(G148gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n525), .B2(G141gat), .ZN(new_n526));
  INV_X1    g325(.A(G141gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(G141gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT79), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT79), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G162gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n237), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(G155gat), .A2(G162gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT2), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n527), .A2(G148gat), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT2), .B1(new_n543), .B2(new_n529), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n544), .A2(new_n536), .A3(new_n538), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n381), .A2(new_n383), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n534), .B2(new_n541), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(new_n381), .A3(new_n383), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(KEYINPUT5), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G225gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT82), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n532), .A2(new_n533), .B1(new_n537), .B2(new_n540), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(new_n545), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n542), .A2(KEYINPUT82), .A3(new_n546), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n378), .A2(new_n384), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT4), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n550), .A2(new_n565), .A3(new_n381), .A4(new_n383), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT83), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n369), .A2(new_n377), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT83), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n565), .A4(new_n550), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n564), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n554), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT5), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT3), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n548), .B1(new_n574), .B2(new_n550), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n550), .A2(new_n574), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n556), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n551), .A2(KEYINPUT4), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n561), .B2(new_n563), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n577), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT5), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G1gat), .B(G29gat), .Z(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G57gat), .B(G85gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n579), .A2(new_n585), .A3(KEYINPUT6), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT89), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT82), .B1(new_n542), .B2(new_n546), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n558), .A2(new_n557), .A3(new_n545), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n562), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n567), .A2(new_n570), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n578), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n555), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT5), .B1(new_n581), .B2(new_n582), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT87), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n605), .A3(new_n585), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n590), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n579), .A2(new_n585), .ZN(new_n608));
  INV_X1    g407(.A(new_n590), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT6), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT35), .B1(new_n592), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n574), .B1(new_n498), .B2(KEYINPUT29), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n596), .B2(new_n597), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n512), .B1(new_n577), .B2(new_n503), .ZN(new_n616));
  INV_X1    g415(.A(G228gat), .ZN(new_n617));
  INV_X1    g416(.A(G233gat), .ZN(new_n618));
  OAI22_X1  g417(.A1(new_n615), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n616), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n617), .B(new_n618), .C1(new_n613), .C2(new_n547), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT85), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G78gat), .B(G106gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT31), .B(G50gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(G22gat), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n620), .A2(new_n621), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n617), .A2(new_n618), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n620), .B2(new_n614), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT85), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n629), .B2(new_n631), .ZN(new_n634));
  INV_X1    g433(.A(G22gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n626), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n628), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n633), .B1(new_n628), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n484), .A2(new_n523), .A3(new_n612), .A4(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n467), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n481), .B2(new_n483), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n609), .B1(new_n602), .B2(new_n603), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT6), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n579), .A2(new_n590), .A3(new_n585), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n591), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n642), .A2(new_n647), .A3(new_n523), .A4(new_n639), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n640), .A2(KEYINPUT90), .B1(new_n648), .B2(KEYINPUT35), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n469), .A2(new_n470), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n481), .A2(new_n483), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n650), .A2(new_n651), .A3(new_n639), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT90), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n652), .A2(new_n653), .A3(new_n523), .A4(new_n612), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n602), .A2(new_n603), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n655), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n590), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT89), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n591), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n610), .B2(new_n607), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n517), .B1(new_n516), .B2(KEYINPUT37), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(KEYINPUT38), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n506), .A2(KEYINPUT88), .A3(new_n498), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n506), .A2(new_n498), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT88), .B1(new_n505), .B2(new_n512), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n663), .B(KEYINPUT37), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n516), .A2(KEYINPUT37), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT38), .B1(new_n668), .B2(new_n661), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n660), .A2(new_n667), .A3(new_n521), .A4(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n549), .A2(new_n551), .A3(new_n572), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT39), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT39), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n676), .A2(KEYINPUT86), .A3(new_n609), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT86), .B1(new_n676), .B2(new_n609), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n681), .B(new_n674), .C1(new_n677), .C2(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n511), .A2(new_n518), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n520), .A2(new_n522), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n686), .A3(new_n607), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n687), .A3(new_n639), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n463), .A2(new_n466), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n482), .B1(new_n689), .B2(new_n478), .ZN(new_n690));
  AND4_X1   g489(.A1(new_n482), .A2(new_n475), .A3(new_n478), .A4(new_n479), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n467), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT36), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n684), .A2(new_n647), .A3(new_n685), .ZN(new_n694));
  INV_X1    g493(.A(new_n639), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT36), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n650), .A2(new_n651), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n693), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n649), .A2(new_n654), .B1(new_n688), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n230), .A2(new_n269), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n230), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(new_n270), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(G229gat), .A2(G233gat), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(KEYINPUT93), .A3(KEYINPUT18), .A4(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n269), .A2(KEYINPUT17), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT17), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n266), .B2(new_n268), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n703), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n710), .A2(KEYINPUT18), .A3(new_n705), .A4(new_n701), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT93), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(G113gat), .B(G141gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(G169gat), .B(G197gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT92), .B(KEYINPUT12), .Z(new_n720));
  XOR2_X1   g519(.A(new_n719), .B(new_n720), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n705), .B(KEYINPUT13), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n230), .A2(new_n269), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n701), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n710), .A2(new_n705), .A3(new_n701), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT18), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n714), .A2(new_n721), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n721), .B1(new_n714), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n352), .B1(new_n700), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n612), .A2(new_n523), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n650), .A2(new_n651), .A3(new_n639), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT90), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n648), .A2(KEYINPUT35), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n654), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n699), .A2(new_n688), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n730), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(KEYINPUT94), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n351), .B1(new_n731), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n647), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT105), .B(G1gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1324gat));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n746));
  INV_X1    g545(.A(new_n351), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT94), .B1(new_n738), .B2(new_n739), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n352), .B(new_n730), .C1(new_n736), .C2(new_n737), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n686), .B(new_n747), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT16), .B(G8gat), .Z(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n746), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT106), .B(new_n746), .C1(new_n750), .C2(new_n752), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n741), .A2(KEYINPUT42), .A3(new_n686), .A4(new_n751), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n750), .A2(G8gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(G1325gat));
  INV_X1    g558(.A(new_n741), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n693), .A2(new_n698), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G15gat), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n484), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n764), .A2(G15gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n760), .B2(new_n765), .ZN(G1326gat));
  NAND2_X1  g565(.A1(new_n741), .A2(new_n695), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT43), .B(G22gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1327gat));
  NAND2_X1  g568(.A1(new_n731), .A2(new_n740), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n345), .A2(new_n245), .A3(new_n306), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT107), .Z(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n647), .A2(G29gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT44), .B1(new_n738), .B2(new_n306), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n780), .B(new_n347), .C1(new_n736), .C2(new_n737), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n244), .B(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n728), .B2(new_n729), .ZN(new_n786));
  INV_X1    g585(.A(new_n713), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n711), .A2(new_n712), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n727), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n721), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n714), .A2(new_n721), .A3(new_n727), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(KEYINPUT108), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n784), .A2(new_n344), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n782), .A2(new_n742), .A3(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n777), .B(new_n778), .C1(new_n252), .C2(new_n796), .ZN(G1328gat));
  NOR2_X1   g596(.A1(new_n523), .A2(G36gat), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n770), .A2(new_n773), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n780), .B1(new_n700), .B2(new_n347), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n738), .A2(KEYINPUT44), .A3(new_n306), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n801), .A2(new_n686), .A3(new_n802), .A4(new_n795), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n799), .A2(new_n800), .B1(G36gat), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n770), .A2(new_n773), .A3(new_n798), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT110), .B1(new_n805), .B2(KEYINPUT46), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(G1329gat));
  NOR2_X1   g607(.A1(new_n764), .A2(G43gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n770), .A2(new_n773), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT47), .B1(new_n810), .B2(KEYINPUT111), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n801), .A2(new_n761), .A3(new_n802), .A4(new_n795), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G43gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n813), .B(new_n810), .C1(KEYINPUT111), .C2(KEYINPUT47), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1330gat));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n695), .A3(new_n802), .A4(new_n795), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G50gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT48), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n639), .A2(G50gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n770), .A2(new_n773), .A3(new_n821), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n819), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(G1331gat));
  NAND3_X1  g624(.A1(new_n307), .A2(new_n344), .A3(new_n794), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n700), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n742), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g628(.A(new_n523), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n833));
  OR2_X1    g632(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n834));
  OR3_X1    g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n832), .B2(new_n833), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1333gat));
  NAND2_X1  g636(.A1(new_n827), .A2(new_n761), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n764), .A2(G71gat), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n838), .A2(G71gat), .B1(new_n827), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g640(.A1(new_n827), .A2(new_n695), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G78gat), .ZN(G1335gat));
  INV_X1    g642(.A(new_n794), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n244), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n345), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n782), .A2(new_n742), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n273), .A2(new_n275), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n851));
  NOR4_X1   g650(.A1(new_n700), .A2(new_n851), .A3(new_n347), .A4(new_n846), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n347), .B1(new_n736), .B2(new_n737), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT51), .B1(new_n853), .B2(new_n845), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n344), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n647), .A2(new_n849), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n850), .B1(new_n855), .B2(new_n856), .ZN(G1336gat));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n801), .A2(new_n686), .A3(new_n802), .A4(new_n847), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G92gat), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n523), .A2(G92gat), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n344), .B(new_n863), .C1(new_n852), .C2(new_n854), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n858), .A2(new_n859), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n860), .A2(new_n862), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n861), .B2(G92gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n860), .B1(new_n868), .B2(new_n864), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(G1337gat));
  NAND3_X1  g669(.A1(new_n738), .A2(new_n306), .A3(new_n845), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n851), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n853), .A2(KEYINPUT51), .A3(new_n845), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n345), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n277), .A3(new_n484), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n782), .A2(new_n761), .A3(new_n847), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n277), .ZN(G1338gat));
  NAND4_X1  g676(.A1(new_n801), .A2(new_n695), .A3(new_n802), .A4(new_n847), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n278), .B1(new_n878), .B2(KEYINPUT114), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n782), .A2(new_n880), .A3(new_n695), .A4(new_n847), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n639), .A2(G106gat), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n878), .A2(G106gat), .ZN(new_n886));
  INV_X1    g685(.A(new_n883), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n855), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(G1339gat));
  NAND2_X1  g689(.A1(new_n331), .A2(new_n322), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n335), .A2(KEYINPUT101), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n335), .A2(new_n892), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n317), .A2(new_n314), .A3(new_n318), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n328), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n897), .A3(KEYINPUT55), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n337), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT55), .B1(new_n894), .B2(new_n897), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n786), .A2(new_n901), .A3(new_n793), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT116), .B1(new_n704), .B2(new_n705), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n723), .A2(new_n701), .A3(new_n722), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n704), .A2(KEYINPUT116), .A3(new_n705), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n719), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n792), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n340), .B2(new_n343), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n347), .B1(new_n902), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n908), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n306), .A2(new_n911), .A3(new_n901), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n784), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n348), .B2(new_n844), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n345), .A2(new_n307), .A3(KEYINPUT115), .A4(new_n794), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n733), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n686), .A2(new_n647), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G113gat), .B1(new_n921), .B2(new_n730), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n742), .B1(new_n913), .B2(new_n917), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n642), .A2(new_n639), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT117), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n523), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n844), .A2(new_n354), .A3(new_n356), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n922), .B1(new_n929), .B2(new_n930), .ZN(G1340gat));
  NOR3_X1   g730(.A1(new_n921), .A2(new_n359), .A3(new_n345), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n523), .A3(new_n344), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n359), .ZN(G1341gat));
  INV_X1    g733(.A(new_n784), .ZN(new_n935));
  OAI21_X1  g734(.A(G127gat), .B1(new_n921), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n244), .A2(new_n220), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n929), .B2(new_n937), .ZN(G1342gat));
  NOR3_X1   g737(.A1(new_n686), .A2(G134gat), .A3(new_n347), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT56), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n928), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  OAI21_X1  g742(.A(G134gat), .B1(new_n921), .B2(new_n347), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(G1343gat));
  INV_X1    g744(.A(KEYINPUT118), .ZN(new_n946));
  INV_X1    g745(.A(new_n920), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n761), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n762), .A2(KEYINPUT118), .A3(new_n920), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n695), .B1(new_n913), .B2(new_n917), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n948), .B(new_n949), .C1(new_n950), .C2(KEYINPUT57), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n344), .A2(new_n911), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n739), .A2(new_n901), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n894), .A2(new_n897), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT55), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n337), .A3(new_n898), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n730), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT119), .B1(new_n909), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n955), .A2(new_n961), .A3(new_n347), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n244), .B1(new_n962), .B2(new_n912), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n695), .B1(new_n963), .B2(new_n917), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n951), .B1(KEYINPUT57), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n527), .B1(new_n965), .B2(new_n844), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n761), .A2(KEYINPUT120), .A3(new_n639), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT120), .B1(new_n761), .B2(new_n639), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n730), .A2(G141gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n523), .A2(new_n970), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n969), .A2(new_n923), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT58), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n527), .B1(new_n965), .B2(new_n739), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n924), .A2(KEYINPUT121), .A3(new_n968), .A4(new_n967), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n976), .B1(new_n969), .B2(new_n923), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n975), .A2(new_n977), .A3(new_n523), .A4(new_n970), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT58), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n973), .B1(new_n974), .B2(new_n980), .ZN(G1344gat));
  NOR2_X1   g780(.A1(new_n345), .A2(G148gat), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n975), .A2(new_n977), .A3(new_n523), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT122), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n639), .A2(KEYINPUT57), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n351), .A2(new_n739), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n963), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n950), .A2(KEYINPUT57), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n949), .A2(new_n344), .A3(new_n948), .ZN(new_n990));
  OAI21_X1  g789(.A(G148gat), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT59), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n525), .A2(KEYINPUT59), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n993), .B1(new_n965), .B2(new_n344), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g795(.A(KEYINPUT123), .B(new_n993), .C1(new_n965), .C2(new_n344), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n984), .B1(new_n996), .B2(new_n997), .ZN(G1345gat));
  NAND2_X1  g797(.A1(new_n975), .A2(new_n977), .ZN(new_n999));
  NOR4_X1   g798(.A1(new_n999), .A2(G155gat), .A3(new_n686), .A4(new_n245), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n237), .B1(new_n965), .B2(new_n784), .ZN(new_n1001));
  OR2_X1    g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1346gat));
  AND2_X1   g801(.A1(new_n965), .A2(new_n306), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n523), .A2(new_n535), .A3(new_n306), .ZN(new_n1004));
  OAI22_X1  g803(.A1(new_n1003), .A2(new_n535), .B1(new_n999), .B2(new_n1004), .ZN(G1347gat));
  NAND3_X1  g804(.A1(new_n919), .A2(new_n647), .A3(new_n686), .ZN(new_n1006));
  NOR3_X1   g805(.A1(new_n1006), .A2(new_n393), .A3(new_n730), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n647), .B1(new_n913), .B2(new_n917), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n1009));
  OR2_X1    g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n523), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1012), .A2(new_n926), .A3(new_n844), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1007), .B1(new_n1013), .B2(new_n393), .ZN(G1348gat));
  OAI21_X1  g813(.A(G176gat), .B1(new_n1006), .B2(new_n345), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1012), .A2(new_n926), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n344), .A2(new_n394), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(G1349gat));
  OAI21_X1  g817(.A(new_n432), .B1(new_n1006), .B2(new_n935), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n244), .A2(new_n429), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1019), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1021), .A2(KEYINPUT60), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT60), .ZN(new_n1023));
  OAI211_X1 g822(.A(new_n1023), .B(new_n1019), .C1(new_n1016), .C2(new_n1020), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1022), .A2(new_n1024), .ZN(G1350gat));
  OAI21_X1  g824(.A(G190gat), .B1(new_n1006), .B2(new_n347), .ZN(new_n1026));
  XNOR2_X1  g825(.A(new_n1026), .B(KEYINPUT61), .ZN(new_n1027));
  NAND4_X1  g826(.A1(new_n1012), .A2(new_n410), .A3(new_n926), .A4(new_n306), .ZN(new_n1028));
  INV_X1    g827(.A(KEYINPUT125), .ZN(new_n1029));
  AND2_X1   g828(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(G1351gat));
  INV_X1    g831(.A(new_n989), .ZN(new_n1033));
  NOR3_X1   g832(.A1(new_n761), .A2(new_n742), .A3(new_n523), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g834(.A1(new_n1035), .A2(new_n730), .ZN(new_n1036));
  XNOR2_X1  g835(.A(KEYINPUT126), .B(G197gat), .ZN(new_n1037));
  NOR2_X1   g836(.A1(new_n761), .A2(new_n639), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1012), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n844), .A2(new_n1037), .ZN(new_n1040));
  OAI22_X1  g839(.A1(new_n1036), .A2(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(G1352gat));
  NOR2_X1   g840(.A1(new_n345), .A2(G204gat), .ZN(new_n1042));
  NAND3_X1  g841(.A1(new_n1012), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  OR2_X1    g842(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1044));
  OAI21_X1  g843(.A(G204gat), .B1(new_n1035), .B2(new_n345), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(G1353gat));
  INV_X1    g846(.A(KEYINPUT63), .ZN(new_n1048));
  NAND4_X1  g847(.A1(new_n987), .A2(new_n988), .A3(new_n244), .A4(new_n1034), .ZN(new_n1049));
  NAND2_X1  g848(.A1(new_n1049), .A2(KEYINPUT127), .ZN(new_n1050));
  INV_X1    g849(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g850(.A(G211gat), .B1(new_n1049), .B2(KEYINPUT127), .ZN(new_n1052));
  OAI21_X1  g851(.A(new_n1048), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g852(.A(KEYINPUT127), .ZN(new_n1054));
  NAND4_X1  g853(.A1(new_n1033), .A2(new_n1054), .A3(new_n244), .A4(new_n1034), .ZN(new_n1055));
  NAND4_X1  g854(.A1(new_n1055), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n1050), .ZN(new_n1056));
  NAND2_X1  g855(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g856(.A1(new_n1012), .A2(new_n493), .A3(new_n244), .A4(new_n1038), .ZN(new_n1058));
  NAND2_X1  g857(.A1(new_n1057), .A2(new_n1058), .ZN(G1354gat));
  OAI21_X1  g858(.A(G218gat), .B1(new_n1035), .B2(new_n347), .ZN(new_n1060));
  NAND2_X1  g859(.A1(new_n306), .A2(new_n494), .ZN(new_n1061));
  OAI21_X1  g860(.A(new_n1060), .B1(new_n1039), .B2(new_n1061), .ZN(G1355gat));
endmodule


