//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1121, new_n1122;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G234));
  NAND2_X1  g027(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n456), .A2(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT69), .Z(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OR3_X1    g044(.A1(new_n469), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT70), .B1(new_n469), .B2(G2105), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n466), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n467), .A2(new_n472), .A3(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n466), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(KEYINPUT71), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  NOR3_X1   g058(.A1(new_n480), .A2(new_n483), .A3(new_n466), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n477), .A2(new_n479), .A3(new_n466), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n486), .A2(G124), .B1(G136), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n487), .A2(new_n495), .A3(G138), .A4(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n477), .A2(new_n479), .A3(G138), .A4(new_n466), .ZN(new_n498));
  XOR2_X1   g073(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n499));
  OAI21_X1  g074(.A(KEYINPUT75), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n464), .A2(KEYINPUT72), .A3(G138), .A4(new_n466), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n503), .A2(new_n504), .A3(new_n507), .A4(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n501), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n466), .A2(G114), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n481), .A2(G126), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G50), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n524), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n525), .A2(new_n527), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n520), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n516), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G51), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n538), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n523), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  INV_X1    g123(.A(G52), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n529), .A2(new_n548), .B1(new_n531), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n547), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(new_n537), .A2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n539), .A2(G43), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n523), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT76), .Z(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(KEYINPUT77), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n531), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(KEYINPUT77), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n520), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(G651), .A2(new_n572), .B1(new_n537), .B2(G91), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n567), .A2(new_n568), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n523), .B1(new_n520), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT78), .ZN(new_n578));
  AOI22_X1  g153(.A1(G87), .A2(new_n537), .B1(new_n539), .B2(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G288));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT79), .B1(new_n529), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n537), .A2(new_n583), .A3(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n520), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n539), .B2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(G85), .A2(new_n537), .B1(new_n539), .B2(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n523), .B2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n529), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G79), .ZN(new_n596));
  OR3_X1    g171(.A1(new_n596), .A2(new_n516), .A3(KEYINPUT80), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT80), .B1(new_n596), .B2(new_n516), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n520), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(new_n539), .B2(G54), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT10), .B1(new_n529), .B2(new_n594), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n595), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G860), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n603), .B1(G559), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT81), .Z(G148));
  OR2_X1    g189(.A1(new_n603), .A2(G559), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n557), .B2(G868), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n485), .A2(KEYINPUT83), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n466), .A2(G111), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n487), .A2(G135), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT83), .B1(new_n485), .B2(new_n619), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n470), .A2(new_n471), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(new_n480), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT13), .B(G2100), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n628), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT15), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2435), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n642), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(new_n643), .B2(new_n645), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  OAI21_X1  g224(.A(KEYINPUT84), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n648), .B2(new_n649), .ZN(new_n652));
  OR4_X1    g227(.A1(KEYINPUT84), .A2(new_n646), .A3(new_n647), .A4(new_n649), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n656), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n627), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT85), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n667), .B(new_n668), .Z(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  OAI22_X1  g252(.A1(new_n675), .A2(KEYINPUT20), .B1(new_n671), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(KEYINPUT20), .B2(new_n675), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n671), .A3(new_n674), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  INV_X1    g257(.A(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1991), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n681), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(G1986), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  NOR2_X1   g267(.A1(G95), .A2(G2105), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  OAI21_X1  g269(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n695));
  INV_X1    g270(.A(G131), .ZN(new_n696));
  OAI22_X1  g271(.A1(new_n694), .A2(new_n695), .B1(new_n473), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n486), .B2(G119), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(new_n691), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT35), .B(G1991), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT88), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT89), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G16), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G6), .B(G305), .S(G16), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n713), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n713), .A2(new_n718), .A3(new_n721), .A4(KEYINPUT90), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n708), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n708), .A3(new_n725), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n707), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n691), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n691), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n729), .A2(KEYINPUT36), .B1(G2078), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n714), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n714), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1961), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G16), .A2(G19), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n557), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1341), .ZN(new_n739));
  NOR2_X1   g314(.A1(G29), .A2(G32), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n487), .A2(G141), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT26), .Z(new_n743));
  INV_X1    g318(.A(G105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n743), .C1(new_n629), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n486), .B2(G129), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT27), .B(G1996), .Z(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n739), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n731), .A2(G2078), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n732), .A2(new_n736), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(KEYINPUT30), .A2(G28), .ZN(new_n753));
  NOR2_X1   g328(.A1(KEYINPUT30), .A2(G28), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n691), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n755), .B(new_n756), .C1(new_n626), .C2(new_n691), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT96), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n691), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  NOR2_X1   g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n764));
  INV_X1    g339(.A(G140), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n763), .A2(new_n764), .B1(new_n473), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n486), .B2(G128), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(new_n691), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(G29), .A2(G33), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n487), .A2(G139), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n775), .C1(new_n466), .C2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n771), .B1(new_n777), .B2(new_n691), .ZN(new_n778));
  INV_X1    g353(.A(G2072), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n770), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G21), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G168), .B2(G16), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n747), .A2(new_n748), .B1(new_n785), .B2(G1966), .ZN(new_n786));
  INV_X1    g361(.A(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(G1966), .ZN(new_n788));
  OR2_X1    g363(.A1(KEYINPUT24), .A2(G34), .ZN(new_n789));
  NAND2_X1  g364(.A1(KEYINPUT24), .A2(G34), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n789), .A2(new_n691), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G160), .B2(new_n691), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n787), .A2(new_n788), .B1(G2084), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n758), .A2(new_n783), .A3(new_n786), .A4(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n707), .ZN(new_n795));
  INV_X1    g370(.A(new_n728), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n726), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n691), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n691), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G2090), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT98), .Z(new_n804));
  NOR2_X1   g379(.A1(new_n792), .A2(G2084), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT97), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n714), .A2(KEYINPUT23), .A3(G20), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT23), .ZN(new_n808));
  INV_X1    g383(.A(G20), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G16), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n810), .C1(new_n609), .C2(new_n714), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n799), .A2(new_n804), .A3(new_n806), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n603), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G16), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G4), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT92), .B(G1348), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n802), .A2(G2090), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n752), .A2(new_n814), .A3(new_n819), .A4(new_n820), .ZN(G311));
  NOR2_X1   g396(.A1(new_n752), .A2(new_n814), .ZN(new_n822));
  INV_X1    g397(.A(new_n819), .ZN(new_n823));
  INV_X1    g398(.A(new_n820), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n520), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G651), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT99), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n539), .A2(G55), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT100), .B(G93), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n830), .B(new_n831), .C1(new_n529), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n557), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n529), .A2(new_n832), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n830), .A2(new_n556), .A3(new_n835), .A4(new_n831), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n815), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n612), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT101), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n833), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n698), .B(KEYINPUT102), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n487), .A2(G142), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n466), .A2(G118), .ZN(new_n851));
  INV_X1    g426(.A(G130), .ZN(new_n852));
  OAI221_X1 g427(.A(new_n849), .B1(new_n850), .B2(new_n851), .C1(new_n485), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n632), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n848), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n514), .B(new_n767), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n777), .B(new_n746), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n855), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G160), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n626), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n493), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(KEYINPUT103), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n858), .Z(new_n865));
  OAI211_X1 g440(.A(new_n847), .B(new_n863), .C1(new_n865), .C2(new_n862), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(G395));
  NAND2_X1  g443(.A1(new_n833), .A2(new_n604), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(G303), .B(G290), .Z(new_n871));
  XNOR2_X1  g446(.A(G305), .B(G288), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT42), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n837), .B(new_n615), .Z(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n603), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(G299), .A2(new_n603), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n877), .A2(KEYINPUT41), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT41), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(KEYINPUT106), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n880), .A2(KEYINPUT106), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n877), .A2(new_n878), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n875), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n875), .B2(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n874), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  INV_X1    g466(.A(new_n874), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n884), .A4(new_n887), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n870), .B1(new_n894), .B2(G868), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT107), .ZN(G295));
  NAND2_X1  g471(.A1(new_n894), .A2(G868), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n869), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n899));
  XNOR2_X1  g474(.A(G301), .B(G286), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n834), .A2(new_n836), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n834), .B2(new_n836), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n837), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n886), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n834), .A2(new_n836), .A3(new_n900), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n881), .A2(new_n909), .A3(new_n882), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n873), .ZN(new_n912));
  OAI211_X1 g487(.A(KEYINPUT109), .B(new_n847), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n910), .A3(new_n912), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n907), .B2(new_n910), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n903), .A2(new_n906), .B1(new_n880), .B2(new_n879), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n909), .A2(new_n877), .A3(new_n878), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n873), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n921), .A2(new_n847), .A3(new_n914), .ZN(new_n922));
  MUX2_X1   g497(.A(new_n918), .B(new_n922), .S(KEYINPUT43), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT44), .ZN(new_n924));
  MUX2_X1   g499(.A(new_n922), .B(new_n918), .S(KEYINPUT43), .Z(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n514), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  XOR2_X1   g506(.A(KEYINPUT110), .B(G40), .Z(new_n932));
  NOR2_X1   g507(.A1(new_n860), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(G1996), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(KEYINPUT46), .ZN(new_n936));
  INV_X1    g511(.A(new_n934), .ZN(new_n937));
  INV_X1    g512(.A(new_n746), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n767), .B(new_n769), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(KEYINPUT46), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT127), .Z(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT47), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n934), .A2(G1996), .A3(new_n938), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT111), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n697), .B(new_n700), .C1(new_n486), .C2(G119), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n938), .A2(G1996), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n937), .B1(new_n939), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(KEYINPUT111), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n767), .A2(new_n769), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n934), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n698), .B(new_n700), .Z(new_n954));
  NAND2_X1  g529(.A1(new_n937), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n946), .A2(new_n949), .A3(new_n950), .A4(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n934), .A2(G1986), .A3(G290), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT48), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n944), .A2(new_n953), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n509), .B2(new_n513), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n933), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n964));
  OR3_X1    g539(.A1(new_n963), .A2(new_n964), .A3(G2078), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n966));
  INV_X1    g541(.A(G1961), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n930), .A2(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n933), .A3(new_n970), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n965), .A2(new_n966), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n966), .B2(new_n965), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(G171), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT113), .B(G8), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(G168), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(KEYINPUT51), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n788), .B1(new_n963), .B2(new_n964), .ZN(new_n979));
  INV_X1    g554(.A(G2084), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n968), .A2(new_n980), .A3(new_n933), .A4(new_n970), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n982), .B2(new_n976), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n979), .B2(new_n981), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT51), .B1(new_n985), .B2(new_n977), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n977), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n974), .B1(new_n990), .B2(KEYINPUT62), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n717), .B1(new_n963), .B2(new_n964), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G2090), .B2(new_n971), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n975), .ZN(new_n994));
  NAND2_X1  g569(.A1(G303), .A2(G8), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT55), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n585), .A2(new_n683), .A3(new_n589), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n537), .A2(G86), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n589), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G1981), .ZN(new_n1001));
  OR2_X1    g576(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n961), .A2(new_n933), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n998), .A2(new_n1001), .A3(KEYINPUT114), .A4(KEYINPUT49), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n975), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G288), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1006), .A2(new_n975), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n976), .B(new_n1010), .C1(new_n961), .C2(new_n933), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1008), .B(new_n1013), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1006), .A2(new_n975), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n1019), .B2(new_n1010), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1020), .A2(KEYINPUT116), .A3(new_n1008), .A4(new_n1013), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n996), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n993), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n997), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n983), .A2(new_n986), .B1(new_n977), .B2(new_n988), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n991), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1024), .A2(new_n1016), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1008), .A2(new_n1009), .A3(new_n710), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n998), .B(KEYINPUT115), .Z(new_n1032));
  AOI21_X1  g607(.A(new_n1019), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g608(.A(G286), .B(new_n976), .C1(new_n979), .C2(new_n981), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n997), .A2(new_n1022), .A3(new_n1024), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n993), .A2(G8), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1016), .B1(new_n1038), .B2(new_n996), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(KEYINPUT63), .A3(new_n1024), .A4(new_n1034), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1033), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1029), .A2(new_n1030), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n969), .B1(new_n514), .B2(new_n929), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT50), .B(G1384), .C1(new_n509), .C2(new_n513), .ZN(new_n1044));
  INV_X1    g619(.A(new_n933), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT117), .B1(new_n1046), .B2(G1956), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n930), .A2(new_n931), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(new_n779), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(new_n933), .A3(new_n962), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n971), .A2(new_n1052), .A3(new_n812), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1047), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(G299), .B(KEYINPUT57), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1348), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1006), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n971), .A2(new_n1057), .B1(new_n769), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n603), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1055), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1047), .A2(new_n1061), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT119), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1048), .A2(new_n933), .A3(new_n962), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT58), .B(G1341), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1068), .A2(G1996), .B1(new_n1058), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n557), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1070), .B2(new_n557), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1058), .A2(new_n769), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT60), .B(new_n1075), .C1(new_n1046), .C2(G1348), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1076), .A2(KEYINPUT121), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1076), .A2(KEYINPUT121), .A3(new_n603), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n603), .B1(new_n1076), .B2(KEYINPUT121), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1059), .A2(KEYINPUT60), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1074), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1064), .A2(new_n1083), .A3(new_n1065), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1067), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1056), .A2(KEYINPUT61), .A3(new_n1062), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT120), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1063), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1026), .A2(new_n1025), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  OAI221_X1 g665(.A(new_n1090), .B1(new_n473), .B2(new_n474), .C1(new_n629), .C2(new_n468), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT122), .B1(new_n475), .B2(new_n472), .ZN(new_n1092));
  INV_X1    g667(.A(new_n467), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(G40), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1048), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n966), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1048), .A2(new_n1096), .A3(KEYINPUT124), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n963), .A2(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT125), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1099), .A2(new_n1104), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1103), .A2(G301), .A3(new_n972), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT54), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n974), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n973), .A2(G301), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1103), .A2(G171), .A3(new_n972), .A4(new_n1105), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(KEYINPUT54), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1089), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1042), .B1(new_n1088), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G290), .B(G1986), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n956), .B1(new_n937), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT112), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n960), .B1(new_n1115), .B2(new_n1118), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g694(.A(G227), .ZN(new_n1121));
  AND3_X1   g695(.A1(new_n866), .A2(new_n654), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g696(.A1(new_n925), .A2(G319), .A3(new_n689), .A4(new_n1122), .ZN(G225));
  INV_X1    g697(.A(G225), .ZN(G308));
endmodule


