//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n209), .A2(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  NAND4_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n209), .A2(KEYINPUT0), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n216), .A2(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(G1), .A2(G13), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G13), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  OR2_X1    g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n204), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G150), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G58), .A2(G68), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n204), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n246), .A2(new_n204), .A3(G1), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n263), .A2(new_n244), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n253), .A2(KEYINPUT9), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n243), .B1(G33), .B2(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n269), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(G226), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G222), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G223), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n280), .B(new_n267), .C1(G77), .C2(new_n276), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n275), .A2(G190), .A3(new_n281), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT10), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n266), .A2(new_n283), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT9), .B1(new_n253), .B2(new_n265), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n285), .A2(KEYINPUT10), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n253), .A2(new_n265), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n282), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n294), .C1(G179), .C2(new_n282), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G68), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n255), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(new_n244), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n301), .A2(KEYINPUT11), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n245), .A2(new_n248), .A3(G68), .A4(new_n251), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n264), .A2(new_n297), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT12), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(KEYINPUT11), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n302), .A2(new_n304), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n278), .A2(G232), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G226), .B2(G1698), .ZN(new_n311));
  INV_X1    g0111(.A(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n309), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n267), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n270), .B1(G238), .B2(new_n274), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT13), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G169), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(KEYINPUT70), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n325), .A2(new_n327), .B1(new_n328), .B2(new_n324), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n325), .A2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n308), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(new_n308), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n333), .C1(new_n334), .C2(new_n324), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n251), .A2(G77), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n249), .A2(new_n336), .B1(G77), .B2(new_n248), .ZN(new_n337));
  INV_X1    g0137(.A(new_n254), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT15), .B(G87), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n255), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n341), .B2(new_n244), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n276), .A2(G232), .A3(new_n278), .ZN(new_n344));
  INV_X1    g0144(.A(G107), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n276), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n267), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n270), .B1(G244), .B2(new_n274), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n342), .B1(new_n349), .B2(new_n293), .ZN(new_n350));
  INV_X1    g0150(.A(new_n349), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n328), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n342), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(G200), .B2(new_n349), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(G190), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n331), .A2(new_n335), .A3(new_n358), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n296), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n254), .B1(new_n203), .B2(G20), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT75), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n362), .A2(new_n250), .B1(new_n248), .B2(new_n338), .ZN(new_n363));
  INV_X1    g0163(.A(G58), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n297), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(new_n260), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(G20), .B1(G159), .B2(new_n257), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n316), .A2(new_n368), .A3(new_n204), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT71), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n314), .A2(G33), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT71), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n204), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT16), .B(new_n367), .C1(new_n377), .C2(new_n297), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n378), .A2(new_n244), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT73), .B1(new_n314), .B2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n312), .A3(KEYINPUT3), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(new_n315), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n376), .A2(G20), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n387));
  NOR2_X1   g0187(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n276), .B2(G20), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n297), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n367), .B1(new_n391), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n380), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n363), .B1(new_n379), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n270), .B1(G232), .B2(new_n274), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n313), .A2(new_n315), .A3(G223), .A4(new_n278), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n313), .A2(new_n315), .A3(G226), .A4(G1698), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT76), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT76), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n276), .A2(new_n404), .A3(G226), .A4(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n401), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n267), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n405), .ZN(new_n409));
  INV_X1    g0209(.A(new_n401), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n334), .B(new_n398), .C1(new_n408), .C2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n398), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n272), .B1(new_n411), .B2(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n406), .A2(new_n407), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(G200), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT17), .B1(new_n397), .B2(new_n418), .ZN(new_n420));
  NOR2_X1   g0220(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n363), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n366), .A2(G20), .ZN(new_n424));
  INV_X1    g0224(.A(G159), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n258), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n386), .A2(new_n390), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G68), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n428), .B2(KEYINPUT74), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT16), .B1(new_n429), .B2(new_n393), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n378), .A2(new_n244), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n423), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(G179), .B(new_n398), .C1(new_n408), .C2(new_n412), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n417), .B2(new_n293), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n422), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n419), .A2(new_n420), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n432), .B2(new_n434), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT78), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n360), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT5), .B(G41), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n267), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G270), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n447), .A2(new_n446), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n267), .A2(new_n268), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n316), .A2(G303), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n313), .A2(new_n315), .A3(G257), .A4(new_n278), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n313), .A2(new_n315), .A3(G264), .A4(G1698), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n455), .A2(KEYINPUT82), .A3(new_n456), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT83), .B1(new_n462), .B2(new_n267), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  AOI211_X1 g0264(.A(new_n464), .B(new_n272), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n454), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n248), .A2(G116), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n204), .C1(G33), .C2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n244), .C1(new_n204), .C2(G116), .ZN(new_n472));
  OR3_X1    g0272(.A1(new_n472), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n312), .A2(G1), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n264), .A2(new_n244), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G116), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n468), .A2(new_n473), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n466), .A2(KEYINPUT21), .A3(G169), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n462), .A2(new_n267), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n464), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n462), .A2(KEYINPUT83), .A3(new_n267), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT86), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n453), .A2(new_n328), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n479), .A4(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n479), .B(new_n486), .C1(new_n463), .C2(new_n465), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT86), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT87), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n480), .A2(new_n487), .A3(new_n489), .A4(KEYINPUT87), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n466), .A2(G169), .A3(new_n479), .ZN(new_n494));
  XOR2_X1   g0294(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n479), .B1(new_n466), .B2(G200), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n334), .B2(new_n466), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n492), .A2(new_n493), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n276), .A2(new_n204), .A3(G87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n276), .A2(new_n502), .A3(new_n204), .A4(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n312), .A2(new_n505), .A3(G20), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n204), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n345), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT24), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n504), .A2(new_n513), .A3(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n244), .ZN(new_n516));
  INV_X1    g0316(.A(new_n477), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT25), .B1(new_n264), .B2(new_n345), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n345), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n517), .A2(new_n345), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n516), .A2(KEYINPUT89), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT89), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n245), .B1(new_n512), .B2(new_n514), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n313), .A2(new_n315), .A3(G257), .A4(G1698), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n313), .A2(new_n315), .A3(G250), .A4(new_n278), .ZN(new_n527));
  INV_X1    g0327(.A(G294), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n312), .C2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n267), .B1(new_n448), .B2(G264), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n452), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G169), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n328), .B2(new_n531), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n522), .A2(new_n525), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT90), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n522), .A2(new_n525), .A3(new_n533), .A4(KEYINPUT90), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n345), .A2(KEYINPUT6), .A3(G97), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT79), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n470), .A2(new_n345), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n541), .A2(new_n542), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G20), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n257), .A2(G77), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n345), .B1(new_n386), .B2(new_n390), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n244), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n313), .A2(new_n315), .A3(G244), .A4(new_n278), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(KEYINPUT80), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(KEYINPUT80), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n276), .A2(G244), .A3(new_n278), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n557), .A2(new_n469), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n267), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n448), .A2(G257), .B1(new_n450), .B2(new_n451), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(G190), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n248), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n477), .B2(G97), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n554), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G200), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n562), .B2(new_n563), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n540), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n566), .ZN(new_n571));
  INV_X1    g0371(.A(new_n553), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n551), .A3(new_n550), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(new_n244), .ZN(new_n574));
  INV_X1    g0374(.A(new_n569), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT81), .A4(new_n564), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n204), .B1(new_n309), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n546), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n313), .A2(new_n315), .A3(new_n204), .A4(G68), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n578), .B1(new_n255), .B2(new_n470), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n244), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n340), .A2(new_n264), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n477), .A2(G87), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n272), .A2(G274), .A3(new_n446), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n203), .A2(G45), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n272), .A2(G250), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n313), .A2(new_n315), .A3(G238), .A4(new_n278), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n313), .A2(new_n315), .A3(G244), .A4(G1698), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n594), .B(new_n595), .C1(new_n312), .C2(new_n505), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n593), .B1(new_n596), .B2(new_n267), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G190), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n589), .B(new_n598), .C1(new_n568), .C2(new_n597), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n328), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n586), .B(new_n587), .C1(new_n517), .C2(new_n340), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(G169), .C2(new_n597), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n524), .A2(new_n520), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n531), .A2(new_n334), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n568), .B1(new_n530), .B2(new_n452), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n574), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n562), .A2(new_n563), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n328), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n562), .A2(new_n563), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n293), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n577), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n539), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n444), .A2(new_n499), .A3(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n335), .A2(new_n354), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n420), .B(new_n419), .C1(new_n331), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n432), .A2(new_n434), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT18), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n438), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n291), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(new_n295), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n496), .A2(new_n489), .A3(new_n480), .A4(new_n487), .ZN(new_n625));
  INV_X1    g0425(.A(new_n604), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n533), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n615), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n602), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  OR3_X1    g0430(.A1(new_n614), .A2(new_n630), .A3(new_n603), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n614), .B2(new_n603), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n624), .B1(new_n444), .B2(new_n635), .ZN(G369));
  NAND2_X1  g0436(.A1(new_n247), .A2(new_n204), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n638), .A2(new_n639), .A3(G213), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G343), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT91), .Z(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n479), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n625), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n499), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n604), .A2(new_n607), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n643), .A2(new_n522), .A3(new_n525), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n536), .A2(new_n649), .A3(new_n537), .A4(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n534), .A2(new_n642), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n539), .A2(new_n655), .A3(new_n649), .A4(new_n642), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n627), .A2(new_n642), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n654), .A2(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n207), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G41), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n581), .A2(G116), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G1), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n212), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(new_n662), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n492), .A2(new_n493), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n536), .A2(new_n496), .A3(new_n537), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n615), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n643), .B1(new_n670), .B2(new_n633), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT29), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n643), .B1(new_n628), .B2(new_n633), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT29), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n486), .B1(new_n463), .B2(new_n465), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n530), .A2(new_n597), .A3(KEYINPUT92), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT92), .B1(new_n530), .B2(new_n597), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n610), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n597), .A2(G179), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n466), .A2(new_n612), .A3(new_n531), .A4(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n677), .A2(new_n680), .A3(new_n676), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT93), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n681), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n679), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n530), .A2(new_n597), .A3(KEYINPUT92), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n612), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n484), .A3(KEYINPUT30), .A4(new_n486), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(KEYINPUT93), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n643), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT31), .B(new_n643), .C1(new_n686), .C2(new_n691), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n615), .A2(new_n536), .A3(new_n537), .A4(new_n642), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n694), .B(new_n695), .C1(new_n499), .C2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n675), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n667), .B1(new_n700), .B2(G1), .ZN(G364));
  INV_X1    g0501(.A(new_n648), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n246), .A2(G20), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n203), .B1(new_n703), .B2(G45), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n661), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(G330), .B2(new_n647), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n207), .A2(new_n276), .ZN(new_n709));
  INV_X1    g0509(.A(G355), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n709), .A2(new_n710), .B1(G116), .B2(new_n207), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n373), .A2(new_n374), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n660), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n445), .B2(new_n212), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n237), .A2(new_n445), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n243), .B1(G20), .B2(new_n293), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n706), .B1(new_n718), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n722), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n204), .A2(G179), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n334), .A3(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n345), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n204), .A2(new_n328), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G190), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n334), .A2(G179), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n204), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n733), .A2(new_n364), .B1(new_n470), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n731), .A2(new_n568), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n729), .B(new_n736), .C1(G50), .C2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n739));
  NOR2_X1   g0539(.A1(G190), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n727), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT94), .B(G159), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n727), .A2(G190), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n580), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n730), .A2(new_n334), .A3(G200), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n276), .B1(new_n748), .B2(new_n297), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n730), .A2(new_n740), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n749), .B1(G77), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n738), .A2(new_n743), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n735), .ZN(new_n754));
  INV_X1    g0554(.A(new_n745), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n754), .A2(G294), .B1(new_n755), .B2(G303), .ZN(new_n756));
  INV_X1    g0556(.A(new_n748), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n276), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n741), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G311), .A2(new_n751), .B1(new_n760), .B2(G329), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n756), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G322), .A2(new_n732), .B1(new_n737), .B2(G326), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n728), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n726), .B1(new_n753), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n725), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n721), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n647), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n708), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(G396));
  INV_X1    g0571(.A(new_n737), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n733), .A2(new_n528), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G107), .B2(new_n755), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n750), .A2(new_n505), .B1(new_n741), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n276), .B(new_n777), .C1(G283), .C2(new_n757), .ZN(new_n778));
  INV_X1    g0578(.A(new_n728), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n754), .A2(G97), .B1(new_n779), .B2(G87), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n775), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n712), .B1(G132), .B2(new_n760), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n735), .A2(new_n364), .B1(new_n745), .B2(new_n261), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n728), .A2(new_n297), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n742), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n757), .A2(G150), .B1(new_n751), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G137), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT96), .B(G143), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(new_n772), .B2(new_n788), .C1(new_n733), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n782), .B(new_n785), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n781), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n722), .ZN(new_n795));
  INV_X1    g0595(.A(new_n706), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n722), .A2(new_n719), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(new_n299), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n643), .A2(new_n355), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n358), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n354), .A2(KEYINPUT97), .A3(new_n643), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT97), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n353), .B2(new_n642), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n795), .B(new_n798), .C1(new_n805), .C2(new_n720), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n673), .B(new_n805), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n807), .A2(new_n698), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT98), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n796), .C1(new_n698), .C2(new_n807), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(KEYINPUT98), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(G384));
  NAND2_X1  g0612(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n243), .A2(new_n204), .A3(new_n505), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n549), .B2(KEYINPUT35), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT36), .Z(new_n819));
  NOR3_X1   g0619(.A1(new_n665), .A2(new_n299), .A3(new_n365), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n261), .B2(G68), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n246), .A2(G1), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT100), .Z(new_n824));
  NAND2_X1  g0624(.A1(new_n643), .A2(new_n308), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n331), .A2(new_n335), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(new_n331), .B2(new_n335), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n697), .A2(new_n805), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n377), .A2(new_n297), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT16), .B1(new_n831), .B2(new_n367), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n423), .B1(new_n832), .B2(new_n431), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n640), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n436), .B2(new_n441), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n397), .A2(new_n418), .B1(new_n833), .B2(new_n640), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n434), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n397), .A2(new_n418), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n432), .A2(new_n640), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n840), .A2(new_n620), .A3(new_n841), .A4(new_n836), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n835), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n834), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT78), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n621), .B2(new_n438), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT17), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n840), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n620), .A2(new_n421), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n418), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n847), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n837), .A2(new_n838), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n842), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT102), .B1(new_n846), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n845), .B1(new_n835), .B2(new_n844), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n855), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT102), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n830), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(KEYINPUT40), .ZN(new_n866));
  INV_X1    g0666(.A(new_n805), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n828), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n697), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT40), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n840), .A2(new_n620), .A3(new_n841), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(KEYINPUT103), .A3(new_n842), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n851), .A2(new_n621), .A3(new_n438), .A4(new_n853), .ZN(new_n874));
  INV_X1    g0674(.A(new_n841), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT103), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n871), .A2(new_n877), .A3(KEYINPUT37), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n845), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n870), .B1(new_n880), .B2(new_n862), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n866), .B1(new_n869), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n443), .A2(new_n697), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(G330), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n882), .A2(new_n883), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n860), .A2(new_n864), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n643), .A2(new_n353), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT101), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n673), .B2(new_n805), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n828), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n842), .A2(KEYINPUT103), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n897), .A2(new_n872), .B1(new_n875), .B2(new_n874), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n898), .B2(new_n878), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n896), .B1(new_n899), .B2(new_n846), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n331), .A2(new_n643), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT39), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n640), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n622), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n895), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n443), .A2(new_n672), .A3(new_n674), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n624), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n888), .A2(new_n911), .B1(new_n203), .B2(new_n703), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n888), .A2(new_n911), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n824), .B1(new_n912), .B2(new_n913), .ZN(G367));
  INV_X1    g0714(.A(KEYINPUT107), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n614), .A2(new_n642), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n577), .A2(new_n614), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n643), .A2(new_n609), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n656), .A2(new_n657), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT45), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n656), .A2(KEYINPUT45), .A3(new_n657), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n656), .B2(new_n657), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n658), .A2(new_n919), .ZN(new_n929));
  INV_X1    g0729(.A(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n925), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n654), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n926), .B(new_n930), .ZN(new_n934));
  INV_X1    g0734(.A(new_n654), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n925), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n655), .A2(new_n642), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n653), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n656), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT106), .B1(new_n647), .B2(G330), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n702), .A2(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n702), .A2(new_n940), .A3(KEYINPUT106), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n700), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n915), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n699), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n949), .A2(KEYINPUT107), .A3(new_n933), .A4(new_n936), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n700), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n661), .B(KEYINPUT41), .Z(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n705), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n656), .A2(new_n919), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n538), .A2(new_n917), .A3(new_n918), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n643), .B1(new_n959), .B2(new_n614), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n957), .B1(new_n961), .B2(KEYINPUT104), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n958), .B2(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n642), .A2(new_n589), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(new_n603), .Z(new_n967));
  INV_X1    g0767(.A(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n965), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n962), .A2(new_n968), .A3(new_n967), .A4(new_n964), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n935), .A2(new_n919), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n974), .A3(new_n972), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n967), .A2(new_n721), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n723), .B1(new_n207), .B2(new_n340), .C1(new_n715), .C2(new_n233), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n772), .A2(new_n789), .B1(new_n364), .B2(new_n745), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G150), .B2(new_n732), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n750), .A2(new_n261), .B1(new_n741), .B2(new_n788), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n316), .B(new_n983), .C1(new_n786), .C2(new_n757), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n754), .A2(G68), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n779), .A2(G77), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n982), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n772), .A2(new_n776), .B1(new_n345), .B2(new_n735), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G97), .B2(new_n779), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n748), .A2(new_n528), .B1(new_n750), .B2(new_n764), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G317), .B2(new_n760), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n713), .B1(G303), .B2(new_n732), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n755), .A2(G116), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT46), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n989), .A2(new_n991), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  OAI211_X1 g0797(.A(new_n706), .B(new_n980), .C1(new_n997), .C2(new_n726), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n955), .A2(new_n978), .B1(new_n979), .B2(new_n998), .ZN(G387));
  NOR2_X1   g0799(.A1(new_n949), .A2(new_n662), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n699), .A2(new_n944), .A3(new_n945), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n653), .A2(new_n721), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n230), .A2(G45), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n445), .B1(new_n297), .B2(new_n299), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n663), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(new_n1005), .B2(KEYINPUT109), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT50), .B1(new_n338), .B2(new_n261), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n338), .A2(KEYINPUT50), .A3(new_n261), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1006), .B1(KEYINPUT109), .B2(new_n1005), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1003), .A2(new_n714), .A3(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(G107), .B2(new_n207), .C1(new_n663), .C2(new_n709), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(new_n723), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n772), .A2(new_n425), .B1(new_n745), .B2(new_n299), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n713), .B1(new_n470), .B2(new_n728), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G68), .A2(new_n751), .B1(new_n760), .B2(G150), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n254), .B2(new_n748), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n735), .A2(new_n340), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n733), .B2(new_n261), .ZN(new_n1018));
  OR4_X1    g0818(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n713), .B1(G326), .B2(new_n760), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n735), .A2(new_n764), .B1(new_n745), .B2(new_n528), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n757), .A2(G311), .B1(new_n751), .B2(G303), .ZN(new_n1022));
  INV_X1    g0822(.A(G322), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(new_n772), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G317), .B2(new_n732), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT110), .Z(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1021), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1020), .B1(new_n505), .B2(new_n728), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1019), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n796), .B(new_n1012), .C1(new_n1033), .C2(new_n722), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1000), .A2(new_n1001), .B1(new_n1002), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n946), .A2(new_n705), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT108), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(G393));
  AOI22_X1  g0838(.A1(G150), .A2(new_n737), .B1(new_n732), .B2(G159), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT51), .Z(new_n1040));
  NAND2_X1  g0840(.A1(new_n754), .A2(G77), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n757), .A2(G50), .B1(new_n751), .B2(new_n338), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n297), .A2(new_n745), .B1(new_n728), .B2(new_n580), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n741), .A2(new_n789), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n712), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT112), .Z(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n732), .B1(new_n737), .B2(G317), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT52), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n316), .B1(new_n741), .B2(new_n1023), .C1(new_n528), .C2(new_n750), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n729), .B(new_n1050), .C1(G283), .C2(new_n755), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n754), .A2(G116), .B1(new_n757), .B2(G303), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT113), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT113), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1043), .A2(new_n1047), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT114), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n726), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n723), .B1(new_n470), .B2(new_n207), .C1(new_n715), .C2(new_n240), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n706), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT111), .Z(new_n1062));
  AND2_X1   g0862(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n919), .A2(new_n721), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n937), .B2(new_n704), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n662), .B1(new_n937), .B2(new_n947), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n951), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT115), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(G390));
  INV_X1    g0870(.A(new_n797), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1041), .B1(new_n772), .B2(new_n764), .C1(new_n505), .C2(new_n733), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G97), .A2(new_n751), .B1(new_n760), .B2(G294), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1073), .B(new_n316), .C1(new_n345), .C2(new_n748), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1072), .A2(new_n1074), .A3(new_n746), .A4(new_n784), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G159), .A2(new_n754), .B1(new_n737), .B2(G128), .ZN(new_n1076));
  INV_X1    g0876(.A(G132), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n733), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT54), .B(G143), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n757), .A2(G137), .B1(new_n751), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(G125), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1081), .B1(new_n1082), .B2(new_n741), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n745), .A2(new_n256), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT53), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1078), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n276), .B1(new_n728), .B2(new_n261), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT120), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1075), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n706), .B1(new_n338), .B2(new_n1071), .C1(new_n1091), .C2(new_n726), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n900), .A2(new_n903), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n719), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n901), .B1(new_n893), .B2(new_n828), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n643), .B(new_n867), .C1(new_n670), .C2(new_n633), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n829), .B1(new_n1096), .B2(new_n892), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n901), .B(KEYINPUT116), .Z(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n880), .B2(new_n862), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1093), .A2(new_n1095), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n697), .A2(new_n829), .A3(G330), .A4(new_n805), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT117), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT39), .B1(new_n880), .B2(new_n862), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT39), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1095), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n880), .A2(new_n862), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1098), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n892), .B1(new_n671), .B2(new_n805), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1106), .B(new_n1107), .C1(new_n1108), .C2(new_n828), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1101), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1105), .A2(new_n1109), .A3(new_n1101), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT118), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT118), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1105), .A2(new_n1109), .A3(new_n1116), .A4(new_n1101), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1102), .A2(new_n1113), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1094), .B1(new_n1118), .B2(new_n705), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n443), .A2(G330), .A3(new_n697), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n908), .A2(new_n1120), .A3(new_n624), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n694), .A2(new_n695), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n696), .A2(new_n499), .ZN(new_n1123));
  OAI211_X1 g0923(.A(G330), .B(new_n805), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n828), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT119), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n1108), .A4(new_n1101), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1108), .A3(new_n1101), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT119), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n893), .B1(new_n1125), .B2(new_n1101), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1121), .B(new_n1127), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1113), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1111), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n661), .B1(new_n1118), .B2(new_n1132), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1119), .B1(new_n1137), .B2(new_n1138), .ZN(G378));
  AOI21_X1  g0939(.A(new_n796), .B1(new_n261), .B2(new_n797), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n745), .A2(new_n299), .B1(new_n741), .B2(new_n764), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n713), .A2(G41), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G58), .C2(new_n779), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT122), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n748), .A2(new_n470), .B1(new_n750), .B2(new_n340), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT123), .Z(new_n1146));
  OAI221_X1 g0946(.A(new_n985), .B1(new_n772), .B2(new_n505), .C1(new_n345), .C2(new_n733), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT58), .Z(new_n1149));
  AOI211_X1 g0949(.A(G33), .B(G41), .C1(new_n760), .C2(G124), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n742), .B2(new_n728), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n748), .A2(new_n1077), .B1(new_n750), .B2(new_n788), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n732), .A2(G128), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n256), .B2(new_n735), .C1(new_n772), .C2(new_n1082), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n755), .C2(new_n1080), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1151), .B1(new_n1156), .B2(KEYINPUT59), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(KEYINPUT59), .B2(new_n1156), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1142), .B(new_n261), .C1(G33), .C2(G41), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT121), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1149), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n292), .A2(new_n640), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n296), .B(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1140), .B1(new_n726), .B2(new_n1161), .C1(new_n1165), .C2(new_n720), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n886), .B1(new_n881), .B2(new_n869), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n865), .B2(KEYINPUT40), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1165), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1167), .B(new_n1165), .C1(new_n865), .C2(KEYINPUT40), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1170), .A2(new_n907), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n907), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1166), .B1(new_n1174), .B2(new_n704), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1136), .A2(new_n1121), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1121), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1118), .B2(new_n1132), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n661), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1176), .B1(new_n1179), .B2(new_n1183), .ZN(G375));
  OAI21_X1  g0984(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1180), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n954), .A3(new_n1131), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1185), .A2(new_n704), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n706), .B1(G68), .B2(new_n1071), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n772), .A2(new_n528), .B1(new_n745), .B2(new_n470), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G283), .B2(new_n732), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n750), .A2(new_n345), .B1(new_n741), .B2(new_n773), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n276), .B(new_n1192), .C1(G116), .C2(new_n757), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n986), .A3(new_n1017), .A4(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n732), .A2(G137), .B1(new_n755), .B2(G159), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n261), .B2(new_n735), .C1(new_n1077), .C2(new_n772), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n712), .B1(G58), .B2(new_n779), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n757), .A2(new_n1080), .B1(new_n760), .B2(G128), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n256), .C2(new_n750), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1194), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1189), .B1(new_n1200), .B2(new_n722), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n829), .B2(new_n720), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1187), .A2(new_n1188), .A3(new_n1202), .ZN(G381));
  NAND3_X1  g1003(.A1(new_n1035), .A2(new_n1037), .A3(new_n770), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(G384), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(G390), .A2(G381), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n979), .A2(new_n998), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n971), .A2(new_n974), .A3(new_n972), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n974), .B1(new_n971), .B2(new_n972), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n699), .B1(new_n948), .B2(new_n950), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n704), .B1(new_n1211), .B2(new_n953), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1207), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1133), .B(new_n705), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1094), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n662), .B1(new_n1217), .B2(new_n1131), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1216), .B1(new_n1218), .B2(new_n1136), .ZN(new_n1219));
  INV_X1    g1019(.A(G375), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1206), .A2(new_n1213), .A3(new_n1219), .A4(new_n1220), .ZN(G407));
  OR3_X1    g1021(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(G407), .A2(G213), .A3(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1024(.A(G213), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(G343), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(G2897), .ZN(new_n1227));
  OAI211_X1 g1027(.A(KEYINPUT125), .B(new_n806), .C1(new_n810), .C2(new_n811), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1188), .A2(new_n1228), .A3(new_n1202), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1186), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1185), .A2(KEYINPUT60), .A3(new_n1180), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1231), .A2(new_n661), .A3(new_n1131), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(G384), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1229), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1227), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1238), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1227), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1236), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G378), .B(new_n1176), .C1(new_n1179), .C2(new_n1183), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1181), .A2(new_n953), .A3(new_n1174), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1219), .B1(new_n1246), .B2(new_n1175), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1226), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1244), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1252), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1068), .B(KEYINPUT115), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G387), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G390), .A2(new_n1213), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n770), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(KEYINPUT126), .A3(new_n1204), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1204), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n1258), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1256), .A2(new_n1257), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1226), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1253), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1251), .A2(new_n1254), .A3(new_n1267), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1268), .A2(new_n1272), .A3(new_n1269), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1268), .B2(new_n1243), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1273), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1271), .B1(new_n1278), .B2(new_n1267), .ZN(G405));
  NAND2_X1  g1079(.A1(G375), .A2(new_n1219), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1245), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1253), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1269), .A2(new_n1280), .A3(new_n1245), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1267), .ZN(G402));
endmodule


