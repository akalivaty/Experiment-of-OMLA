//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933;
  XNOR2_X1  g000(.A(KEYINPUT68), .B(G128), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G146), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n187), .A2(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .A4(G128), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n199), .C2(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(G134), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(new_n202), .B2(G134), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n199), .A3(G137), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n204), .A2(new_n208), .A3(new_n209), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n199), .A2(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n199), .B2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n198), .A2(new_n213), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n205), .A2(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n209), .B1(new_n224), .B2(new_n204), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n204), .A2(new_n208), .A3(new_n212), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .A3(G131), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n221), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(G131), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n222), .A3(new_n213), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT69), .A3(new_n228), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n191), .A2(new_n192), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n235), .B2(new_n236), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n220), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(G116), .B(G119), .Z(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT28), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n232), .A2(KEYINPUT69), .A3(new_n228), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n232), .B2(new_n228), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n239), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AND4_X1   g062(.A1(KEYINPUT28), .A2(new_n248), .A3(new_n244), .A4(new_n219), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n240), .A2(new_n244), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n254));
  INV_X1    g068(.A(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n256), .B(new_n257), .Z(new_n258));
  NAND4_X1  g072(.A1(new_n250), .A2(KEYINPUT29), .A3(new_n251), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G902), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(KEYINPUT72), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n240), .A2(new_n244), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n248), .A2(KEYINPUT30), .A3(new_n219), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n232), .A2(new_n228), .A3(new_n239), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT30), .B1(new_n269), .B2(new_n219), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n243), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT70), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n268), .A2(new_n274), .A3(new_n243), .A4(new_n271), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n267), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(new_n258), .ZN(new_n277));
  INV_X1    g091(.A(new_n245), .ZN(new_n278));
  INV_X1    g092(.A(new_n249), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n269), .A2(new_n219), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n243), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n258), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n277), .A2(KEYINPUT29), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G472), .B1(new_n265), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n266), .A2(new_n258), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n273), .B2(new_n275), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n288), .A2(new_n289), .B1(new_n283), .B2(new_n282), .ZN(new_n290));
  INV_X1    g104(.A(new_n287), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n270), .B1(new_n240), .B2(KEYINPUT30), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n274), .B1(new_n292), .B2(new_n243), .ZN(new_n293));
  INV_X1    g107(.A(new_n275), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT31), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT71), .B1(new_n288), .B2(new_n289), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n290), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  NOR2_X1   g114(.A1(G472), .A2(G902), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n286), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G137), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT68), .B(G128), .Z(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT73), .A3(G119), .ZN(new_n310));
  INV_X1    g124(.A(G119), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G128), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n187), .B2(new_n311), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT24), .B(G110), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n309), .A2(KEYINPUT23), .A3(G119), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n311), .A2(G128), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(new_n312), .C1(KEYINPUT23), .C2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n317), .B1(G110), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT74), .A2(G125), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G146), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n326), .A2(new_n332), .A3(new_n190), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n321), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n321), .A2(KEYINPUT75), .A3(new_n330), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n324), .A2(new_n190), .A3(new_n328), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n315), .A2(new_n316), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n320), .A2(G110), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT76), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  INV_X1    g159(.A(new_n343), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n345), .B(new_n346), .C1(new_n336), .C2(new_n337), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n308), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n343), .A3(new_n307), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n260), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT25), .ZN(new_n351));
  INV_X1    g165(.A(G217), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(new_n260), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n348), .A2(new_n349), .A3(new_n354), .A4(new_n260), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n348), .A2(new_n349), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n353), .A2(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT77), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n356), .A2(KEYINPUT77), .A3(new_n359), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(new_n188), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G131), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n364), .B(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n209), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  MUX2_X1   g183(.A(new_n369), .B(new_n366), .S(KEYINPUT17), .Z(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n330), .A3(new_n339), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT18), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n367), .B1(new_n372), .B2(new_n209), .ZN(new_n373));
  INV_X1    g187(.A(new_n323), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n333), .B1(new_n374), .B2(new_n190), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n373), .B(new_n375), .C1(new_n372), .C2(new_n366), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT93), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT94), .B(G104), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n371), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n371), .B2(new_n377), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n260), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G475), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n326), .A2(new_n332), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n374), .B2(new_n386), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n369), .B(new_n330), .C1(G146), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n380), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(G475), .B1(new_n392), .B2(new_n381), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n260), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT20), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n393), .B2(new_n260), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n385), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G116), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G116), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT14), .A3(G122), .ZN(new_n404));
  INV_X1    g218(.A(new_n400), .ZN(new_n405));
  OAI211_X1 g219(.A(G107), .B(new_n404), .C1(new_n405), .C2(KEYINPUT14), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n187), .A2(new_n188), .ZN(new_n407));
  INV_X1    g221(.A(G128), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G143), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(new_n199), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n407), .A2(G134), .A3(new_n409), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n402), .B(new_n406), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n199), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n400), .B(new_n401), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n188), .A2(KEYINPUT13), .A3(G128), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT95), .ZN(new_n417));
  INV_X1    g231(.A(new_n409), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT13), .B1(new_n187), .B2(new_n188), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n414), .B(new_n415), .C1(new_n420), .C2(new_n199), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT9), .B(G234), .Z(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n424), .A2(new_n352), .A3(G953), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n413), .B2(new_n421), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n260), .ZN(new_n430));
  AND2_X1   g244(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n431));
  NOR2_X1   g245(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n432));
  OAI21_X1  g246(.A(G478), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n430), .B(new_n433), .Z(new_n434));
  NOR2_X1   g248(.A1(new_n399), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n437));
  XNOR2_X1  g251(.A(G104), .B(G107), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n255), .ZN(new_n439));
  INV_X1    g253(.A(G104), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT3), .B1(new_n440), .B2(G107), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n401), .A3(G104), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(G107), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n255), .A4(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n440), .A2(G107), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n401), .A2(G104), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT82), .B(G101), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n191), .A2(new_n192), .A3(G128), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n189), .A2(G128), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n450), .A2(new_n194), .B1(new_n451), .B2(new_n235), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n436), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n448), .A2(new_n445), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n235), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n195), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n454), .A2(KEYINPUT83), .A3(new_n456), .A4(new_n439), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n197), .A2(new_n449), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n230), .A2(new_n233), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT84), .B1(new_n460), .B2(KEYINPUT12), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n439), .A2(new_n445), .A3(new_n448), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT83), .B1(new_n462), .B2(new_n456), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n449), .A2(new_n452), .A3(new_n436), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n246), .B2(new_n247), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n465), .A2(KEYINPUT12), .A3(new_n228), .A4(new_n232), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n461), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT10), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n197), .A2(new_n449), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT80), .A3(G101), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT4), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n475), .B2(new_n445), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n239), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(KEYINPUT81), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(KEYINPUT81), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n473), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n234), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n458), .A2(new_n472), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n253), .A2(G227), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(G140), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT78), .B(G110), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n471), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n492));
  INV_X1    g306(.A(new_n485), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n471), .A2(new_n496), .A3(new_n485), .A4(new_n490), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n260), .ZN(new_n500));
  NAND2_X1  g314(.A1(G469), .A2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n471), .A2(new_n485), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n489), .B(KEYINPUT79), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n493), .A2(new_n494), .ZN(new_n505));
  OAI211_X1 g319(.A(G469), .B(new_n504), .C1(new_n505), .C2(new_n489), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G221), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n423), .B2(new_n260), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G952), .ZN(new_n511));
  AOI211_X1 g325(.A(G953), .B(new_n511), .C1(G234), .C2(G237), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT21), .B(G898), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n260), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G214), .B1(G237), .B2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n235), .A2(new_n236), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(new_n238), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G125), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n197), .A2(new_n331), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n521), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G224), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(G953), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(KEYINPUT7), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n526), .B2(new_n528), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT5), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n311), .A3(G116), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT86), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n541), .B(G113), .C1(new_n539), .C2(new_n241), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n241), .A2(new_n242), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n462), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n462), .B1(new_n542), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n533), .A2(new_n535), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT91), .A4(new_n547), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n243), .B1(new_n477), .B2(new_n478), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n544), .A3(new_n536), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n529), .B(new_n532), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n544), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n536), .B(KEYINPUT87), .Z(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n553), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT88), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n557), .A2(new_n556), .A3(new_n558), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n553), .B2(new_n559), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n555), .B(new_n562), .C1(new_n564), .C2(new_n561), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n260), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n554), .A2(new_n260), .A3(new_n565), .A4(new_n567), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n520), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND4_X1   g385(.A1(new_n435), .A2(new_n507), .A3(new_n510), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n304), .A2(new_n363), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  NAND2_X1  g388(.A1(new_n299), .A2(new_n260), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n575), .A2(G472), .B1(new_n301), .B2(new_n299), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n356), .A2(KEYINPUT77), .A3(new_n359), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n360), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n507), .A2(new_n510), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n427), .A2(KEYINPUT33), .A3(new_n428), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n422), .A2(KEYINPUT98), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT99), .A3(new_n425), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n422), .B2(new_n426), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n422), .B(KEYINPUT98), .C1(new_n585), .C2(new_n426), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n582), .B1(new_n588), .B2(KEYINPUT33), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G478), .ZN(new_n590));
  NAND2_X1  g404(.A1(G478), .A2(G902), .ZN(new_n591));
  INV_X1    g405(.A(G478), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n429), .A2(new_n592), .A3(new_n260), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT100), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n590), .A2(new_n596), .A3(new_n591), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n399), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n569), .A2(new_n602), .A3(new_n570), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n566), .A2(KEYINPUT97), .A3(new_n568), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n517), .A3(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n601), .A2(new_n516), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n581), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G104), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  INV_X1    g424(.A(new_n398), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n393), .A2(new_n260), .A3(new_n397), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n611), .A2(new_n612), .B1(G475), .B2(new_n384), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n434), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n605), .A2(new_n516), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n581), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  OR2_X1    g432(.A1(new_n344), .A2(new_n347), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n308), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n358), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n356), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n572), .A2(new_n576), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT37), .B(G110), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G12));
  NOR3_X1   g440(.A1(new_n580), .A2(new_n605), .A3(new_n614), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT102), .B(G900), .Z(new_n628));
  AOI21_X1  g442(.A(new_n512), .B1(new_n515), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n627), .A2(new_n304), .A3(new_n623), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n623), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n299), .A2(new_n301), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT32), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n634), .B1(new_n638), .B2(new_n286), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n639), .A2(KEYINPUT103), .A3(new_n627), .A4(new_n630), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  XNOR2_X1  g456(.A(new_n629), .B(KEYINPUT39), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n580), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT40), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n267), .A2(new_n258), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n251), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n276), .B2(new_n283), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n649));
  AOI21_X1  g463(.A(G902), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n636), .A2(new_n637), .B1(G472), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n623), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n569), .A2(new_n570), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n399), .A2(new_n434), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n645), .A2(new_n657), .A3(new_n518), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  NAND4_X1  g476(.A1(new_n399), .A2(new_n595), .A3(new_n597), .A4(new_n630), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT107), .ZN(new_n664));
  INV_X1    g478(.A(new_n605), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n304), .A2(new_n664), .A3(new_n665), .A4(new_n623), .ZN(new_n666));
  INV_X1    g480(.A(new_n580), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n190), .ZN(G48));
  AOI21_X1  g483(.A(new_n579), .B1(new_n638), .B2(new_n286), .ZN(new_n670));
  INV_X1    g484(.A(new_n500), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n499), .B1(new_n498), .B2(new_n260), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n671), .A2(new_n672), .A3(new_n509), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n670), .A2(new_n606), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT41), .B(G113), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NAND3_X1  g490(.A1(new_n670), .A2(new_n615), .A3(new_n673), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  NOR3_X1   g492(.A1(new_n399), .A2(new_n434), .A3(new_n516), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n639), .A2(new_n665), .A3(new_n673), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  NOR4_X1   g495(.A1(new_n671), .A2(new_n672), .A3(new_n509), .A4(new_n516), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n605), .A2(new_n658), .ZN(new_n683));
  INV_X1    g497(.A(new_n301), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n258), .B1(new_n250), .B2(new_n251), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n295), .B2(KEYINPUT31), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n288), .A2(new_n289), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n575), .B2(G472), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n356), .A2(new_n359), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(G472), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n299), .B2(new_n260), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n694), .A2(new_n690), .A3(new_n695), .A4(new_n688), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n682), .B(new_n683), .C1(new_n692), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  NAND3_X1  g512(.A1(new_n689), .A2(new_n623), .A3(new_n673), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n595), .A2(new_n597), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(KEYINPUT107), .A3(new_n399), .A4(new_n630), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n663), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n699), .A2(new_n605), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n331), .ZN(G27));
  AND3_X1   g520(.A1(new_n569), .A2(new_n570), .A3(new_n517), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n507), .A2(new_n510), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n507), .A2(new_n707), .A3(KEYINPUT109), .A4(new_n510), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n304), .A3(new_n363), .A4(new_n664), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n304), .A2(KEYINPUT42), .A3(new_n691), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n704), .B1(new_n710), .B2(new_n711), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n713), .A2(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n209), .ZN(G33));
  NAND3_X1  g532(.A1(new_n613), .A2(new_n434), .A3(new_n630), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n670), .A2(new_n721), .A3(new_n712), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n199), .ZN(G36));
  NAND2_X1  g538(.A1(new_n700), .A2(new_n599), .ZN(new_n725));
  NAND2_X1  g539(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n577), .A3(new_n623), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(KEYINPUT44), .A3(new_n577), .A4(new_n623), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n707), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n504), .B1(new_n505), .B2(new_n489), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G469), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT46), .B1(new_n739), .B2(new_n501), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n671), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n501), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n510), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n643), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n732), .A2(KEYINPUT112), .A3(new_n707), .A4(new_n733), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n736), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  INV_X1    g562(.A(new_n304), .ZN(new_n749));
  INV_X1    g563(.A(new_n707), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n704), .A2(new_n363), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n510), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT47), .B1(new_n743), .B2(new_n510), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n749), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  NAND2_X1  g569(.A1(new_n511), .A2(new_n253), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT118), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n652), .A2(new_n512), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n363), .A2(new_n673), .A3(new_n707), .ZN(new_n761));
  OR4_X1    g575(.A1(new_n399), .A2(new_n760), .A3(new_n700), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n692), .A2(new_n696), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n729), .A2(new_n512), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n673), .ZN(new_n766));
  OR3_X1    g580(.A1(new_n766), .A2(new_n517), .A3(new_n656), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n763), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n765), .A2(new_n673), .A3(new_n707), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n623), .A3(new_n689), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n759), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n752), .A2(new_n753), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n671), .A2(new_n672), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n509), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n750), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n764), .A2(new_n765), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n758), .B(KEYINPUT51), .C1(new_n774), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n771), .A2(new_n773), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n758), .A2(KEYINPUT51), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n705), .B1(new_n666), .B2(new_n667), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n658), .B(new_n605), .C1(KEYINPUT113), .C2(new_n629), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n629), .A2(KEYINPUT113), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n653), .A2(new_n788), .A3(new_n667), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n641), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n787), .A2(new_n641), .A3(KEYINPUT52), .A4(new_n790), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(KEYINPUT114), .A3(new_n792), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n507), .A2(new_n510), .A3(new_n571), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n435), .B1(new_n598), .B2(new_n399), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n363), .A2(new_n576), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n573), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n680), .A3(new_n624), .A4(new_n697), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n674), .A2(new_n677), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n712), .A2(new_n664), .A3(new_n689), .ZN(new_n805));
  INV_X1    g619(.A(new_n708), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n434), .A2(new_n629), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n304), .A2(new_n613), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n634), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n717), .A2(new_n809), .A3(new_n723), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n804), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n796), .A2(new_n797), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n793), .A2(new_n795), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n811), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT54), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n804), .A2(new_n810), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n793), .B2(new_n795), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n819), .B1(new_n821), .B2(KEYINPUT53), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n796), .A2(new_n811), .A3(KEYINPUT53), .A4(new_n797), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n816), .A2(KEYINPUT115), .A3(new_n813), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n749), .A2(new_n690), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n772), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT48), .Z(new_n830));
  OAI211_X1 g644(.A(G952), .B(new_n253), .C1(new_n766), .C2(new_n605), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n786), .A2(new_n818), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n760), .A2(new_n761), .A3(new_n601), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n757), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n776), .B(KEYINPUT49), .Z(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n690), .A3(new_n509), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n656), .A2(new_n725), .A3(new_n518), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n652), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n839), .ZN(G75));
  NAND2_X1  g654(.A1(new_n511), .A2(G953), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT119), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n825), .A2(G210), .A3(G902), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n562), .B1(new_n564), .B2(new_n561), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(new_n555), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT55), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n849), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n843), .B1(new_n850), .B2(new_n851), .ZN(G51));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n825), .A2(new_n853), .A3(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n853), .B1(new_n825), .B2(KEYINPUT54), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n854), .A2(new_n855), .A3(new_n826), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n501), .B(KEYINPUT57), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n498), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n825), .A2(G469), .A3(G902), .A4(new_n738), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n843), .B1(new_n858), .B2(new_n859), .ZN(G54));
  NAND4_X1  g674(.A1(new_n825), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n392), .A2(new_n381), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n861), .A2(new_n865), .A3(new_n863), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n861), .B2(new_n863), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n843), .B(new_n864), .C1(new_n866), .C2(new_n867), .ZN(G60));
  XOR2_X1   g682(.A(new_n591), .B(KEYINPUT59), .Z(new_n869));
  NOR3_X1   g683(.A1(new_n856), .A2(new_n589), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n827), .B2(new_n818), .ZN(new_n871));
  INV_X1    g685(.A(new_n589), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n842), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n870), .A2(new_n873), .ZN(G63));
  XNOR2_X1  g688(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n352), .A2(new_n260), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n825), .A2(new_n621), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n842), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n357), .B1(new_n825), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(G66));
  OAI21_X1  g697(.A(G953), .B1(new_n514), .B2(new_n530), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n804), .B2(G953), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n847), .B1(G898), .B2(new_n253), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(G69));
  XOR2_X1   g701(.A(new_n292), .B(new_n388), .Z(new_n888));
  AND2_X1   g702(.A1(new_n747), .A2(new_n754), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n745), .A2(new_n683), .A3(new_n828), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n717), .A2(new_n723), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT125), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n787), .A2(new_n641), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT124), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n253), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n253), .A2(G900), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n897), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n888), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n661), .A2(new_n895), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n644), .A2(new_n750), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n670), .A3(new_n799), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n889), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n888), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n253), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(G227), .A2(G900), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(G953), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n912), .B(new_n914), .ZN(G72));
  NOR2_X1   g729(.A1(new_n276), .A2(new_n283), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n906), .A2(new_n804), .A3(new_n889), .A4(new_n908), .ZN(new_n918));
  NAND2_X1  g732(.A1(G472), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT63), .Z(new_n920));
  AOI21_X1  g734(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n891), .A2(new_n896), .ZN(new_n924));
  INV_X1    g738(.A(new_n804), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n646), .B1(new_n293), .B2(new_n294), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n843), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n817), .A2(new_n917), .A3(new_n920), .A4(new_n927), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n922), .A2(new_n923), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT127), .B1(new_n932), .B2(new_n921), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(G57));
endmodule


