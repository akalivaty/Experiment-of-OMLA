//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT68), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n464), .A2(KEYINPUT69), .A3(new_n465), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G125), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT70), .A4(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n471), .B1(new_n483), .B2(G2105), .ZN(G160));
  INV_X1    g059(.A(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n464), .B2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT71), .Z(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n466), .B2(G136), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n488), .A2(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n473), .C2(new_n474), .ZN(new_n494));
  OR2_X1    g069(.A1(KEYINPUT72), .A2(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT72), .A2(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n485), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n485), .C1(new_n473), .C2(new_n474), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n485), .A2(G138), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n475), .A3(new_n476), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n501), .B2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT74), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n511), .A2(G88), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n520), .A2(G651), .B1(G50), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n514), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT75), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT7), .Z(new_n531));
  NOR2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n522), .A2(new_n534), .A3(new_n523), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(G543), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n511), .A2(new_n513), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n532), .A2(new_n537), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT77), .B(G90), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n536), .A2(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n542), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n552), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(G171));
  NAND2_X1  g129(.A1(new_n536), .A2(G43), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n548), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n511), .A2(new_n513), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n555), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT79), .Z(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n518), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n559), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n533), .A2(G53), .A3(G543), .A4(new_n535), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  NAND2_X1  g153(.A1(new_n536), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n511), .A2(G87), .A3(new_n513), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n511), .A2(G86), .A3(new_n513), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n518), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n518), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n533), .A2(G543), .A3(new_n535), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n592), .B1(new_n593), .B2(new_n594), .C1(new_n559), .C2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  AND3_X1   g175(.A1(G301), .A2(KEYINPUT81), .A3(G868), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n559), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n594), .A2(KEYINPUT82), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n594), .B2(KEYINPUT82), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n518), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n607), .A2(new_n609), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT81), .B1(G301), .B2(G868), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n601), .B1(new_n616), .B2(new_n617), .ZN(G284));
  AOI21_X1  g193(.A(new_n601), .B1(new_n616), .B2(new_n617), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n615), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g197(.A(new_n614), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n560), .A2(new_n615), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n614), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n486), .A2(G123), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n485), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(G135), .B2(new_n466), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n475), .A2(new_n476), .A3(new_n468), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(new_n636), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(KEYINPUT83), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(KEYINPUT83), .ZN(new_n642));
  OAI221_X1 g217(.A(new_n635), .B1(new_n636), .B2(new_n639), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT84), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n636), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2096), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(new_n685), .B(new_n684), .S(new_n677), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT86), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n688), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n691), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n674), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n689), .A2(new_n691), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n699), .A3(new_n673), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n697), .A2(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G24), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G290), .B2(G16), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n705), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n693), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n704), .A2(new_n705), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n710), .A2(G1986), .A3(new_n706), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n702), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n702), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G6), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G305), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT32), .B(G1981), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n702), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n702), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n717), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n717), .A2(new_n722), .A3(new_n729), .A4(new_n726), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT87), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT87), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(G25), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n486), .A2(G119), .ZN(new_n737));
  OR2_X1    g312(.A1(G95), .A2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(G2104), .C1(G107), .C2(new_n485), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G131), .B2(new_n466), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n736), .B1(new_n741), .B2(new_n735), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT88), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT35), .B(G1991), .Z(new_n744));
  XOR2_X1   g319(.A(new_n743), .B(new_n744), .Z(new_n745));
  NAND3_X1  g320(.A1(new_n728), .A2(new_n730), .A3(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(KEYINPUT90), .B(KEYINPUT36), .C1(new_n712), .C2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n748), .A2(new_n749), .A3(new_n711), .A4(new_n709), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G286), .A2(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n702), .A2(G21), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n731), .A2(G33), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n485), .A2(G103), .A3(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT92), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT25), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n466), .A2(G139), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n475), .A2(new_n476), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n761), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n760), .C1(new_n762), .C2(new_n485), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G2072), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n734), .A2(G27), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G164), .B2(new_n734), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n764), .A2(new_n765), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n754), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  AOI21_X1  g348(.A(KEYINPUT96), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND3_X1   g349(.A1(new_n772), .A2(KEYINPUT96), .A3(new_n773), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n755), .B(new_n771), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n702), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n734), .A2(G35), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT99), .Z(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G162), .B2(new_n734), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(KEYINPUT29), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(new_n783), .C1(G162), .C2(new_n734), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G2090), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n781), .B1(new_n789), .B2(KEYINPUT100), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n561), .A2(G16), .ZN(new_n791));
  OR2_X1    g366(.A1(G16), .A2(G19), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1341), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n788), .A2(G2090), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n734), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT91), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT28), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n466), .A2(G140), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n486), .A2(G128), .ZN(new_n801));
  OR2_X1    g376(.A1(G104), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G116), .C2(new_n485), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G29), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n797), .A2(new_n798), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n799), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT30), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n811), .A2(KEYINPUT94), .A3(G28), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n813));
  INV_X1    g388(.A(G28), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(KEYINPUT30), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n731), .B1(new_n811), .B2(G28), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n812), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n810), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n634), .B2(new_n735), .ZN(new_n821));
  NAND3_X1  g396(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT26), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n466), .A2(G141), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n486), .A2(G129), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n468), .A2(G105), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n731), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n731), .B2(G32), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT27), .B(G1996), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n821), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n794), .A2(new_n795), .A3(new_n809), .A4(new_n833), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n776), .A2(new_n790), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(G160), .A2(G29), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT24), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(G34), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(G34), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n734), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(G2084), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT98), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n623), .A2(G16), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G4), .B2(G16), .ZN(new_n844));
  INV_X1    g419(.A(G1348), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n836), .A2(G2084), .A3(new_n840), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n764), .A2(new_n765), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT93), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT93), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n846), .B(new_n847), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n702), .A2(G5), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G171), .B2(new_n702), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT97), .B(G1961), .Z(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n843), .B(G1348), .C1(G4), .C2(G16), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n854), .ZN(new_n857));
  INV_X1    g432(.A(G2090), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n785), .A2(KEYINPUT100), .A3(new_n858), .A4(new_n787), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n835), .A2(new_n842), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n751), .A2(KEYINPUT102), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT102), .B1(new_n751), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(G311));
  NAND2_X1  g440(.A1(new_n751), .A2(new_n862), .ZN(G150));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  INV_X1    g442(.A(G67), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n518), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G651), .ZN(new_n870));
  INV_X1    g445(.A(G55), .ZN(new_n871));
  INV_X1    g446(.A(G93), .ZN(new_n872));
  OAI221_X1 g447(.A(new_n870), .B1(new_n871), .B2(new_n594), .C1(new_n559), .C2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT103), .B(G860), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n623), .A2(G559), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT38), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n560), .A2(new_n873), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n560), .A2(new_n873), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n879), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT39), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n884), .A2(new_n885), .A3(new_n874), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(new_n884), .B2(new_n874), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n877), .B1(new_n886), .B2(new_n887), .ZN(G145));
  XNOR2_X1  g463(.A(new_n741), .B(KEYINPUT107), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n638), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n763), .B(new_n827), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n506), .A2(new_n501), .ZN(new_n893));
  INV_X1    g468(.A(new_n499), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n804), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n466), .A2(G142), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT105), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n486), .A2(G130), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n485), .A2(KEYINPUT106), .A3(G118), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT106), .B1(new_n485), .B2(G118), .ZN(new_n901));
  OR2_X1    g476(.A1(G106), .A2(G2105), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(G2104), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n896), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n890), .A2(new_n891), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n892), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n892), .B2(new_n906), .ZN(new_n908));
  XNOR2_X1  g483(.A(G160), .B(new_n634), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g490(.A(new_n882), .B(new_n627), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n614), .B(G299), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n614), .A2(G299), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n614), .A2(G299), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n916), .A2(new_n917), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n916), .A2(KEYINPUT108), .A3(new_n919), .A4(new_n922), .ZN(new_n927));
  AND4_X1   g502(.A1(KEYINPUT109), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(G290), .A2(new_n719), .ZN(new_n932));
  XNOR2_X1  g507(.A(G166), .B(G288), .ZN(new_n933));
  AOI21_X1  g508(.A(G305), .B1(new_n598), .B2(new_n599), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n935), .A2(KEYINPUT42), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT42), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n928), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  NOR4_X1   g515(.A1(new_n929), .A2(new_n937), .A3(new_n930), .A4(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n873), .A2(new_n615), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(G295));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n943), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n882), .A2(new_n553), .A3(new_n551), .ZN(new_n948));
  NAND3_X1  g523(.A1(G171), .A2(new_n881), .A3(new_n880), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(G286), .ZN(new_n951));
  INV_X1    g526(.A(new_n917), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(G168), .A3(new_n949), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n948), .A2(G168), .A3(new_n949), .ZN(new_n955));
  AOI21_X1  g530(.A(G168), .B1(new_n948), .B2(new_n949), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n919), .A2(new_n922), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n935), .A2(new_n936), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n954), .B(new_n960), .C1(new_n957), .C2(new_n958), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n947), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n951), .B2(new_n953), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n955), .A2(new_n956), .A3(new_n917), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n947), .A2(new_n967), .A3(new_n912), .A4(new_n963), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n946), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n912), .A3(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(new_n947), .A3(new_n963), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(new_n482), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n479), .B2(new_n480), .ZN(new_n976));
  OAI211_X1 g551(.A(G40), .B(new_n470), .C1(new_n976), .C2(new_n485), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(G164), .B2(G1384), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n828), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT110), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n741), .B(new_n744), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n804), .B(new_n808), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n981), .B2(new_n828), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n980), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n985), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(G290), .B(G1986), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n980), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n978), .A2(G1384), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT117), .B1(G164), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n895), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n979), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n773), .B1(new_n1000), .B2(new_n977), .ZN(new_n1001));
  INV_X1    g576(.A(new_n977), .ZN(new_n1002));
  INV_X1    g577(.A(G2084), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(G164), .B2(G1384), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n895), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n994), .B(G8), .C1(new_n1011), .C2(G286), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G286), .A2(G8), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1016), .B(new_n1013), .C1(new_n1001), .C2(new_n1010), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1012), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1011), .A2(G8), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(KEYINPUT51), .A3(new_n1013), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT62), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1014), .B(KEYINPUT122), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT62), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1020), .A4(new_n1012), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n583), .A2(new_n1026), .A3(new_n587), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n583), .B2(new_n587), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT113), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n895), .A2(new_n1006), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(G160), .A2(G40), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT113), .B(new_n1034), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1030), .A2(new_n1033), .A3(G8), .A4(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n579), .A2(G1976), .A3(new_n580), .A4(new_n581), .ZN(new_n1037));
  OAI211_X1 g612(.A(G8), .B(new_n1037), .C1(new_n977), .C2(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1033), .A2(G8), .A3(new_n1037), .A4(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1036), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(G164), .B2(new_n996), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n895), .A2(KEYINPUT111), .A3(new_n995), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n979), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n725), .B1(new_n1048), .B2(new_n977), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1002), .A2(new_n858), .A3(new_n1009), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1044), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1043), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1031), .A2(new_n1007), .ZN(new_n1058));
  NOR2_X1   g633(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT115), .B1(G164), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n895), .A2(new_n1062), .A3(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1002), .A2(new_n858), .A3(new_n1058), .A4(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1044), .B1(new_n1049), .B2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1066), .A2(KEYINPUT116), .A3(new_n1055), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT116), .B1(new_n1066), .B2(new_n1055), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1057), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NOR4_X1   g646(.A1(new_n1000), .A2(new_n977), .A3(new_n1071), .A4(G2078), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT123), .B(G1961), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n979), .A2(new_n1046), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n1002), .A3(new_n1047), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1071), .B1(new_n1077), .B2(G2078), .ZN(new_n1078));
  AOI21_X1  g653(.A(G301), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1022), .A2(new_n1025), .A3(new_n1070), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1033), .A2(G8), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1036), .A2(new_n1040), .A3(new_n714), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1027), .B(KEYINPUT114), .Z(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1044), .B(new_n1054), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1043), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1061), .A2(new_n1063), .B1(new_n1031), .B2(new_n1007), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1002), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n575), .B(KEYINPUT9), .Z(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n1091), .C2(new_n573), .ZN(new_n1092));
  OR2_X1    g667(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1093));
  NAND2_X1  g668(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n574), .A2(new_n576), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1076), .A2(new_n1002), .A3(new_n1047), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1090), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n845), .B1(new_n1100), .B2(new_n977), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1002), .A2(new_n808), .A3(new_n1032), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n623), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1956), .B1(new_n1087), .B2(new_n1002), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1097), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1048), .A2(new_n977), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT60), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n623), .B1(new_n1103), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n614), .A4(new_n1102), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1048), .A2(G1996), .A3(new_n977), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(G1341), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n1002), .B2(new_n1032), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n561), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT59), .B(new_n561), .C1(new_n1116), .C2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1109), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1115), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1099), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1090), .A2(new_n1096), .A3(KEYINPUT121), .A4(new_n1098), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1110), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G171), .B(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(G2105), .B1(new_n976), .B2(KEYINPUT124), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(KEYINPUT124), .B2(new_n976), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n470), .A2(KEYINPUT53), .A3(G40), .A4(new_n768), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1135), .A2(new_n1048), .A3(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1133), .A2(new_n1074), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1138), .A2(new_n1078), .B1(new_n1139), .B2(new_n1133), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1023), .A2(new_n1020), .A3(new_n1012), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1070), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1080), .B(new_n1086), .C1(new_n1131), .C2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1036), .A2(new_n1042), .A3(new_n1039), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1085), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1019), .A2(G286), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1049), .A2(new_n1065), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G8), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1149), .B2(new_n1054), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1145), .B(new_n1146), .C1(new_n1150), .C2(new_n1067), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1151), .A2(KEYINPUT118), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT118), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1155));
  AND4_X1   g730(.A1(KEYINPUT63), .A2(new_n1145), .A3(new_n1146), .A4(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n993), .B1(new_n1143), .B2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n980), .A2(new_n598), .A3(new_n693), .A4(new_n599), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1162));
  XNOR2_X1  g737(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT46), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n988), .A2(new_n828), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n982), .A2(new_n1165), .B1(new_n980), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(new_n983), .B2(KEYINPUT46), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n982), .A2(KEYINPUT125), .A3(new_n1165), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1167), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT47), .ZN(new_n1172));
  AND4_X1   g747(.A1(new_n744), .A2(new_n985), .A3(new_n741), .A4(new_n990), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n804), .A2(G2067), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n980), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1164), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1158), .A2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g752(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1179));
  AOI21_X1  g753(.A(new_n1179), .B1(new_n697), .B2(new_n700), .ZN(new_n1180));
  OAI211_X1 g754(.A(new_n914), .B(new_n1180), .C1(new_n964), .C2(new_n968), .ZN(G225));
  INV_X1    g755(.A(G225), .ZN(G308));
endmodule


