//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n468), .A2(G136), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT66), .Z(new_n485));
  AOI21_X1  g060(.A(new_n473), .B1(new_n466), .B2(new_n467), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n483), .B(new_n485), .C1(G124), .C2(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(new_n486), .A2(G126), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n473), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n466), .A2(new_n467), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n473), .A2(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n474), .A2(new_n496), .A3(G138), .A4(new_n473), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n506), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  INV_X1    g092(.A(G89), .ZN(new_n518));
  OAI221_X1 g093(.A(new_n516), .B1(new_n510), .B2(new_n517), .C1(new_n518), .C2(new_n508), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT67), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n501), .A2(new_n523), .A3(new_n502), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT68), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR3_X1    g102(.A1(new_n525), .A2(KEYINPUT68), .A3(new_n526), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(G168));
  INV_X1    g104(.A(new_n510), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n503), .A2(new_n507), .ZN(new_n531));
  AOI22_X1  g106(.A1(G52), .A2(new_n530), .B1(new_n531), .B2(G90), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n522), .A2(new_n524), .A3(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT69), .B1(new_n535), .B2(G651), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n537));
  AOI211_X1 g112(.A(new_n537), .B(new_n505), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n532), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G171));
  NAND3_X1  g115(.A1(new_n522), .A2(new_n524), .A3(G56), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n505), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n508), .A2(new_n544), .B1(new_n510), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT70), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n503), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n520), .A2(new_n521), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT72), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT71), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n510), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n507), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n564), .A2(new_n566), .B1(G91), .B2(new_n531), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n539), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g145(.A(KEYINPUT73), .B(new_n532), .C1(new_n536), .C2(new_n538), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  AOI22_X1  g149(.A1(G49), .A2(new_n530), .B1(new_n531), .B2(G87), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n522), .A2(new_n524), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n576), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G288));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n508), .A2(new_n579), .B1(new_n510), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n503), .A2(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT74), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n505), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n508), .A2(new_n588), .B1(new_n510), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n525), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n590), .B1(new_n593), .B2(G651), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  NAND3_X1  g173(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n508), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n599), .A2(new_n602), .B1(G54), .B2(new_n530), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n556), .B2(new_n558), .ZN(new_n605));
  AND2_X1   g180(.A1(G79), .A2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT76), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  MUX2_X1   g186(.A(G301), .B(new_n610), .S(new_n611), .Z(G284));
  MUX2_X1   g187(.A(G301), .B(new_n610), .S(new_n611), .Z(G321));
  NAND2_X1  g188(.A1(G299), .A2(new_n611), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G168), .B2(new_n611), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(G168), .B2(new_n611), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n609), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n547), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n611), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n610), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n474), .A2(new_n463), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT12), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT12), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n474), .A2(new_n626), .A3(new_n463), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n468), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n486), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n473), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(G14), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT77), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT78), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT79), .Z(new_n664));
  INV_X1    g239(.A(new_n658), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n660), .A3(new_n662), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n659), .A2(new_n661), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n662), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n658), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT80), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(new_n686), .B(new_n685), .S(new_n678), .Z(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  MUX2_X1   g275(.A(G23), .B(G288), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT33), .Z(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G1976), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT81), .B(G16), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G1971), .Z(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G6), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n586), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT82), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n703), .A2(new_n704), .A3(new_n709), .A4(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n706), .A2(G24), .ZN(new_n719));
  INV_X1    g294(.A(G290), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n706), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G1986), .Z(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G25), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n468), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n486), .A2(G119), .ZN(new_n726));
  OR2_X1    g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n723), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n717), .A2(new_n718), .A3(new_n722), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n723), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n723), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G2090), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT89), .B1(G29), .B2(G32), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n463), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT26), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n744), .B(new_n746), .C1(G141), .C2(new_n468), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n486), .A2(G129), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT88), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n723), .ZN(new_n751));
  MUX2_X1   g326(.A(new_n743), .B(KEYINPUT89), .S(new_n751), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n723), .A2(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT25), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G139), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n469), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n474), .A2(G127), .ZN(new_n761));
  NAND2_X1  g336(.A1(G115), .A2(G2104), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n473), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT87), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n755), .B1(new_n765), .B2(new_n723), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G2072), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n705), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n742), .A2(new_n754), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G164), .A2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G27), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G34), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n479), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2084), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n784), .A2(new_n723), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n637), .B2(new_n723), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n781), .B2(new_n782), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n774), .A2(new_n775), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n776), .A2(new_n783), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n741), .B2(G2090), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n705), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n547), .B2(new_n705), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1341), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n710), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n710), .ZN(new_n797));
  INV_X1    g372(.A(G1966), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n710), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n710), .ZN(new_n801));
  INV_X1    g376(.A(G1961), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n792), .A2(new_n795), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n609), .A2(new_n710), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G4), .B2(new_n710), .ZN(new_n806));
  INV_X1    g381(.A(G1348), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n723), .A2(G26), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT28), .Z(new_n811));
  NAND3_X1  g386(.A1(new_n474), .A2(G128), .A3(G2105), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT84), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n486), .A2(new_n814), .A3(G128), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n473), .A2(G116), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT85), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT85), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(G140), .B2(new_n468), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n816), .A2(new_n821), .A3(KEYINPUT86), .ZN(new_n822));
  AOI21_X1  g397(.A(KEYINPUT86), .B1(new_n816), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n811), .B1(new_n825), .B2(G29), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2067), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n808), .A2(new_n809), .A3(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n772), .A2(new_n804), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n736), .A2(new_n738), .A3(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n508), .A2(new_n832), .B1(new_n510), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n525), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n834), .B1(new_n837), .B2(G651), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT92), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n609), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT91), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT90), .B(KEYINPUT38), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n838), .A2(new_n547), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n839), .B2(new_n547), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n846), .B(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n840), .B1(new_n850), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n842), .B1(new_n851), .B2(new_n852), .ZN(G145));
  NAND2_X1  g428(.A1(new_n816), .A2(new_n821), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT86), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n816), .A2(new_n821), .A3(KEYINPUT86), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n495), .A2(new_n497), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n489), .A2(new_n490), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n486), .B2(G126), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(KEYINPUT93), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT93), .B1(new_n858), .B2(new_n860), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n856), .B(new_n857), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(new_n860), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n867), .B(new_n861), .C1(new_n822), .C2(new_n823), .ZN(new_n868));
  INV_X1    g443(.A(new_n750), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n864), .B2(new_n868), .ZN(new_n871));
  OAI22_X1  g446(.A1(new_n870), .A2(new_n871), .B1(new_n763), .B2(new_n760), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n864), .A2(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n750), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n765), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n730), .A2(new_n628), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n729), .A2(new_n625), .A3(new_n627), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n468), .A2(G142), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT94), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  INV_X1    g457(.A(G118), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(G2105), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(G130), .B2(new_n486), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n877), .A2(new_n878), .A3(new_n881), .A4(new_n885), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT95), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT95), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n872), .A2(new_n876), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n479), .B(new_n637), .ZN(new_n893));
  XOR2_X1   g468(.A(G162), .B(new_n893), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n872), .A2(new_n876), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n887), .A2(new_n888), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n897), .A3(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n896), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n892), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n891), .B1(new_n872), .B2(new_n876), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT97), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n891), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n874), .A2(new_n765), .A3(new_n875), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n764), .B1(new_n874), .B2(new_n875), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n892), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n915), .B2(new_n894), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n892), .A2(new_n895), .ZN(new_n917));
  AOI211_X1 g492(.A(KEYINPUT96), .B(new_n899), .C1(new_n872), .C2(new_n876), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n901), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT97), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g498(.A(new_n621), .B(new_n848), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n608), .A2(G299), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n603), .A2(new_n562), .A3(new_n607), .A4(new_n567), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT98), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT41), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n925), .A2(new_n930), .A3(new_n926), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n925), .B2(new_n926), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n924), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n927), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n924), .A2(new_n937), .ZN(new_n938));
  OR3_X1    g513(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT42), .ZN(new_n939));
  XNOR2_X1  g514(.A(G303), .B(G288), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G290), .A2(new_n586), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(G290), .A2(new_n586), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n940), .A3(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT42), .B1(new_n936), .B2(new_n938), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n939), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n939), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(G868), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G868), .B2(new_n839), .ZN(G295));
  OAI21_X1  g529(.A(new_n953), .B1(G868), .B2(new_n839), .ZN(G331));
  NAND3_X1  g530(.A1(new_n570), .A2(G168), .A3(new_n571), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT99), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n539), .B2(G168), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n570), .A2(new_n957), .A3(G168), .A4(new_n571), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n959), .A2(new_n848), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n848), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n934), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n849), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n959), .A2(new_n848), .A3(new_n960), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n937), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n967), .A3(new_n948), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT100), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n963), .A2(new_n967), .A3(new_n948), .A4(KEYINPUT100), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  INV_X1    g548(.A(new_n933), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n961), .B2(new_n962), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT101), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT101), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n974), .C1(new_n961), .C2(new_n962), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n967), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n973), .B1(new_n979), .B2(new_n949), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n970), .A2(new_n971), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n963), .A2(new_n967), .ZN(new_n983));
  AOI21_X1  g558(.A(G37), .B1(new_n983), .B2(new_n949), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT44), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n984), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT43), .B1(new_n979), .B2(new_n949), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n987), .A2(KEYINPUT43), .B1(new_n972), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(KEYINPUT44), .B2(new_n989), .ZN(G397));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n858), .B2(new_n860), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G40), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n471), .A2(new_n477), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n994), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n798), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n995), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1003), .A2(new_n1005), .A3(new_n782), .A4(new_n1000), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n992), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n991), .B1(new_n1007), .B2(G286), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G168), .A2(new_n992), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT122), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1007), .B2(KEYINPUT121), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1003), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1012), .A2(new_n782), .B1(new_n1001), .B2(new_n798), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n992), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1008), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1007), .A2(KEYINPUT51), .A3(new_n1009), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1016), .A2(KEYINPUT62), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT107), .B(KEYINPUT55), .Z(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(G303), .B(G8), .C1(KEYINPUT107), .C2(KEYINPUT55), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1023), .A2(KEYINPUT108), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT108), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT106), .B(G2090), .Z(new_n1028));
  NAND2_X1  g603(.A1(new_n1012), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n472), .A2(G40), .A3(new_n478), .ZN(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n865), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1032), .B2(new_n996), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n1031), .A4(new_n861), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1971), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT105), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1029), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT105), .B(G1971), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1027), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n995), .A2(new_n1000), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n575), .A2(new_n577), .A3(G1976), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(G8), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n582), .A2(new_n584), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G651), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n531), .A2(G86), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n530), .A2(G48), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(G1981), .B1(new_n581), .B2(new_n585), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n992), .B1(new_n995), .B2(new_n1000), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1050), .A3(KEYINPUT49), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT109), .B(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n1054), .A3(new_n1041), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1043), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT113), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1043), .A2(new_n1056), .A3(new_n1059), .A4(new_n1062), .ZN(new_n1063));
  AND4_X1   g638(.A1(new_n1000), .A2(new_n1003), .A3(new_n1005), .A4(new_n1028), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n1035), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1061), .A2(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1033), .A2(new_n1034), .A3(new_n775), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1003), .A2(new_n1005), .A3(new_n1000), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1068), .A2(new_n1069), .B1(new_n802), .B2(new_n1070), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n1001), .A2(new_n1069), .A3(G2078), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1073), .A2(KEYINPUT123), .A3(new_n572), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT123), .B1(new_n1073), .B2(new_n572), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1039), .B(new_n1067), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT62), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1019), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1040), .A2(G2067), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1070), .B2(new_n807), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(new_n608), .ZN(new_n1081));
  XOR2_X1   g656(.A(G299), .B(KEYINPUT57), .Z(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1070), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1033), .A2(new_n1034), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1082), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT116), .Z(new_n1093));
  AND2_X1   g668(.A1(new_n1080), .A2(new_n608), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT60), .B1(new_n1094), .B2(new_n1081), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(KEYINPUT61), .A3(new_n1087), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n608), .A2(KEYINPUT60), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1080), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT61), .B1(new_n1091), .B2(new_n1087), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT117), .B(G1996), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1033), .A2(new_n1034), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT118), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1033), .A2(new_n1034), .A3(new_n1106), .A4(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1040), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(KEYINPUT119), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT119), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n547), .B(new_n1102), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1101), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1113), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1111), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1102), .B1(new_n1117), .B2(new_n547), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1093), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1030), .A2(new_n1069), .A3(G2078), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n862), .A2(new_n863), .A3(G1384), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1034), .B(new_n1121), .C1(new_n1122), .C2(new_n997), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1071), .A2(G301), .A3(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT54), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1070), .A2(new_n802), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n1123), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT125), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1071), .A2(new_n1131), .A3(new_n1123), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(G171), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1071), .A2(G301), .A3(new_n1072), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(KEYINPUT54), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1014), .B1(new_n1013), .B2(new_n992), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1007), .A2(KEYINPUT121), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1010), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1017), .B1(new_n1138), .B2(new_n1008), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1067), .A2(new_n1039), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1126), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1078), .B1(new_n1119), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G288), .A2(G1976), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1056), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1049), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT111), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(KEYINPUT111), .A3(new_n1049), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1054), .B(KEYINPUT110), .Z(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1039), .B2(new_n1060), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1152), .A2(KEYINPUT112), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(KEYINPUT112), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1013), .A2(new_n992), .A3(G286), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1067), .A2(new_n1039), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT114), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT114), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1067), .A2(new_n1039), .A3(new_n1160), .A4(new_n1156), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1066), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(G8), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1060), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1039), .A2(KEYINPUT63), .A3(new_n1167), .A4(new_n1156), .ZN(new_n1168));
  OAI22_X1  g743(.A1(new_n1159), .A2(new_n1163), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1155), .A2(new_n1169), .A3(KEYINPUT115), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1168), .A2(new_n1166), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1173), .B2(new_n1158), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1143), .A2(new_n1170), .A3(new_n1176), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1122), .A2(new_n1030), .A3(new_n997), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1178), .A2(G1996), .A3(new_n750), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT104), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n824), .B(G2067), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(G1996), .B2(new_n750), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1181), .A2(new_n1182), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n730), .A2(new_n732), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n730), .A2(new_n732), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1178), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT103), .ZN(new_n1190));
  AND3_X1   g765(.A1(G290), .A2(new_n1190), .A3(G1986), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1178), .ZN(new_n1192));
  OR2_X1    g767(.A1(G290), .A2(G1986), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1190), .B1(G290), .B2(G1986), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1191), .B(new_n1192), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1177), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1192), .B1(new_n869), .B2(new_n1183), .ZN(new_n1198));
  OR3_X1    g773(.A1(new_n1192), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT46), .B1(new_n1192), .B2(G1996), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT47), .Z(new_n1202));
  NOR2_X1   g777(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1202), .B1(new_n1189), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n825), .A2(G2067), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1192), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1205), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1197), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g787(.A1(G227), .A2(new_n460), .ZN(new_n1214));
  AND3_X1   g788(.A1(new_n1214), .A2(new_n656), .A3(new_n699), .ZN(new_n1215));
  AND3_X1   g789(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g792(.A(KEYINPUT127), .B1(new_n989), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n1214), .A2(new_n699), .A3(new_n656), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1220), .B1(new_n910), .B2(new_n921), .ZN(new_n1221));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n1222));
  AND2_X1   g796(.A1(new_n972), .A2(new_n988), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n973), .B1(new_n982), .B2(new_n984), .ZN(new_n1224));
  OAI211_X1 g798(.A(new_n1221), .B(new_n1222), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AND2_X1   g799(.A1(new_n1219), .A2(new_n1225), .ZN(G308));
  NAND2_X1  g800(.A1(new_n1219), .A2(new_n1225), .ZN(G225));
endmodule


