//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1228, new_n1229, new_n1230, new_n1231;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n451));
  OR2_X1    g026(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n450), .A2(new_n451), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AND2_X1   g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n459), .A2(new_n460), .B1(G567), .B2(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT66), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n469), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G137), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n471), .A2(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g060(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G112), .B2(new_n472), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n479), .A2(G136), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND3_X1  g067(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(G114), .B2(new_n472), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n465), .A2(G138), .A3(new_n472), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n479), .A2(new_n500), .A3(G138), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n504));
  OAI211_X1 g079(.A(KEYINPUT69), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n505), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(KEYINPUT70), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n528), .B1(new_n519), .B2(new_n520), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n529), .A3(G543), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT71), .B(G51), .Z(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT7), .Z(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n514), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n521), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n514), .A2(G89), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n533), .A2(new_n538), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  OAI21_X1  g117(.A(G543), .B1(new_n503), .B2(new_n504), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(new_n512), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n521), .B1(new_n544), .B2(new_n505), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n527), .A2(new_n529), .A3(G543), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n545), .A2(G90), .B1(new_n546), .B2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n544), .B2(new_n505), .ZN(new_n549));
  AND2_X1   g124(.A1(G77), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AND2_X1   g128(.A1(new_n514), .A2(G56), .ZN(new_n554));
  AND2_X1   g129(.A1(G68), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT72), .B(G81), .Z(new_n557));
  NAND3_X1  g132(.A1(new_n514), .A2(new_n539), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n527), .A2(new_n529), .A3(G43), .A4(G543), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n544), .B2(new_n505), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT74), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n514), .A2(G65), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n574), .A2(new_n577), .A3(G651), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n546), .A2(new_n579), .A3(G53), .ZN(new_n580));
  INV_X1    g155(.A(G53), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT9), .B1(new_n530), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n580), .A2(new_n582), .B1(G91), .B2(new_n545), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(G299));
  NAND2_X1  g159(.A1(new_n545), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n546), .A2(G49), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n514), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n521), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n592), .A2(KEYINPUT75), .A3(G651), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n591), .B2(new_n516), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n590), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n516), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n546), .A2(G47), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n514), .A2(new_n539), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n530), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n514), .A2(G66), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n608), .B1(new_n611), .B2(G651), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n514), .A2(G92), .A3(new_n539), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n545), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n606), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n606), .B1(new_n619), .B2(G868), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(G299), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(G168), .ZN(G297));
  XOR2_X1   g199(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n465), .A2(new_n470), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n479), .A2(G135), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT77), .Z(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n639), .A2(new_n640), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n641), .A2(new_n643), .B1(new_n489), .B2(G123), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n635), .A2(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(G2096), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n636), .A2(new_n646), .A3(new_n647), .A4(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT80), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2451), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT81), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2454), .ZN(new_n667));
  INV_X1    g242(.A(new_n664), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n655), .A2(new_n668), .A3(new_n656), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G14), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n665), .B2(new_n669), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(KEYINPUT17), .A3(new_n677), .ZN(new_n682));
  INV_X1    g257(.A(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n689), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1956), .B(G2474), .Z(new_n700));
  XOR2_X1   g275(.A(G1961), .B(G1966), .Z(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(new_n703), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n699), .A2(new_n702), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT20), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n696), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(G1991), .B(G1996), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n708), .A2(new_n710), .A3(new_n696), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n712), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n695), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n718), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n720), .A2(new_n694), .A3(new_n716), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(G229));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G32), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n470), .A2(G105), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT26), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n726), .B(new_n728), .C1(G141), .C2(new_n479), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n489), .A2(G129), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT98), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n729), .A2(new_n731), .A3(KEYINPUT99), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n725), .B1(new_n737), .B2(new_n724), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT100), .Z(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n743), .B2(KEYINPUT24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT24), .B2(new_n743), .ZN(new_n745));
  INV_X1    g320(.A(G160), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n724), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT25), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n479), .A2(G139), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n465), .A2(G127), .ZN(new_n755));
  AND2_X1   g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  OAI21_X1  g331(.A(G2105), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT97), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n752), .B(new_n754), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n724), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n724), .B2(G33), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n749), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n750), .B2(new_n762), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n742), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT101), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT104), .B(KEYINPUT23), .ZN(new_n768));
  INV_X1    g343(.A(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n768), .B(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G35), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G162), .B2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT103), .B(KEYINPUT29), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2090), .ZN(new_n778));
  NAND2_X1  g353(.A1(G286), .A2(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n769), .A2(G21), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n778), .B1(G1966), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n747), .A2(new_n748), .ZN(new_n784));
  NOR2_X1   g359(.A1(G27), .A2(G29), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G164), .B2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n784), .B1(G2078), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n724), .A2(G26), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT96), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n489), .A2(G128), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n793));
  INV_X1    g368(.A(G116), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G2105), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G140), .B2(new_n479), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n786), .A2(G2078), .ZN(new_n801));
  INV_X1    g376(.A(G28), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT30), .ZN(new_n803));
  AOI21_X1  g378(.A(G29), .B1(new_n802), .B2(KEYINPUT30), .ZN(new_n804));
  OR2_X1    g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n801), .B(new_n807), .C1(new_n724), .C2(new_n645), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n787), .A2(new_n800), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G171), .A2(new_n769), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G5), .B2(new_n769), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  INV_X1    g387(.A(G1966), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n781), .ZN(new_n814));
  AND4_X1   g389(.A1(new_n773), .A2(new_n783), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G19), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n564), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G1341), .Z(new_n819));
  NOR2_X1   g394(.A1(G4), .A2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT93), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n618), .B2(new_n769), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n811), .A2(new_n812), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n824), .B(new_n826), .C1(new_n741), .C2(new_n739), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n767), .A2(new_n815), .A3(new_n819), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n769), .A2(G6), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n596), .B2(new_n769), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT89), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT32), .B(G1981), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n830), .A2(KEYINPUT89), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(KEYINPUT89), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n832), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n834), .A2(KEYINPUT90), .A3(new_n837), .ZN(new_n841));
  NOR2_X1   g416(.A1(G16), .A2(G23), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT91), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G288), .B2(new_n769), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT33), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1976), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n769), .A2(G22), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G166), .B2(new_n769), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1971), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n840), .A2(new_n841), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT34), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT34), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n840), .A2(new_n853), .A3(new_n841), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n724), .A2(G25), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n489), .A2(G119), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n472), .A2(G107), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n479), .A2(KEYINPUT86), .A3(G131), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT86), .B1(new_n479), .B2(G131), .ZN(new_n860));
  OAI221_X1 g435(.A(new_n856), .B1(new_n857), .B2(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT87), .Z(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n855), .B1(new_n863), .B2(new_n724), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT35), .B(G1991), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT88), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n864), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n769), .A2(G24), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n604), .B2(new_n769), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G1986), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n852), .A2(new_n854), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT36), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n852), .A2(new_n874), .A3(new_n854), .A4(new_n871), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n828), .B1(new_n876), .B2(new_n877), .ZN(G311));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  AND4_X1   g454(.A1(new_n767), .A2(new_n815), .A3(new_n819), .A4(new_n827), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(G150));
  NAND2_X1  g456(.A1(new_n619), .A2(G559), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n558), .A2(new_n560), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT73), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT106), .B(G93), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n514), .A2(new_n539), .A3(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n527), .A2(new_n529), .A3(G55), .A4(G543), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  INV_X1    g467(.A(G67), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n544), .B2(new_n505), .ZN(new_n894));
  AND2_X1   g469(.A1(G80), .A2(G543), .ZN(new_n895));
  OAI21_X1  g470(.A(G651), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n891), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(KEYINPUT105), .B(G651), .C1(new_n894), .C2(new_n895), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n887), .A2(new_n897), .A3(new_n556), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n895), .B1(new_n514), .B2(G67), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n892), .B1(new_n900), .B2(new_n516), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n889), .A2(new_n890), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n563), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n883), .B(new_n905), .Z(new_n906));
  AND2_X1   g481(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n907), .A2(new_n908), .A3(G860), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n903), .A2(G860), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT37), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n909), .A2(new_n911), .ZN(G145));
  XNOR2_X1  g487(.A(G160), .B(new_n491), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(new_n645), .Z(new_n914));
  NAND3_X1  g489(.A1(new_n759), .A2(KEYINPUT107), .A3(new_n760), .ZN(new_n915));
  INV_X1    g490(.A(new_n797), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n861), .B(new_n633), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n737), .A2(G164), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n479), .A2(G142), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n489), .A2(G130), .ZN(new_n927));
  OR2_X1    g502(.A1(G106), .A2(G2105), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G164), .B1(new_n734), .B2(new_n735), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n930), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n493), .A2(new_n496), .ZN(new_n935));
  INV_X1    g510(.A(new_n501), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n500), .B1(new_n479), .B2(G138), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n736), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n934), .B1(new_n939), .B2(new_n931), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n924), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n923), .A2(new_n921), .B1(new_n933), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n914), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n942), .A2(new_n943), .A3(new_n914), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g524(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n899), .B2(new_n904), .ZN(new_n952));
  OR3_X1    g527(.A1(new_n950), .A2(new_n952), .A3(new_n628), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT41), .ZN(new_n954));
  AND4_X1   g529(.A1(new_n578), .A2(new_n612), .A3(new_n583), .A4(new_n617), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n578), .A2(new_n583), .B1(new_n612), .B2(new_n617), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G299), .A2(new_n618), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n578), .A2(new_n612), .A3(new_n583), .A4(new_n617), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(KEYINPUT41), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n628), .B1(new_n950), .B2(new_n952), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n953), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n955), .A2(new_n956), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n953), .B2(new_n962), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n963), .A2(new_n965), .A3(KEYINPUT42), .ZN(new_n966));
  NAND2_X1  g541(.A1(G305), .A2(new_n604), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n596), .A2(G290), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(G303), .B(G288), .Z(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(G303), .B(G288), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n967), .A3(new_n968), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT42), .B1(new_n963), .B2(new_n965), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n966), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n966), .B2(new_n975), .ZN(new_n977));
  OAI21_X1  g552(.A(G868), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n903), .A2(new_n622), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(G295));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n979), .ZN(G331));
  NAND2_X1  g556(.A1(G301), .A2(G286), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n536), .B1(new_n544), .B2(new_n505), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n532), .A2(new_n983), .A3(new_n535), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n984), .A2(new_n540), .A3(new_n551), .A4(new_n547), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n556), .A2(new_n887), .B1(new_n897), .B2(new_n898), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n563), .A2(new_n903), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n982), .A2(new_n985), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n899), .A3(new_n904), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n964), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n904), .B2(new_n899), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(KEYINPUT109), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n990), .A2(new_n899), .A3(new_n995), .A4(new_n904), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n993), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n992), .B1(new_n997), .B2(new_n961), .ZN(new_n998));
  AOI21_X1  g573(.A(G37), .B1(new_n998), .B2(new_n974), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n971), .A2(new_n973), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(new_n992), .C1(new_n997), .C2(new_n961), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT43), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n989), .A2(new_n964), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n994), .B2(new_n996), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n961), .B1(new_n989), .B2(new_n991), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n974), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AND4_X1   g581(.A1(KEYINPUT43), .A2(new_n1006), .A3(new_n945), .A4(new_n1001), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT44), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n999), .B2(new_n1001), .ZN(new_n1011));
  AND4_X1   g586(.A1(new_n1010), .A2(new_n1006), .A3(new_n945), .A4(new_n1001), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1008), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(G397));
  NAND2_X1  g592(.A1(G303), .A2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n471), .A2(new_n482), .A3(G40), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n938), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G2090), .B1(new_n1028), .B2(KEYINPUT120), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n471), .A2(new_n482), .A3(G40), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G164), .A2(G1384), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1025), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n1023), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(G164), .B2(G1384), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n938), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1024), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1029), .A2(new_n1034), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT116), .B(G8), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1022), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1035), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1039), .A2(KEYINPUT114), .A3(new_n1035), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1023), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n938), .A2(new_n1026), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT115), .B1(new_n1050), .B2(KEYINPUT50), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1047), .B(new_n1032), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1046), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(G8), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1042), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1050), .A2(new_n1030), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1058), .A2(new_n1041), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G288), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1057), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1058), .A2(new_n1041), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(KEYINPUT117), .C1(new_n1060), .C2(G288), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1062), .B(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n593), .A2(new_n595), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n589), .A2(new_n521), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n592), .A2(G651), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1069), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G1981), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1059), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1068), .B1(new_n1071), .B2(new_n1069), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n596), .B2(new_n1068), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1079), .B2(KEYINPUT49), .ZN(new_n1080));
  AND4_X1   g655(.A1(new_n1077), .A2(new_n1070), .A3(KEYINPUT49), .A4(new_n1073), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT119), .B(new_n1076), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1070), .A2(KEYINPUT49), .A3(new_n1073), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT118), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1079), .A2(new_n1077), .A3(KEYINPUT49), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n1087), .B2(new_n1076), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1056), .B(new_n1066), .C1(new_n1083), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1039), .B2(G2078), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G301), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G2078), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(KEYINPUT122), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(KEYINPUT122), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT53), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1092), .A2(new_n1094), .B1(new_n1039), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1032), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n812), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1039), .A2(G2078), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(KEYINPUT53), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n812), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1039), .A2(G2078), .B1(KEYINPUT121), .B2(new_n1090), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1091), .A2(new_n1101), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G168), .A2(new_n1041), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT51), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n748), .B(new_n1032), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1039), .A2(new_n813), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1111), .B1(new_n1114), .B2(new_n1041), .ZN(new_n1115));
  AOI211_X1 g690(.A(G168), .B(new_n1041), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1116));
  INV_X1    g691(.A(G8), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT51), .B1(new_n1118), .B2(new_n1110), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1109), .B(new_n1115), .C1(new_n1116), .C2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT123), .B1(new_n1089), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1076), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1065), .B1(new_n1124), .B2(new_n1082), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1115), .B1(new_n1119), .B2(new_n1116), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1101), .A2(new_n1091), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1125), .A2(new_n1130), .A3(new_n1131), .A4(new_n1056), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G299), .B(KEYINPUT57), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1028), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1037), .A2(new_n1024), .A3(new_n1038), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n618), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1100), .A2(new_n823), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1058), .A2(new_n799), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1140), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1141), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(new_n1139), .A3(KEYINPUT61), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT58), .B(G1341), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1039), .A2(G1996), .B1(new_n1058), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n564), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT59), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1143), .A2(KEYINPUT60), .A3(new_n1144), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n618), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1148), .A2(new_n1150), .A3(new_n1154), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT60), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1155), .A2(new_n1158), .A3(new_n618), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1146), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1121), .A2(new_n1132), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n1114), .A2(G286), .A3(new_n1041), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1089), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1055), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1163), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1053), .A2(G8), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1022), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1125), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1126), .B(KEYINPUT62), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1089), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(G171), .A4(new_n1107), .ZN(new_n1173));
  NOR2_X1   g748(.A1(G288), .A2(G1976), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1070), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1176), .A2(new_n1063), .B1(new_n1125), .B2(new_n1165), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1161), .A2(new_n1170), .A3(new_n1173), .A4(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1037), .A2(new_n1030), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(G1996), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1180), .B1(new_n736), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1181), .B2(new_n736), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n797), .B(G2067), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT112), .B1(new_n1184), .B2(new_n1179), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1184), .A2(KEYINPUT112), .A3(new_n1179), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1183), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT113), .Z(new_n1188));
  INV_X1    g763(.A(new_n866), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n861), .B(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1188), .B1(new_n1180), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(G1986), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n604), .A2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT111), .Z(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1195), .B1(new_n1192), .B2(new_n604), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1191), .B1(new_n1179), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1178), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1179), .B1(new_n1184), .B2(new_n736), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT124), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT46), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  XOR2_X1   g778(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1204));
  XNOR2_X1  g779(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1194), .A2(new_n1179), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT48), .Z(new_n1207));
  OAI21_X1  g782(.A(new_n1205), .B1(new_n1191), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1188), .A2(new_n863), .A3(new_n1189), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n916), .A2(new_n799), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1180), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1198), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g788(.A1(new_n1006), .A2(new_n1001), .A3(new_n1010), .A4(new_n945), .ZN(new_n1215));
  AND2_X1   g789(.A1(new_n999), .A2(new_n1001), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1215), .B1(new_n1216), .B2(new_n1010), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1218));
  NOR2_X1   g792(.A1(G227), .A2(new_n463), .ZN(new_n1219));
  OAI21_X1  g793(.A(new_n1219), .B1(new_n671), .B2(new_n672), .ZN(new_n1220));
  OAI21_X1  g794(.A(new_n1218), .B1(G229), .B2(new_n1220), .ZN(new_n1221));
  NOR3_X1   g795(.A1(G401), .A2(new_n463), .A3(G227), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n1222), .A2(new_n722), .A3(KEYINPUT126), .ZN(new_n1223));
  AOI22_X1  g797(.A1(new_n1221), .A2(new_n1223), .B1(new_n946), .B2(new_n947), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n1217), .A2(new_n1224), .A3(KEYINPUT127), .ZN(new_n1225));
  AOI21_X1  g799(.A(KEYINPUT127), .B1(new_n1217), .B2(new_n1224), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
  NAND2_X1  g801(.A1(new_n1217), .A2(new_n1224), .ZN(new_n1228));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g804(.A1(new_n1217), .A2(new_n1224), .A3(KEYINPUT127), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n1230), .A2(new_n1231), .ZN(G225));
endmodule


