//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT74), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT74), .A3(G128), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n192), .A2(new_n194), .B1(G119), .B2(new_n191), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT24), .B(G110), .Z(new_n196));
  OR3_X1    g010(.A1(new_n195), .A2(KEYINPUT77), .A3(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT77), .B1(new_n195), .B2(new_n196), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT23), .B1(new_n191), .B2(G119), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT76), .B1(new_n191), .B2(G119), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n199), .B(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n197), .B(new_n198), .C1(G110), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(KEYINPUT16), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT64), .A2(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n202), .A2(new_n208), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n195), .A2(new_n196), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT75), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n201), .A2(G110), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n210), .B1(new_n221), .B2(new_n205), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n208), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G953), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(G221), .A3(G234), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT78), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(new_n230), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT79), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n231), .B2(new_n232), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n216), .A2(new_n224), .A3(new_n233), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n188), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n240), .A2(new_n241), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n189), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n238), .A2(new_n239), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n189), .A2(G902), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n246), .B(KEYINPUT80), .Z(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT32), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n226), .A3(G210), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT27), .Z(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G137), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  AOI22_X1  g075(.A1(KEYINPUT66), .A2(new_n261), .B1(new_n259), .B2(G137), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT11), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n260), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT11), .A2(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n269), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(G131), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n271), .ZN(new_n273));
  INV_X1    g087(.A(new_n260), .ZN(new_n274));
  OAI22_X1  g088(.A1(new_n263), .A2(KEYINPUT11), .B1(new_n269), .B2(G134), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G131), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT0), .B(G128), .ZN(new_n281));
  INV_X1    g095(.A(G143), .ZN(new_n282));
  INV_X1    g096(.A(new_n212), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT64), .A2(G146), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n282), .A2(G146), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n281), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n211), .A2(KEYINPUT65), .A3(G143), .A4(new_n212), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n283), .A2(new_n284), .A3(new_n282), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT65), .B1(new_n282), .B2(G146), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n280), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n269), .A2(G134), .ZN(new_n297));
  OAI21_X1  g111(.A(G131), .B1(new_n297), .B2(new_n260), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n211), .A2(G143), .A3(new_n212), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n191), .B1(new_n299), .B2(KEYINPUT1), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n286), .B1(new_n213), .B2(new_n282), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n299), .A2(new_n291), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(new_n289), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n298), .B(new_n279), .C1(new_n302), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G119), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT2), .B(G113), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n307), .A3(new_n311), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n258), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n256), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n296), .A2(new_n307), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n296), .B2(new_n307), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n312), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n256), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n314), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n323), .A3(new_n314), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT31), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT68), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n330), .A3(KEYINPUT31), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n326), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(G472), .A2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n251), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n318), .A2(new_n325), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n327), .A2(new_n330), .A3(KEYINPUT31), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n330), .B1(new_n327), .B2(KEYINPUT31), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n333), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT71), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n251), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(KEYINPUT32), .A3(new_n333), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n296), .A2(new_n307), .A3(new_n311), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n311), .B1(new_n296), .B2(new_n307), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n257), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n314), .A2(new_n316), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n323), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n308), .A2(KEYINPUT30), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n296), .A2(new_n307), .A3(new_n319), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n346), .B1(new_n354), .B2(new_n312), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n350), .B(new_n351), .C1(new_n355), .C2(new_n323), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n313), .A2(new_n314), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n317), .B1(new_n357), .B2(KEYINPUT28), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n256), .A2(new_n351), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n345), .B1(new_n361), .B2(G472), .ZN(new_n362));
  INV_X1    g176(.A(G472), .ZN(new_n363));
  AOI211_X1 g177(.A(KEYINPUT72), .B(new_n363), .C1(new_n356), .C2(new_n360), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n336), .A2(new_n343), .A3(new_n344), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT73), .ZN(new_n367));
  INV_X1    g181(.A(new_n362), .ZN(new_n368));
  INV_X1    g182(.A(new_n364), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n368), .A2(new_n369), .A3(new_n344), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT73), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n336), .A4(new_n343), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n250), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  OAI21_X1  g188(.A(G221), .B1(new_n374), .B2(G902), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G107), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G104), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OAI22_X1  g196(.A1(new_n379), .A2(new_n380), .B1(new_n382), .B2(G107), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n377), .A2(KEYINPUT82), .A3(KEYINPUT3), .A4(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n382), .A2(G107), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n378), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT85), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n392), .A3(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n302), .A2(new_n306), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n390), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n191), .B1(new_n287), .B2(KEYINPUT1), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n293), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n397), .B(new_n398), .C1(new_n306), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n306), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n293), .B2(new_n399), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n398), .B1(new_n404), .B2(new_n397), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n396), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT12), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n400), .A2(new_n306), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT84), .B1(new_n409), .B2(new_n390), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n410), .A2(new_n401), .B1(new_n394), .B2(new_n395), .ZN(new_n411));
  INV_X1    g225(.A(new_n280), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n402), .B2(new_n405), .ZN(new_n416));
  INV_X1    g230(.A(new_n395), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n391), .A2(KEYINPUT86), .A3(new_n393), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT86), .B1(new_n391), .B2(new_n393), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT10), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n381), .A2(new_n385), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT83), .A3(G101), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n424), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n295), .A3(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n416), .A2(new_n421), .A3(new_n412), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n414), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G140), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT81), .ZN(new_n431));
  INV_X1    g245(.A(G227), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G953), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n431), .B(new_n433), .Z(new_n434));
  NAND2_X1  g248(.A1(new_n417), .A2(KEYINPUT10), .ZN(new_n435));
  INV_X1    g249(.A(new_n420), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n436), .B2(new_n418), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT10), .B1(new_n410), .B2(new_n401), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n425), .A2(new_n295), .A3(new_n426), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n434), .B1(new_n440), .B2(new_n412), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n416), .A2(new_n421), .A3(new_n427), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n280), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n429), .A2(new_n434), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G469), .B1(new_n444), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  INV_X1    g260(.A(new_n434), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n428), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n407), .B2(new_n413), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n443), .B2(new_n428), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n446), .B(new_n188), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n376), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G214), .B1(G237), .B2(G902), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT87), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n226), .A2(G952), .ZN(new_n457));
  INV_X1    g271(.A(G234), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n252), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n188), .B(new_n226), .C1(G234), .C2(G237), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(G898), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G122), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT89), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n466), .B(KEYINPUT8), .Z(new_n467));
  INV_X1    g281(.A(new_n309), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n468), .A2(new_n310), .ZN(new_n469));
  INV_X1    g283(.A(G113), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT88), .B(KEYINPUT5), .Z(new_n471));
  AND2_X1   g285(.A1(new_n193), .A2(G116), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT5), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(new_n468), .ZN(new_n475));
  AND4_X1   g289(.A1(new_n469), .A2(new_n391), .A3(new_n393), .A4(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n468), .B2(new_n471), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n469), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n397), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n467), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G125), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n295), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n395), .A2(new_n482), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n226), .A2(G224), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT7), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n484), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(KEYINPUT7), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(KEYINPUT90), .A3(new_n489), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n479), .B1(new_n419), .B2(new_n420), .ZN(new_n495));
  INV_X1    g309(.A(new_n466), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n425), .A2(new_n312), .A3(new_n426), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n478), .B1(new_n436), .B2(new_n418), .ZN(new_n501));
  INV_X1    g315(.A(new_n497), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n466), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n498), .A3(KEYINPUT6), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n488), .B(new_n485), .Z(new_n505));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n506), .B(new_n466), .C1(new_n501), .C2(new_n502), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n499), .A2(new_n500), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n500), .B1(new_n499), .B2(new_n508), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n456), .B(new_n464), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n374), .A2(new_n187), .A3(G953), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G122), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G116), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n377), .B1(new_n515), .B2(KEYINPUT14), .ZN(new_n516));
  XNOR2_X1  g330(.A(G116), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(G128), .B(G143), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT94), .ZN(new_n521));
  XNOR2_X1  g335(.A(G128), .B(G143), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n259), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n524), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G134), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n519), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(G128), .A3(new_n282), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n530), .B(G134), .C1(new_n520), .C2(new_n529), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n517), .B(new_n377), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n531), .A2(new_n525), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n513), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n525), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n518), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n525), .A3(new_n532), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n512), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n539), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n252), .A2(new_n226), .A3(G214), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n282), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT18), .A3(G131), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n215), .B1(new_n210), .B2(new_n206), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n544), .B(G143), .ZN(new_n548));
  NAND2_X1  g362(.A1(KEYINPUT18), .A2(G131), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(G131), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n278), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n545), .A2(KEYINPUT17), .A3(G131), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n222), .A3(new_n208), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n551), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G113), .B(G122), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(new_n382), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n560), .B(new_n551), .C1(new_n555), .C2(new_n557), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n188), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G475), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n206), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n206), .B1(KEYINPUT91), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT92), .B1(new_n572), .B2(new_n213), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n569), .A2(new_n574), .A3(new_n214), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n552), .A2(new_n553), .B1(G146), .B2(new_n207), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n567), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n563), .B1(new_n578), .B2(new_n560), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT20), .ZN(new_n580));
  NOR2_X1   g394(.A1(G475), .A2(G902), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n566), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n543), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n453), .A2(new_n511), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n373), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  OAI21_X1  g403(.A(G472), .B1(new_n332), .B2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n341), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n452), .A3(new_n249), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n528), .A2(new_n533), .A3(new_n513), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n512), .B1(new_n536), .B2(new_n537), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT33), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n534), .A2(new_n597), .A3(new_n538), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(G478), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n540), .A2(new_n188), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n539), .B2(new_n540), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n579), .A2(new_n581), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT20), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n606), .B2(new_n566), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT95), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n593), .A2(new_n511), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G104), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n566), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n565), .A2(KEYINPUT97), .A3(G475), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n606), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n543), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n593), .A2(new_n511), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT98), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G107), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  AOI21_X1  g436(.A(KEYINPUT36), .B1(new_n234), .B2(new_n236), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n225), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n247), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT99), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n627), .A3(new_n247), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n244), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n591), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n511), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n452), .A4(new_n585), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  NAND2_X1  g448(.A1(new_n367), .A2(new_n372), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n456), .B1(new_n509), .B2(new_n510), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n629), .ZN(new_n637));
  INV_X1    g451(.A(G900), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n461), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n459), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n453), .A2(new_n618), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n635), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  XNOR2_X1  g458(.A(new_n640), .B(KEYINPUT39), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n452), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n342), .B1(new_n341), .B2(new_n251), .ZN(new_n649));
  AOI211_X1 g463(.A(KEYINPUT71), .B(KEYINPUT32), .C1(new_n340), .C2(new_n333), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n344), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n355), .A2(new_n256), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n357), .A2(new_n323), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(G902), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n363), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n509), .ZN(new_n660));
  INV_X1    g474(.A(new_n510), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(KEYINPUT38), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT38), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n509), .B2(new_n510), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n244), .A2(new_n626), .A3(new_n628), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n543), .A2(new_n584), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n455), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n648), .A2(new_n659), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT100), .B(G143), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G45));
  NAND2_X1  g486(.A1(new_n607), .A2(new_n640), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n453), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n366), .A2(KEYINPUT73), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n371), .B1(new_n651), .B2(new_n370), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n637), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  NOR2_X1   g492(.A1(new_n511), .A2(new_n608), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n443), .A2(new_n428), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n680), .A2(new_n434), .B1(new_n441), .B2(new_n414), .ZN(new_n681));
  OAI21_X1  g495(.A(G469), .B1(new_n681), .B2(G902), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n451), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n684), .B(G469), .C1(new_n681), .C2(G902), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n679), .A2(new_n686), .A3(new_n375), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n373), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NOR2_X1   g504(.A1(new_n511), .A2(new_n618), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n686), .A3(new_n375), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n373), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  INV_X1    g508(.A(new_n686), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n376), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n586), .A2(new_n463), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n635), .A2(new_n696), .A3(new_n637), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  XNOR2_X1  g513(.A(new_n668), .B(KEYINPUT102), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n511), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n363), .B1(new_n340), .B2(new_n188), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n358), .A2(new_n323), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(new_n325), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n334), .B1(new_n704), .B2(new_n328), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n250), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n701), .A2(new_n686), .A3(new_n375), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  OR2_X1    g522(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n705), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n590), .A3(new_n667), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n590), .A3(KEYINPUT103), .A4(new_n667), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n376), .B(new_n636), .C1(new_n683), .C2(new_n685), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NOR3_X1   g534(.A1(new_n509), .A2(new_n510), .A3(new_n455), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n452), .A2(new_n710), .A3(new_n709), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n373), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n724));
  AOI21_X1  g538(.A(new_n250), .B1(new_n370), .B2(new_n335), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n722), .A2(KEYINPUT42), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n723), .A2(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n278), .ZN(G33));
  NAND4_X1  g542(.A1(new_n635), .A2(new_n249), .A3(new_n642), .A4(new_n721), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n584), .B2(new_n602), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n599), .A2(new_n601), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n606), .A3(new_n733), .A4(new_n566), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n629), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n591), .A3(KEYINPUT44), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n721), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n736), .B2(new_n591), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n443), .A2(new_n428), .A3(new_n447), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n412), .A2(new_n440), .B1(new_n407), .B2(new_n413), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n742), .B(KEYINPUT45), .C1(new_n743), .C2(new_n447), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n429), .A2(new_n434), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(KEYINPUT106), .A3(KEYINPUT45), .A4(new_n742), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  INV_X1    g563(.A(new_n742), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n447), .B1(new_n414), .B2(new_n428), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n746), .A2(G469), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n451), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n741), .A2(new_n759), .A3(new_n375), .A4(new_n645), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  XOR2_X1   g575(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT46), .B1(new_n753), .B2(new_n754), .ZN(new_n765));
  INV_X1    g579(.A(new_n451), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n763), .B1(new_n767), .B2(new_n376), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n249), .A2(new_n673), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n635), .A2(new_n739), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n759), .A2(new_n375), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  NAND2_X1  g588(.A1(new_n695), .A2(KEYINPUT49), .ZN(new_n775));
  INV_X1    g589(.A(new_n584), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n249), .A2(new_n456), .A3(new_n375), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT108), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n776), .A3(new_n732), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT109), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n666), .A2(new_n659), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n780), .B(new_n781), .C1(KEYINPUT49), .C2(new_n695), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n695), .A2(new_n459), .A3(new_n376), .A4(new_n739), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n651), .A3(new_n249), .A4(new_n658), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n584), .A3(new_n732), .ZN(new_n786));
  INV_X1    g600(.A(new_n735), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n706), .A2(new_n460), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n696), .A2(new_n789), .A3(new_n455), .A4(new_n665), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n715), .A2(new_n716), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n784), .A2(new_n793), .A3(new_n787), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n795));
  NAND2_X1  g609(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n768), .A2(new_n772), .B1(new_n376), .B2(new_n686), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n789), .A2(new_n721), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n783), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT51), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n784), .A2(new_n725), .A3(new_n787), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT48), .Z(new_n804));
  NAND2_X1  g618(.A1(new_n789), .A2(new_n718), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n457), .B(new_n805), .C1(new_n785), .C2(new_n608), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n783), .B(new_n808), .C1(new_n797), .C2(new_n800), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n802), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n636), .A2(new_n700), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n667), .A2(new_n641), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n452), .A2(KEYINPUT111), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT111), .B1(new_n452), .B2(new_n812), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n659), .B(new_n811), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n643), .A2(new_n677), .A3(new_n719), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n637), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n367), .B2(new_n372), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n820), .A2(new_n642), .B1(new_n718), .B2(new_n717), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(KEYINPUT52), .A3(new_n677), .A4(new_n815), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n667), .A2(new_n542), .A3(new_n617), .A4(new_n640), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n453), .A2(new_n739), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n635), .A2(new_n825), .B1(new_n793), .B2(new_n722), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n729), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(new_n729), .A3(KEYINPUT110), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n373), .B1(new_n687), .B2(new_n692), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n586), .B1(new_n776), .B2(new_n732), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n511), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n249), .A3(new_n452), .A4(new_n592), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n707), .A2(new_n835), .A3(new_n632), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n698), .A3(new_n836), .A4(new_n588), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n727), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n823), .A2(new_n831), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  INV_X1    g656(.A(new_n821), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n843), .B2(KEYINPUT52), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n823), .A2(new_n831), .A3(new_n838), .A4(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n841), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n840), .B1(new_n821), .B2(new_n817), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n823), .A2(new_n831), .A3(new_n838), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n842), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT112), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n841), .A2(new_n848), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n841), .A2(new_n842), .A3(new_n845), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n810), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT115), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n782), .B1(new_n856), .B2(new_n858), .ZN(G75));
  NAND2_X1  g673(.A1(new_n841), .A2(new_n845), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(G210), .A3(G902), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n504), .A2(new_n507), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(new_n505), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(new_n861), .B2(new_n862), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n226), .A2(G952), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G51));
  XOR2_X1   g683(.A(new_n754), .B(KEYINPUT57), .Z(new_n870));
  AOI21_X1  g684(.A(new_n842), .B1(new_n841), .B2(new_n845), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n846), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n450), .B2(new_n449), .ZN(new_n873));
  INV_X1    g687(.A(new_n753), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n860), .A2(G902), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n868), .B1(new_n873), .B2(new_n875), .ZN(G54));
  NAND2_X1  g690(.A1(KEYINPUT58), .A2(G475), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT116), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n860), .A2(G902), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n579), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n868), .ZN(G60));
  NAND2_X1  g697(.A1(new_n596), .A2(new_n598), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT117), .Z(new_n885));
  XNOR2_X1  g699(.A(new_n600), .B(KEYINPUT59), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n846), .B2(new_n871), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(KEYINPUT118), .B(new_n887), .C1(new_n846), .C2(new_n871), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n868), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n886), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n850), .A2(new_n855), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n885), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n892), .A2(new_n895), .ZN(G63));
  NAND2_X1  g710(.A1(G217), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT60), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n841), .B2(new_n845), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n624), .B(KEYINPUT119), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n868), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n901), .B(new_n902), .C1(new_n245), .C2(new_n899), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT61), .Z(G66));
  INV_X1    g718(.A(new_n462), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n226), .B1(new_n905), .B2(G224), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n837), .B2(new_n226), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n863), .B1(G898), .B2(new_n226), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n907), .B(new_n908), .Z(G69));
  NOR2_X1   g723(.A1(new_n767), .A2(new_n376), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n645), .A3(new_n725), .A4(new_n811), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n729), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n727), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n821), .A2(new_n760), .A3(new_n677), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n913), .A2(new_n916), .A3(new_n773), .A4(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n226), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n354), .B(new_n572), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(G900), .B2(G953), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n773), .A2(new_n760), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n670), .A2(new_n821), .A3(new_n677), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n646), .A2(new_n833), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n373), .A2(new_n721), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n670), .A2(new_n821), .A3(new_n935), .A4(new_n677), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n926), .A2(new_n928), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n226), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n922), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n924), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n432), .B2(new_n638), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT123), .Z(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n924), .A2(new_n939), .A3(new_n942), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(G72));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n947));
  XNOR2_X1  g761(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n363), .A2(new_n188), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n947), .B(new_n951), .C1(new_n937), .C2(new_n837), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n653), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n925), .B1(new_n933), .B2(new_n932), .ZN(new_n954));
  INV_X1    g768(.A(new_n837), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n954), .A2(new_n955), .A3(new_n936), .A4(new_n928), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n947), .B1(new_n956), .B2(new_n951), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT126), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n937), .B2(new_n837), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n653), .A4(new_n952), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n355), .A2(new_n256), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n851), .A2(new_n654), .A3(new_n964), .A4(new_n951), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n955), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n964), .B1(new_n970), .B2(new_n951), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n971), .B2(new_n868), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n950), .B1(new_n920), .B2(new_n955), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT127), .B(new_n902), .C1(new_n973), .C2(new_n964), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n966), .B1(new_n972), .B2(new_n974), .ZN(G57));
endmodule


