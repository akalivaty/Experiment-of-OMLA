

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785;

  NOR2_X1 U379 ( .A1(n526), .A2(n726), .ZN(n684) );
  NOR2_X1 U380 ( .A1(n529), .A2(n527), .ZN(n699) );
  OR2_X1 U381 ( .A1(n520), .A2(n530), .ZN(n728) );
  NAND2_X1 U382 ( .A1(n400), .A2(n402), .ZN(n726) );
  NOR2_X1 U383 ( .A1(n699), .A2(n701), .ZN(n715) );
  BUF_X1 U384 ( .A(n521), .Z(n729) );
  INV_X2 U385 ( .A(G953), .ZN(n778) );
  OR2_X2 U386 ( .A1(n650), .A2(n689), .ZN(n554) );
  XNOR2_X1 U387 ( .A(n758), .B(n462), .ZN(n485) );
  NAND2_X1 U388 ( .A1(n548), .A2(n395), .ZN(n394) );
  AND2_X1 U389 ( .A1(n569), .A2(n568), .ZN(n370) );
  XNOR2_X1 U390 ( .A(n726), .B(KEYINPUT6), .ZN(n584) );
  XNOR2_X1 U391 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U392 ( .A1(n398), .A2(n397), .ZN(n538) );
  NAND2_X1 U393 ( .A1(n396), .A2(n394), .ZN(n398) );
  AND2_X1 U394 ( .A1(n684), .A2(n357), .ZN(n397) );
  OR2_X1 U395 ( .A1(n638), .A2(n403), .ZN(n402) );
  AND2_X1 U396 ( .A1(n399), .A2(n361), .ZN(n400) );
  INV_X1 U397 ( .A(n520), .ZN(n385) );
  INV_X1 U398 ( .A(n530), .ZN(n392) );
  AND2_X1 U399 ( .A1(n628), .A2(n627), .ZN(n630) );
  XNOR2_X1 U400 ( .A(G146), .B(G125), .ZN(n473) );
  XNOR2_X1 U401 ( .A(n511), .B(n457), .ZN(n774) );
  XNOR2_X1 U402 ( .A(KEYINPUT4), .B(G131), .ZN(n457) );
  NAND2_X1 U403 ( .A1(n420), .A2(n383), .ZN(n382) );
  INV_X1 U404 ( .A(KEYINPUT24), .ZN(n470) );
  XNOR2_X1 U405 ( .A(G119), .B(G128), .ZN(n471) );
  XNOR2_X1 U406 ( .A(n498), .B(n474), .ZN(n775) );
  XNOR2_X1 U407 ( .A(KEYINPUT96), .B(KEYINPUT11), .ZN(n494) );
  XNOR2_X1 U408 ( .A(n473), .B(KEYINPUT10), .ZN(n498) );
  XNOR2_X1 U409 ( .A(G131), .B(G143), .ZN(n492) );
  XNOR2_X1 U410 ( .A(n774), .B(G146), .ZN(n393) );
  XNOR2_X1 U411 ( .A(G104), .B(G110), .ZN(n459) );
  NOR2_X1 U412 ( .A1(n728), .A2(n523), .ZN(n524) );
  XNOR2_X1 U413 ( .A(n425), .B(n424), .ZN(n504) );
  INV_X1 U414 ( .A(G475), .ZN(n424) );
  NOR2_X1 U415 ( .A1(n661), .A2(G902), .ZN(n425) );
  NOR2_X1 U416 ( .A1(n413), .A2(n729), .ZN(n412) );
  NOR2_X1 U417 ( .A1(n588), .A2(n416), .ZN(n413) );
  AND2_X1 U418 ( .A1(n588), .A2(n416), .ZN(n414) );
  NOR2_X1 U419 ( .A1(n536), .A2(n415), .ZN(n395) );
  INV_X1 U420 ( .A(n591), .ZN(n407) );
  NOR2_X1 U421 ( .A1(n591), .A2(n416), .ZN(n410) );
  NOR2_X1 U422 ( .A1(n652), .A2(n785), .ZN(n371) );
  INV_X1 U423 ( .A(KEYINPUT34), .ZN(n422) );
  XNOR2_X1 U424 ( .A(n467), .B(KEYINPUT21), .ZN(n720) );
  XOR2_X1 U425 ( .A(KEYINPUT5), .B(G137), .Z(n481) );
  INV_X1 U426 ( .A(n631), .ZN(n378) );
  XNOR2_X1 U427 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n441) );
  NOR2_X1 U428 ( .A1(n521), .A2(n391), .ZN(n390) );
  XNOR2_X1 U429 ( .A(G902), .B(KEYINPUT15), .ZN(n631) );
  NOR2_X1 U430 ( .A1(n584), .A2(n583), .ZN(n585) );
  AND2_X1 U431 ( .A1(n514), .A2(n403), .ZN(n401) );
  XNOR2_X1 U432 ( .A(n456), .B(n647), .ZN(n511) );
  NAND2_X1 U433 ( .A1(n379), .A2(n375), .ZN(n380) );
  NOR2_X1 U434 ( .A1(n777), .A2(n376), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n428), .B(n427), .ZN(n751) );
  INV_X1 U436 ( .A(KEYINPUT41), .ZN(n427) );
  NOR2_X1 U437 ( .A1(n713), .A2(n714), .ZN(n428) );
  XNOR2_X1 U438 ( .A(n423), .B(KEYINPUT35), .ZN(n542) );
  XNOR2_X1 U439 ( .A(n434), .B(n502), .ZN(n759) );
  XNOR2_X1 U440 ( .A(n775), .B(n386), .ZN(n655) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n472), .B(n469), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n426), .B(n499), .ZN(n661) );
  XNOR2_X1 U444 ( .A(n503), .B(n498), .ZN(n426) );
  BUF_X1 U445 ( .A(n672), .Z(n666) );
  XNOR2_X1 U446 ( .A(n463), .B(n368), .ZN(n367) );
  XNOR2_X1 U447 ( .A(n460), .B(n369), .ZN(n368) );
  AND2_X1 U448 ( .A1(n634), .A2(G953), .ZN(n679) );
  INV_X1 U449 ( .A(G140), .ZN(n645) );
  XNOR2_X1 U450 ( .A(n372), .B(KEYINPUT40), .ZN(n652) );
  AND2_X1 U451 ( .A1(n625), .A2(n699), .ZN(n372) );
  INV_X1 U452 ( .A(G122), .ZN(n653) );
  XNOR2_X1 U453 ( .A(n522), .B(n364), .ZN(n702) );
  XNOR2_X1 U454 ( .A(n525), .B(KEYINPUT94), .ZN(n526) );
  NAND2_X1 U455 ( .A1(n405), .A2(n412), .ZN(n404) );
  INV_X1 U456 ( .A(n394), .ZN(n651) );
  AND2_X1 U457 ( .A1(n447), .A2(G210), .ZN(n356) );
  XNOR2_X1 U458 ( .A(KEYINPUT79), .B(n715), .ZN(n357) );
  AND2_X1 U459 ( .A1(n589), .A2(n414), .ZN(n358) );
  OR2_X1 U460 ( .A1(n412), .A2(n591), .ZN(n359) );
  AND2_X1 U461 ( .A1(n374), .A2(n378), .ZN(n360) );
  INV_X1 U462 ( .A(n729), .ZN(n415) );
  NAND2_X1 U463 ( .A1(G902), .A2(G472), .ZN(n361) );
  AND2_X1 U464 ( .A1(n548), .A2(n729), .ZN(n362) );
  NOR2_X1 U465 ( .A1(n579), .A2(n523), .ZN(n363) );
  XOR2_X1 U466 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n364) );
  INV_X1 U467 ( .A(n590), .ZN(n416) );
  INV_X1 U468 ( .A(KEYINPUT2), .ZN(n376) );
  AND2_X1 U469 ( .A1(n421), .A2(n384), .ZN(n365) );
  XNOR2_X1 U470 ( .A(n393), .B(n367), .ZN(n667) );
  XNOR2_X1 U471 ( .A(n523), .B(KEYINPUT1), .ZN(n521) );
  INV_X1 U472 ( .A(n763), .ZN(n379) );
  NAND2_X1 U473 ( .A1(n382), .A2(n365), .ZN(n381) );
  NAND2_X1 U474 ( .A1(n381), .A2(n518), .ZN(n423) );
  NAND2_X1 U475 ( .A1(n366), .A2(n376), .ZN(n374) );
  XNOR2_X1 U476 ( .A(n630), .B(n629), .ZN(n366) );
  INV_X1 U477 ( .A(n474), .ZN(n369) );
  NAND2_X1 U478 ( .A1(n370), .A2(n710), .ZN(n573) );
  NAND2_X1 U479 ( .A1(n370), .A2(n593), .ZN(n644) );
  XNOR2_X1 U480 ( .A(n371), .B(n582), .ZN(n614) );
  NAND2_X1 U481 ( .A1(n764), .A2(n376), .ZN(n373) );
  NAND2_X1 U482 ( .A1(n360), .A2(n373), .ZN(n377) );
  NOR2_X1 U483 ( .A1(n763), .A2(n777), .ZN(n706) );
  NOR2_X4 U484 ( .A1(n708), .A2(n377), .ZN(n672) );
  XNOR2_X2 U485 ( .A(n380), .B(KEYINPUT75), .ZN(n708) );
  INV_X1 U486 ( .A(n491), .ZN(n383) );
  NAND2_X1 U487 ( .A1(n491), .A2(n422), .ZN(n384) );
  AND2_X1 U488 ( .A1(n520), .A2(n577), .ZN(n552) );
  NAND2_X1 U489 ( .A1(n385), .A2(n392), .ZN(n391) );
  NAND2_X1 U490 ( .A1(n505), .A2(G221), .ZN(n388) );
  XNOR2_X1 U491 ( .A(n390), .B(n389), .ZN(n488) );
  INV_X1 U492 ( .A(KEYINPUT103), .ZN(n389) );
  XNOR2_X1 U493 ( .A(n393), .B(n486), .ZN(n638) );
  NAND2_X1 U494 ( .A1(n357), .A2(n702), .ZN(n396) );
  XNOR2_X2 U495 ( .A(n534), .B(n533), .ZN(n548) );
  NAND2_X1 U496 ( .A1(n638), .A2(n401), .ZN(n399) );
  INV_X1 U497 ( .A(G472), .ZN(n403) );
  NOR2_X1 U498 ( .A1(n404), .A2(n358), .ZN(n704) );
  NAND2_X1 U499 ( .A1(n411), .A2(n590), .ZN(n405) );
  NAND2_X1 U500 ( .A1(n408), .A2(n406), .ZN(n605) );
  NAND2_X1 U501 ( .A1(n358), .A2(n407), .ZN(n406) );
  AND2_X1 U502 ( .A1(n409), .A2(n359), .ZN(n408) );
  NAND2_X1 U503 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U504 ( .A(n589), .ZN(n411) );
  NAND2_X1 U505 ( .A1(n673), .A2(n631), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n419), .B(n417), .ZN(n673) );
  XNOR2_X1 U507 ( .A(n418), .B(n442), .ZN(n417) );
  XNOR2_X1 U508 ( .A(n444), .B(n473), .ZN(n418) );
  XNOR2_X1 U509 ( .A(n759), .B(n485), .ZN(n419) );
  NOR2_X1 U510 ( .A1(n749), .A2(n422), .ZN(n420) );
  NAND2_X1 U511 ( .A1(n749), .A2(n422), .ZN(n421) );
  NAND2_X1 U512 ( .A1(n363), .A2(n751), .ZN(n581) );
  NAND2_X1 U513 ( .A1(n529), .A2(n528), .ZN(n713) );
  NOR2_X1 U514 ( .A1(n728), .A2(n729), .ZN(n429) );
  AND2_X1 U515 ( .A1(n636), .A2(n635), .ZN(G63) );
  INV_X1 U516 ( .A(KEYINPUT101), .ZN(n537) );
  INV_X1 U517 ( .A(KEYINPUT74), .ZN(n629) );
  XNOR2_X1 U518 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U519 ( .A(KEYINPUT63), .ZN(n642) );
  BUF_X1 U520 ( .A(n542), .Z(n654) );
  XNOR2_X2 U521 ( .A(G122), .B(G113), .ZN(n432) );
  INV_X1 U522 ( .A(G104), .ZN(n431) );
  XNOR2_X2 U523 ( .A(n432), .B(n431), .ZN(n502) );
  XNOR2_X2 U524 ( .A(G116), .B(G107), .ZN(n509) );
  XNOR2_X1 U525 ( .A(KEYINPUT16), .B(G110), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n509), .B(n433), .ZN(n434) );
  XNOR2_X2 U527 ( .A(G119), .B(KEYINPUT3), .ZN(n436) );
  INV_X1 U528 ( .A(n436), .ZN(n435) );
  NAND2_X1 U529 ( .A1(KEYINPUT70), .A2(n435), .ZN(n439) );
  INV_X1 U530 ( .A(KEYINPUT70), .ZN(n437) );
  NAND2_X1 U531 ( .A1(n437), .A2(n436), .ZN(n438) );
  NAND2_X1 U532 ( .A1(n439), .A2(n438), .ZN(n758) );
  XNOR2_X1 U533 ( .A(KEYINPUT68), .B(G101), .ZN(n462) );
  NAND2_X1 U534 ( .A1(n778), .A2(G224), .ZN(n440) );
  XNOR2_X1 U535 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X2 U536 ( .A(G143), .B(G128), .ZN(n456) );
  XNOR2_X1 U537 ( .A(KEYINPUT18), .B(KEYINPUT89), .ZN(n443) );
  XNOR2_X1 U538 ( .A(n456), .B(n443), .ZN(n444) );
  INV_X1 U539 ( .A(G902), .ZN(n514) );
  INV_X1 U540 ( .A(G237), .ZN(n445) );
  NAND2_X1 U541 ( .A1(n514), .A2(n445), .ZN(n447) );
  XNOR2_X2 U542 ( .A(n446), .B(n356), .ZN(n622) );
  NAND2_X1 U543 ( .A1(n447), .A2(G214), .ZN(n709) );
  NAND2_X1 U544 ( .A1(n622), .A2(n709), .ZN(n448) );
  XNOR2_X1 U545 ( .A(n448), .B(KEYINPUT85), .ZN(n587) );
  XNOR2_X1 U546 ( .A(n587), .B(KEYINPUT19), .ZN(n594) );
  NOR2_X1 U547 ( .A1(G898), .A2(n778), .ZN(n449) );
  XNOR2_X1 U548 ( .A(KEYINPUT90), .B(n449), .ZN(n761) );
  NAND2_X1 U549 ( .A1(n761), .A2(G902), .ZN(n450) );
  NAND2_X1 U550 ( .A1(n778), .A2(G952), .ZN(n564) );
  NAND2_X1 U551 ( .A1(n450), .A2(n564), .ZN(n452) );
  NAND2_X1 U552 ( .A1(G237), .A2(G234), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n451), .B(KEYINPUT14), .ZN(n744) );
  NAND2_X1 U554 ( .A1(n452), .A2(n744), .ZN(n453) );
  OR2_X2 U555 ( .A1(n594), .A2(n453), .ZN(n455) );
  XNOR2_X1 U556 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n454) );
  XNOR2_X2 U557 ( .A(n455), .B(n454), .ZN(n532) );
  INV_X1 U558 ( .A(n532), .ZN(n491) );
  INV_X1 U559 ( .A(G134), .ZN(n647) );
  NAND2_X1 U560 ( .A1(n778), .A2(G227), .ZN(n458) );
  XNOR2_X1 U561 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U562 ( .A(n645), .B(G137), .ZN(n474) );
  XNOR2_X1 U563 ( .A(G107), .B(KEYINPUT76), .ZN(n461) );
  XNOR2_X1 U564 ( .A(n462), .B(n461), .ZN(n463) );
  OR2_X2 U565 ( .A1(n667), .A2(G902), .ZN(n465) );
  INV_X1 U566 ( .A(G469), .ZN(n464) );
  XNOR2_X2 U567 ( .A(n465), .B(n464), .ZN(n523) );
  NAND2_X1 U568 ( .A1(G234), .A2(n631), .ZN(n466) );
  XNOR2_X1 U569 ( .A(KEYINPUT20), .B(n466), .ZN(n475) );
  NAND2_X1 U570 ( .A1(G221), .A2(n475), .ZN(n467) );
  XNOR2_X1 U571 ( .A(n720), .B(KEYINPUT92), .ZN(n530) );
  NAND2_X1 U572 ( .A1(G234), .A2(n778), .ZN(n468) );
  XOR2_X1 U573 ( .A(KEYINPUT8), .B(n468), .Z(n505) );
  XOR2_X1 U574 ( .A(G110), .B(KEYINPUT23), .Z(n469) );
  NAND2_X1 U575 ( .A1(n655), .A2(n514), .ZN(n479) );
  XOR2_X1 U576 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n477) );
  NAND2_X1 U577 ( .A1(G217), .A2(n475), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U579 ( .A(n479), .B(n478), .ZN(n520) );
  XNOR2_X1 U580 ( .A(G113), .B(G116), .ZN(n480) );
  XNOR2_X1 U581 ( .A(n481), .B(n480), .ZN(n483) );
  NOR2_X1 U582 ( .A1(G953), .A2(G237), .ZN(n500) );
  NAND2_X1 U583 ( .A1(n500), .A2(G210), .ZN(n482) );
  XNOR2_X1 U584 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U586 ( .A(n584), .ZN(n487) );
  NAND2_X1 U587 ( .A1(n488), .A2(n487), .ZN(n490) );
  XNOR2_X1 U588 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n489) );
  XNOR2_X2 U589 ( .A(n490), .B(n489), .ZN(n749) );
  XOR2_X1 U590 ( .A(KEYINPUT12), .B(G140), .Z(n493) );
  XNOR2_X1 U591 ( .A(n493), .B(n492), .ZN(n497) );
  XOR2_X1 U592 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n495) );
  XNOR2_X1 U593 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U594 ( .A(n497), .B(n496), .Z(n499) );
  NAND2_X1 U595 ( .A1(G214), .A2(n500), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n504), .B(KEYINPUT13), .ZN(n529) );
  INV_X1 U598 ( .A(n529), .ZN(n517) );
  XOR2_X1 U599 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n507) );
  NAND2_X1 U600 ( .A1(G217), .A2(n505), .ZN(n506) );
  XNOR2_X1 U601 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U602 ( .A(n508), .B(KEYINPUT99), .Z(n513) );
  XNOR2_X1 U603 ( .A(n509), .B(n653), .ZN(n510) );
  XNOR2_X1 U604 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n632) );
  NAND2_X1 U606 ( .A1(n632), .A2(n514), .ZN(n516) );
  INV_X1 U607 ( .A(G478), .ZN(n515) );
  XNOR2_X1 U608 ( .A(n516), .B(n515), .ZN(n528) );
  INV_X1 U609 ( .A(n528), .ZN(n527) );
  NAND2_X1 U610 ( .A1(n517), .A2(n527), .ZN(n592) );
  INV_X1 U611 ( .A(n592), .ZN(n518) );
  NAND2_X1 U612 ( .A1(n542), .A2(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U613 ( .A(n519), .B(KEYINPUT84), .ZN(n540) );
  AND2_X1 U614 ( .A1(n429), .A2(n726), .ZN(n734) );
  NAND2_X1 U615 ( .A1(n532), .A2(n734), .ZN(n522) );
  XOR2_X1 U616 ( .A(KEYINPUT93), .B(n524), .Z(n569) );
  NAND2_X1 U617 ( .A1(n532), .A2(n569), .ZN(n525) );
  AND2_X1 U618 ( .A1(n529), .A2(n527), .ZN(n701) );
  NOR2_X1 U619 ( .A1(n713), .A2(n530), .ZN(n531) );
  NAND2_X1 U620 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U621 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n533) );
  INV_X1 U622 ( .A(KEYINPUT100), .ZN(n535) );
  XNOR2_X1 U623 ( .A(n520), .B(n535), .ZN(n722) );
  NAND2_X1 U624 ( .A1(n584), .A2(n722), .ZN(n536) );
  XNOR2_X1 U625 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U627 ( .A(n541), .B(KEYINPUT83), .ZN(n559) );
  OR2_X1 U628 ( .A1(n722), .A2(n729), .ZN(n544) );
  INV_X1 U629 ( .A(KEYINPUT102), .ZN(n543) );
  XNOR2_X1 U630 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U631 ( .A1(n545), .A2(n584), .ZN(n546) );
  XNOR2_X1 U632 ( .A(n546), .B(KEYINPUT77), .ZN(n547) );
  NAND2_X1 U633 ( .A1(n548), .A2(n547), .ZN(n551) );
  INV_X1 U634 ( .A(KEYINPUT64), .ZN(n549) );
  XNOR2_X1 U635 ( .A(n549), .B(KEYINPUT32), .ZN(n550) );
  XNOR2_X1 U636 ( .A(n551), .B(n550), .ZN(n650) );
  AND2_X1 U637 ( .A1(n362), .A2(n552), .ZN(n689) );
  NOR2_X1 U638 ( .A1(n654), .A2(n554), .ZN(n553) );
  OR2_X1 U639 ( .A1(n553), .A2(KEYINPUT44), .ZN(n557) );
  INV_X1 U640 ( .A(n554), .ZN(n555) );
  NAND2_X1 U641 ( .A1(n555), .A2(KEYINPUT44), .ZN(n556) );
  NAND2_X1 U642 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U643 ( .A1(n559), .A2(n558), .ZN(n561) );
  INV_X1 U644 ( .A(KEYINPUT45), .ZN(n560) );
  XNOR2_X2 U645 ( .A(n561), .B(n560), .ZN(n763) );
  NAND2_X1 U646 ( .A1(n726), .A2(n709), .ZN(n562) );
  XNOR2_X1 U647 ( .A(n562), .B(KEYINPUT30), .ZN(n567) );
  NOR2_X1 U648 ( .A1(G900), .A2(n778), .ZN(n563) );
  NAND2_X1 U649 ( .A1(n563), .A2(G902), .ZN(n565) );
  NAND2_X1 U650 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U651 ( .A1(n566), .A2(n744), .ZN(n574) );
  NOR2_X1 U652 ( .A1(n567), .A2(n574), .ZN(n568) );
  INV_X1 U653 ( .A(n622), .ZN(n570) );
  XOR2_X1 U654 ( .A(KEYINPUT73), .B(KEYINPUT38), .Z(n571) );
  XNOR2_X1 U655 ( .A(n570), .B(n571), .ZN(n710) );
  XNOR2_X1 U656 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n572) );
  XNOR2_X1 U657 ( .A(n573), .B(n572), .ZN(n625) );
  NAND2_X1 U658 ( .A1(n710), .A2(n709), .ZN(n714) );
  INV_X1 U659 ( .A(n726), .ZN(n577) );
  NOR2_X1 U660 ( .A1(n720), .A2(n574), .ZN(n575) );
  XOR2_X1 U661 ( .A(KEYINPUT69), .B(n575), .Z(n576) );
  NAND2_X1 U662 ( .A1(n520), .A2(n576), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n577), .A2(n583), .ZN(n578) );
  XOR2_X1 U664 ( .A(KEYINPUT28), .B(n578), .Z(n579) );
  XOR2_X1 U665 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n580) );
  XNOR2_X1 U666 ( .A(n581), .B(n580), .ZN(n785) );
  XNOR2_X1 U667 ( .A(KEYINPUT82), .B(KEYINPUT46), .ZN(n582) );
  XNOR2_X1 U668 ( .A(n585), .B(KEYINPUT104), .ZN(n586) );
  NAND2_X1 U669 ( .A1(n586), .A2(n699), .ZN(n618) );
  XNOR2_X1 U670 ( .A(n618), .B(KEYINPUT107), .ZN(n589) );
  BUF_X1 U671 ( .A(n587), .Z(n588) );
  XNOR2_X1 U672 ( .A(KEYINPUT108), .B(KEYINPUT36), .ZN(n590) );
  NOR2_X1 U673 ( .A1(KEYINPUT78), .A2(KEYINPUT47), .ZN(n591) );
  NOR2_X1 U674 ( .A1(n592), .A2(n570), .ZN(n593) );
  XOR2_X1 U675 ( .A(n644), .B(KEYINPUT80), .Z(n603) );
  BUF_X1 U676 ( .A(n594), .Z(n595) );
  INV_X1 U677 ( .A(n595), .ZN(n596) );
  NAND2_X1 U678 ( .A1(n363), .A2(n596), .ZN(n696) );
  NAND2_X1 U679 ( .A1(n715), .A2(KEYINPUT79), .ZN(n597) );
  NAND2_X1 U680 ( .A1(KEYINPUT78), .A2(n597), .ZN(n600) );
  OR2_X1 U681 ( .A1(n715), .A2(KEYINPUT79), .ZN(n598) );
  NOR2_X1 U682 ( .A1(KEYINPUT47), .A2(n598), .ZN(n599) );
  NOR2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n696), .A2(n601), .ZN(n602) );
  NOR2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n612) );
  INV_X1 U687 ( .A(n696), .ZN(n607) );
  INV_X1 U688 ( .A(KEYINPUT78), .ZN(n606) );
  NOR2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U690 ( .A1(n608), .A2(n715), .ZN(n610) );
  INV_X1 U691 ( .A(KEYINPUT47), .ZN(n609) );
  NOR2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n616) );
  INV_X1 U695 ( .A(KEYINPUT48), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n616), .B(n615), .ZN(n628) );
  INV_X1 U697 ( .A(n709), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n619), .A2(n729), .ZN(n621) );
  XNOR2_X1 U700 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n620) );
  XNOR2_X1 U701 ( .A(n621), .B(n620), .ZN(n624) );
  BUF_X1 U702 ( .A(n622), .Z(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n646) );
  INV_X1 U704 ( .A(n625), .ZN(n626) );
  INV_X1 U705 ( .A(n701), .ZN(n690) );
  NOR2_X1 U706 ( .A1(n626), .A2(n690), .ZN(n648) );
  NOR2_X1 U707 ( .A1(n646), .A2(n648), .ZN(n627) );
  INV_X1 U708 ( .A(n630), .ZN(n777) );
  NAND2_X1 U709 ( .A1(n666), .A2(G478), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n636) );
  INV_X1 U711 ( .A(G952), .ZN(n634) );
  INV_X1 U712 ( .A(n679), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n672), .A2(G472), .ZN(n640) );
  XNOR2_X1 U714 ( .A(KEYINPUT87), .B(KEYINPUT62), .ZN(n637) );
  XNOR2_X1 U715 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n641) );
  NOR2_X2 U717 ( .A1(n641), .A2(n679), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(G57) );
  XNOR2_X1 U719 ( .A(n644), .B(G143), .ZN(G45) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(G42) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(G36) );
  XOR2_X1 U722 ( .A(G119), .B(KEYINPUT126), .Z(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(G21) );
  XOR2_X1 U724 ( .A(G101), .B(n651), .Z(G3) );
  XOR2_X1 U725 ( .A(n652), .B(G131), .Z(G33) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(G24) );
  NAND2_X1 U727 ( .A1(n666), .A2(G217), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n655), .B(KEYINPUT121), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U730 ( .A1(n658), .A2(n679), .ZN(G66) );
  NAND2_X1 U731 ( .A1(n672), .A2(G475), .ZN(n663) );
  XOR2_X1 U732 ( .A(KEYINPUT66), .B(KEYINPUT88), .Z(n659) );
  XNOR2_X1 U733 ( .A(n659), .B(KEYINPUT59), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X2 U735 ( .A1(n664), .A2(n679), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n665), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U737 ( .A1(n666), .A2(G469), .ZN(n670) );
  XOR2_X1 U738 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n668) );
  XNOR2_X1 U739 ( .A(n667), .B(n668), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U741 ( .A1(n671), .A2(n679), .ZN(G54) );
  NAND2_X1 U742 ( .A1(n672), .A2(G210), .ZN(n678) );
  BUF_X1 U743 ( .A(n673), .Z(n674) );
  XNOR2_X1 U744 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n675), .B(KEYINPUT55), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n674), .B(n676), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n678), .B(n677), .ZN(n680) );
  NOR2_X2 U748 ( .A1(n680), .A2(n679), .ZN(n682) );
  XOR2_X1 U749 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n681) );
  XNOR2_X1 U750 ( .A(n682), .B(n681), .ZN(G51) );
  NAND2_X1 U751 ( .A1(n684), .A2(n699), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(G104), .ZN(G6) );
  XOR2_X1 U753 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n686) );
  NAND2_X1 U754 ( .A1(n684), .A2(n701), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n686), .B(n685), .ZN(n688) );
  XOR2_X1 U756 ( .A(G107), .B(KEYINPUT27), .Z(n687) );
  XNOR2_X1 U757 ( .A(n688), .B(n687), .ZN(G9) );
  XOR2_X1 U758 ( .A(G110), .B(n689), .Z(G12) );
  NOR2_X1 U759 ( .A1(n696), .A2(n690), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n692) );
  XNOR2_X1 U761 ( .A(G128), .B(KEYINPUT111), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n694), .B(n693), .ZN(G30) );
  INV_X1 U764 ( .A(n699), .ZN(n695) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U766 ( .A(KEYINPUT112), .B(n697), .Z(n698) );
  XNOR2_X1 U767 ( .A(G146), .B(n698), .ZN(G48) );
  NAND2_X1 U768 ( .A1(n702), .A2(n699), .ZN(n700) );
  XNOR2_X1 U769 ( .A(n700), .B(G113), .ZN(G15) );
  NAND2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n703), .B(G116), .ZN(G18) );
  XNOR2_X1 U772 ( .A(n704), .B(G125), .ZN(n705) );
  XNOR2_X1 U773 ( .A(n705), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U774 ( .A1(n706), .A2(KEYINPUT2), .ZN(n707) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n748) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT116), .ZN(n712) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U781 ( .A1(n718), .A2(n749), .ZN(n719) );
  XNOR2_X1 U782 ( .A(n719), .B(KEYINPUT117), .ZN(n740) );
  INV_X1 U783 ( .A(n720), .ZN(n721) );
  NOR2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U785 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n723) );
  XNOR2_X1 U786 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U787 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U788 ( .A(KEYINPUT114), .B(n727), .Z(n732) );
  NAND2_X1 U789 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U790 ( .A(KEYINPUT50), .B(n730), .Z(n731) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U792 ( .A(n733), .B(KEYINPUT115), .ZN(n736) );
  INV_X1 U793 ( .A(n734), .ZN(n735) );
  NAND2_X1 U794 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U795 ( .A(KEYINPUT51), .B(n737), .Z(n738) );
  NAND2_X1 U796 ( .A1(n738), .A2(n751), .ZN(n739) );
  NAND2_X1 U797 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U798 ( .A(n741), .B(KEYINPUT118), .ZN(n742) );
  XNOR2_X1 U799 ( .A(n742), .B(KEYINPUT52), .ZN(n743) );
  NAND2_X1 U800 ( .A1(n743), .A2(G952), .ZN(n746) );
  INV_X1 U801 ( .A(n744), .ZN(n745) );
  NOR2_X1 U802 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U803 ( .A1(n748), .A2(n747), .ZN(n754) );
  INV_X1 U804 ( .A(n749), .ZN(n750) );
  NAND2_X1 U805 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U806 ( .A(n752), .B(KEYINPUT119), .Z(n753) );
  NAND2_X1 U807 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U808 ( .A1(G953), .A2(n755), .ZN(n757) );
  XNOR2_X1 U809 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n756) );
  XNOR2_X1 U810 ( .A(n757), .B(n756), .ZN(G75) );
  XNOR2_X1 U811 ( .A(n758), .B(G101), .ZN(n760) );
  XNOR2_X1 U812 ( .A(n760), .B(n759), .ZN(n762) );
  NOR2_X1 U813 ( .A1(n762), .A2(n761), .ZN(n773) );
  XOR2_X1 U814 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n771) );
  BUF_X1 U815 ( .A(n763), .Z(n764) );
  NOR2_X1 U816 ( .A1(n764), .A2(G953), .ZN(n765) );
  XOR2_X1 U817 ( .A(KEYINPUT122), .B(n765), .Z(n769) );
  NAND2_X1 U818 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U819 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U820 ( .A1(n767), .A2(G898), .ZN(n768) );
  NAND2_X1 U821 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U822 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U823 ( .A(n773), .B(n772), .ZN(G69) );
  XNOR2_X1 U824 ( .A(n774), .B(KEYINPUT125), .ZN(n776) );
  XNOR2_X1 U825 ( .A(n776), .B(n775), .ZN(n780) );
  XNOR2_X1 U826 ( .A(n777), .B(n780), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n779), .A2(n778), .ZN(n784) );
  XNOR2_X1 U828 ( .A(n780), .B(G227), .ZN(n781) );
  NAND2_X1 U829 ( .A1(n781), .A2(G900), .ZN(n782) );
  NAND2_X1 U830 ( .A1(n782), .A2(G953), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n784), .A2(n783), .ZN(G72) );
  XOR2_X1 U832 ( .A(G137), .B(n785), .Z(G39) );
endmodule

