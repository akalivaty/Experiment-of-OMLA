//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226,
    new_n1227;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G137), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT66), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  AOI211_X1 g044(.A(new_n469), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR3_X1   g049(.A1(new_n468), .A2(new_n470), .A3(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(new_n467), .B2(G112), .ZN(new_n476));
  INV_X1    g051(.A(G100), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n467), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT68), .Z(new_n479));
  NAND2_X1  g054(.A1(new_n461), .A2(new_n463), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n467), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(KEYINPUT67), .A3(G136), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n479), .A2(new_n482), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NOR2_X1   g064(.A1(new_n460), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G102), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n471), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(new_n467), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n467), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n471), .A2(KEYINPUT4), .A3(G138), .A4(new_n467), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n501), .B(new_n503), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT69), .B(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n509), .A2(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G166));
  INV_X1    g091(.A(new_n513), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(new_n509), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(KEYINPUT70), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n508), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n527), .B2(new_n521), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n518), .B(new_n520), .C1(new_n524), .C2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n506), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n509), .A2(new_n533), .B1(new_n513), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n506), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n509), .A2(new_n539), .B1(new_n513), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(G78), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT72), .B1(new_n550), .B2(new_n500), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n552), .A2(G78), .A3(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n501), .A2(new_n503), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n551), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n517), .A2(G91), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n557), .A2(new_n558), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT73), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n556), .A2(G651), .B1(new_n517), .B2(G91), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n559), .B(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G166), .ZN(G303));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n509), .A2(new_n572), .B1(new_n513), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n577), .B(G651), .C1(new_n504), .C2(G74), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n554), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n509), .A2(new_n587), .B1(new_n513), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n583), .A2(KEYINPUT75), .A3(G651), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT76), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n586), .A2(new_n590), .A3(new_n594), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n554), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n509), .A2(new_n604), .B1(new_n513), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G290));
  INV_X1    g183(.A(G79), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT78), .B1(new_n609), .B2(new_n500), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT78), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n611), .A2(G79), .A3(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n610), .B(new_n612), .C1(new_n554), .C2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(new_n526), .B2(G54), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT10), .B1(new_n513), .B2(new_n616), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n513), .A2(KEYINPUT10), .A3(new_n616), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G171), .ZN(G284));
  OAI21_X1  g197(.A(new_n621), .B1(new_n620), .B2(G171), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT79), .Z(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(G868), .B2(new_n626), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(G868), .B2(new_n626), .ZN(G280));
  INV_X1    g203(.A(G860), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n619), .B1(G559), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT80), .ZN(G148));
  OR2_X1    g206(.A1(new_n619), .A2(G559), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n471), .A2(new_n490), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n481), .A2(G123), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n483), .A2(G135), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n481), .A2(KEYINPUT81), .A3(G123), .ZN(new_n646));
  NAND4_X1  g221(.A1(new_n642), .A2(new_n643), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(G2096), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n639), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2435), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2438), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2451), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2443), .B(G2446), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G14), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(KEYINPUT17), .B2(new_n674), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n670), .A2(new_n671), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n677), .B(new_n678), .C1(KEYINPUT17), .C2(new_n674), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n673), .B(KEYINPUT84), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n679), .C1(new_n678), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n649), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G2100), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n686), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n695), .B(new_n696), .C1(new_n694), .C2(new_n693), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  INV_X1    g275(.A(G1981), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n703), .B(new_n706), .ZN(G229));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G32), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n483), .A2(G141), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n481), .A2(G129), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n490), .A2(G105), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT26), .Z(new_n714));
  NAND4_X1  g289(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT89), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(new_n708), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT27), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1996), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n721), .A2(KEYINPUT23), .A3(G20), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n723));
  INV_X1    g298(.A(G20), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G16), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n725), .C1(new_n626), .C2(new_n721), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(G1956), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n542), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G19), .ZN(new_n729));
  INV_X1    g304(.A(G1341), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n721), .A2(G5), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G171), .B2(new_n721), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n729), .A2(new_n730), .B1(G1961), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(G1961), .ZN(new_n734));
  AND2_X1   g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  NOR2_X1   g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n735), .A2(new_n736), .A3(G29), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n471), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n469), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  INV_X1    g314(.A(G125), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n473), .B1(new_n480), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2105), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n466), .A2(KEYINPUT66), .A3(new_n467), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2084), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n733), .A2(new_n734), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n721), .A2(G4), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n721), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1348), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT90), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n708), .A2(G26), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n481), .A2(G128), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n483), .A2(G140), .ZN(new_n757));
  NOR2_X1   g332(.A1(G104), .A2(G2105), .ZN(new_n758));
  OAI21_X1  g333(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(G29), .ZN(new_n761));
  MUX2_X1   g336(.A(new_n755), .B(new_n761), .S(KEYINPUT28), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n727), .A2(new_n747), .A3(new_n754), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G28), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n766), .A2(new_n767), .A3(new_n708), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(new_n708), .B2(new_n647), .C1(new_n729), .C2(new_n730), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n708), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n708), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT91), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n721), .A2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G168), .B2(new_n721), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1966), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n764), .A2(new_n769), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n721), .A2(G23), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n579), .B2(new_n721), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT87), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n781), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G22), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G166), .B2(G16), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT88), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G1971), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n788), .A2(G1971), .A3(new_n789), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n784), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G305), .A2(new_n721), .ZN(new_n795));
  NOR2_X1   g370(.A1(G6), .A2(G16), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n795), .A2(KEYINPUT32), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT32), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n797), .A2(new_n701), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n701), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n794), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(KEYINPUT34), .B(new_n794), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n721), .A2(G24), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G290), .B2(G16), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(new_n705), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n705), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n708), .A2(G25), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n481), .A2(G119), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n483), .A2(G131), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n708), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT35), .B(G1991), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n808), .A2(new_n809), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n779), .B1(new_n805), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g398(.A(KEYINPUT36), .B(new_n821), .C1(new_n803), .C2(new_n804), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n720), .B(new_n778), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n490), .A2(G103), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT25), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n483), .A2(G139), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n827), .B(new_n828), .C1(new_n467), .C2(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G33), .B(new_n830), .S(G29), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2072), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n708), .A2(G35), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G162), .B2(new_n708), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G2090), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n825), .A2(new_n832), .A3(new_n837), .ZN(G311));
  OR3_X1    g413(.A1(new_n825), .A2(new_n832), .A3(new_n837), .ZN(G150));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n554), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G651), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT94), .B(G93), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n517), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n526), .A2(G55), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  OR2_X1    g426(.A1(new_n849), .A2(new_n542), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n542), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n749), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT95), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n629), .B1(new_n857), .B2(KEYINPUT39), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n744), .B(KEYINPUT96), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n488), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n647), .ZN(new_n865));
  INV_X1    g440(.A(new_n715), .ZN(new_n866));
  MUX2_X1   g441(.A(new_n716), .B(new_n866), .S(new_n830), .Z(new_n867));
  NAND2_X1  g442(.A1(G114), .A2(G2104), .ZN(new_n868));
  INV_X1    g443(.A(G126), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n480), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n870), .A2(G2105), .B1(G102), .B2(new_n490), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n496), .A2(new_n497), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n496), .B2(new_n497), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n760), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n867), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n481), .A2(G130), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n483), .A2(G142), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n637), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(new_n816), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n816), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n877), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n865), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(KEYINPUT98), .A3(new_n886), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n877), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT100), .B1(new_n877), .B2(new_n887), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n890), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT99), .B1(new_n877), .B2(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n895), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n877), .A2(new_n894), .A3(KEYINPUT99), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n865), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g479(.A1(new_n849), .A2(new_n620), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n854), .B(new_n632), .Z(new_n906));
  NAND3_X1  g481(.A1(G299), .A2(KEYINPUT101), .A3(new_n749), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n749), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n564), .A2(new_n568), .A3(new_n619), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n906), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n910), .A2(new_n911), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n913), .B2(new_n907), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n914), .B1(new_n906), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT42), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n593), .A2(G166), .A3(new_n595), .ZN(new_n922));
  AOI21_X1  g497(.A(G166), .B1(new_n593), .B2(new_n595), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n579), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n596), .A2(G303), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n593), .A2(G166), .A3(new_n595), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(G288), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n928));
  XNOR2_X1  g503(.A(G290), .B(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n924), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n924), .B2(new_n927), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n921), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n905), .B1(new_n933), .B2(new_n620), .ZN(G295));
  OAI21_X1  g509(.A(new_n905), .B1(new_n933), .B2(new_n620), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n930), .B2(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n924), .A2(new_n927), .ZN(new_n938));
  INV_X1    g513(.A(new_n929), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n924), .A2(new_n927), .A3(new_n929), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(KEYINPUT104), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n523), .B(KEYINPUT70), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(new_n518), .A3(G301), .A4(new_n520), .ZN(new_n945));
  NAND2_X1  g520(.A1(G286), .A2(G171), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n853), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n849), .A2(new_n542), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n852), .A2(new_n853), .A3(new_n946), .A4(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n918), .B2(new_n916), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n950), .A2(new_n951), .A3(new_n907), .A4(new_n913), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n943), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n932), .A2(new_n953), .A3(new_n954), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n957), .A2(new_n898), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n898), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n913), .A2(new_n917), .A3(new_n907), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT105), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n913), .A2(new_n907), .A3(new_n966), .A4(new_n917), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n952), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(KEYINPUT106), .A3(new_n952), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n954), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n962), .B1(new_n973), .B2(new_n943), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n961), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT44), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n960), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n943), .A2(new_n955), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n959), .B1(new_n980), .B2(new_n962), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n977), .A2(new_n978), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n978), .B1(new_n977), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(KEYINPUT127), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n875), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n739), .A2(new_n743), .A3(G40), .A4(new_n742), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT108), .Z(new_n993));
  INV_X1    g568(.A(G2067), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n760), .B(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n996), .B2(new_n866), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n992), .A2(G1996), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n993), .A2(new_n997), .B1(new_n717), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n815), .A2(new_n818), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n816), .A2(new_n819), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(G290), .B(new_n705), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(new_n992), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n875), .A2(new_n1006), .A3(new_n988), .ZN(new_n1007));
  INV_X1    g582(.A(G2090), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n988), .B1(new_n493), .B2(new_n498), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n991), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n990), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n875), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1971), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT55), .B(G8), .C1(new_n507), .C2(new_n515), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G166), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1020), .B(new_n1021), .C1(KEYINPUT55), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT45), .B(new_n988), .C1(new_n493), .C2(new_n498), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n498), .A2(KEYINPUT97), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n496), .A2(new_n497), .A3(new_n872), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1030), .B2(new_n871), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n991), .B(new_n1027), .C1(new_n1031), .C2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(G1966), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G2084), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1007), .A2(new_n1035), .A3(new_n991), .A4(new_n1010), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1022), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1026), .A2(KEYINPUT63), .A3(G168), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n579), .A2(G1976), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT111), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n875), .A2(G160), .A3(G40), .A4(new_n988), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1041), .A2(new_n1042), .A3(G8), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n1041), .B2(G8), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1024), .B(G8), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n590), .A2(new_n584), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G1981), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n586), .A2(new_n590), .A3(new_n701), .A4(new_n591), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1053), .B(new_n1054), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT112), .B(G1976), .Z(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1040), .B(new_n1057), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1046), .A2(new_n1047), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n1038), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1059), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1016), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1022), .B1(new_n1062), .B2(new_n1011), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT63), .B1(new_n1063), .B2(new_n1024), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1037), .A2(G168), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1061), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1006), .B1(new_n875), .B2(new_n988), .ZN(new_n1069));
  OAI211_X1 g644(.A(G160), .B(G40), .C1(new_n1009), .C2(KEYINPUT50), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1071), .A2(new_n1008), .B1(new_n1072), .B2(new_n791), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1022), .B1(new_n1073), .B2(KEYINPUT113), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1069), .A2(new_n1070), .A3(G2090), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n1016), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1024), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1078), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1060), .B(new_n1068), .C1(new_n1079), .C2(KEYINPUT63), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1047), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1039), .B(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1041), .A2(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT110), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1041), .A2(new_n1042), .A3(G8), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1055), .B(new_n1058), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1976), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1055), .A2(new_n1091), .A3(new_n579), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1050), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1081), .A2(new_n1090), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(G286), .A2(G8), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1007), .A2(new_n991), .A3(new_n1010), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1035), .A2(new_n1100), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1096), .B(new_n1099), .C1(new_n1101), .C2(new_n1022), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1099), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1027), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n989), .A2(new_n990), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1036), .B1(new_n1105), .B2(G1966), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1103), .B(G8), .C1(new_n1106), .C2(G286), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(KEYINPUT121), .B(new_n1096), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1096), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT62), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1078), .A2(new_n1059), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1105), .A2(KEYINPUT53), .A3(new_n773), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1072), .B2(G2078), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1007), .A2(new_n991), .A3(new_n1010), .ZN(new_n1119));
  INV_X1    g694(.A(G1961), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1116), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(G171), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n1101), .B2(new_n1096), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1107), .A4(new_n1102), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1114), .A2(new_n1115), .A3(new_n1123), .A4(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1080), .A2(new_n1095), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1348), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1119), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n493), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1133));
  NOR4_X1   g708(.A1(new_n1133), .A2(new_n990), .A3(G1384), .A4(G2067), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT115), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1041), .B2(G2067), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n619), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(KEYINPUT120), .B(new_n619), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1131), .A2(new_n1119), .B1(new_n1134), .B2(KEYINPUT115), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1137), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT120), .B1(new_n1148), .B2(new_n619), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1140), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1014), .A2(new_n1015), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1071), .B2(G1956), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n563), .B(KEYINPUT57), .Z(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1155), .B(new_n1153), .C1(new_n1071), .C2(G1956), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT61), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n542), .A2(KEYINPUT119), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1014), .A2(new_n1015), .A3(new_n996), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT117), .B(G1341), .Z(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT58), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1041), .A2(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1161), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1162), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1170), .B(new_n1160), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1159), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1157), .A2(KEYINPUT116), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT116), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1175));
  OAI211_X1 g750(.A(KEYINPUT61), .B(new_n1158), .C1(new_n1173), .C2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1146), .A2(new_n1151), .A3(new_n1172), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1138), .A2(new_n749), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1158), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1102), .B(new_n1107), .C1(new_n1112), .C2(new_n1109), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1025), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1121), .A2(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1186), .A2(new_n1118), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n989), .A2(new_n990), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1188), .A2(KEYINPUT53), .A3(new_n773), .A4(new_n1015), .ZN(new_n1189));
  XNOR2_X1  g764(.A(G171), .B(KEYINPUT54), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1119), .A2(KEYINPUT123), .A3(new_n1120), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1190), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1187), .A2(new_n1192), .B1(new_n1122), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1182), .A2(new_n1061), .A3(new_n1184), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(KEYINPUT124), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1115), .A2(new_n1197), .A3(new_n1182), .A4(new_n1194), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1181), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1005), .B1(new_n1130), .B2(new_n1199), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n992), .A2(G1986), .A3(G290), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT48), .Z(new_n1202));
  NAND2_X1  g777(.A1(new_n1003), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n993), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n760), .A2(G2067), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n999), .B2(new_n1000), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1203), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n995), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n993), .B1(new_n715), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n998), .B(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1213), .B(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1207), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1216), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n987), .B1(new_n1200), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1080), .A2(new_n1095), .A3(new_n1129), .ZN(new_n1219));
  AND2_X1   g794(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1219), .B1(new_n1181), .B2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g796(.A(KEYINPUT127), .B(new_n1216), .C1(new_n1221), .C2(new_n1005), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1218), .A2(new_n1222), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g798(.A1(new_n903), .A2(G319), .A3(new_n667), .ZN(new_n1225));
  NOR2_X1   g799(.A1(new_n1225), .A2(G229), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n979), .A2(new_n981), .ZN(new_n1227));
  NAND3_X1  g801(.A1(new_n1226), .A2(new_n683), .A3(new_n1227), .ZN(G225));
  INV_X1    g802(.A(G225), .ZN(G308));
endmodule


