//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n469), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n473), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n470), .A2(G136), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT66), .Z(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n464), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n474), .B1(new_n468), .B2(new_n469), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n483), .A2(new_n485), .B1(G124), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n474), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT69), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT68), .A2(KEYINPUT4), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT68), .A2(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n470), .A2(new_n495), .A3(G138), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  MUX2_X1   g076(.A(G102), .B(G114), .S(G2105), .Z(new_n502));
  AOI22_X1  g077(.A1(G126), .A2(new_n486), .B1(new_n502), .B2(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n511), .A2(KEYINPUT72), .A3(new_n512), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n512), .A2(G543), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n519), .A2(KEYINPUT70), .A3(G50), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT70), .B1(new_n519), .B2(G50), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  AND3_X1   g102(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n528));
  AOI211_X1 g103(.A(new_n527), .B(new_n528), .C1(G51), .C2(new_n519), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n517), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n519), .A2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(new_n516), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n533), .B1(new_n522), .B2(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n522), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n519), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n517), .A2(G81), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n519), .A2(G53), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n557), .A2(new_n558), .B1(new_n522), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n517), .A2(G91), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n560), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G166), .ZN(G303));
  OR2_X1    g139(.A1(new_n511), .A2(G74), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G49), .B2(new_n519), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n535), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n566), .B(KEYINPUT75), .C1(new_n567), .C2(new_n535), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n511), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G48), .B2(new_n519), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n515), .A2(G86), .A3(new_n516), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n522), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT76), .Z(new_n582));
  XOR2_X1   g157(.A(KEYINPUT78), .B(G85), .Z(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT77), .B(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n517), .A2(new_n583), .B1(new_n519), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(G290));
  NAND3_X1  g161(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n535), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n574), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n519), .A2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n591), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  NOR2_X1   g179(.A1(G286), .A2(new_n601), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n560), .A2(new_n561), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n601), .B2(new_n606), .ZN(G297));
  AOI21_X1  g182(.A(new_n605), .B1(new_n601), .B2(new_n606), .ZN(G280));
  AOI21_X1  g183(.A(new_n598), .B1(new_n587), .B2(new_n590), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NOR2_X1   g186(.A1(new_n548), .A2(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n600), .A2(G559), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n470), .A2(G2104), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  MUX2_X1   g196(.A(G99), .B(G111), .S(G2105), .Z(new_n622));
  AOI22_X1  g197(.A1(G123), .A2(new_n486), .B1(new_n622), .B2(G2104), .ZN(new_n623));
  INV_X1    g198(.A(G135), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n471), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(G156));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2427), .ZN(new_n631));
  INV_X1    g206(.A(G2430), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n640), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n641), .A2(G14), .A3(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  INV_X1    g225(.A(new_n646), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n647), .B1(new_n653), .B2(new_n644), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n645), .B2(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n645), .A2(new_n648), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n651), .B1(new_n656), .B2(KEYINPUT17), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n650), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT80), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  OR2_X1    g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n669), .B(new_n671), .C1(new_n664), .C2(new_n670), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT83), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT82), .ZN(new_n677));
  XOR2_X1   g252(.A(G1981), .B(G1986), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G24), .ZN(new_n682));
  XOR2_X1   g257(.A(G290), .B(KEYINPUT86), .Z(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G1986), .Z(new_n685));
  NOR2_X1   g260(.A1(G16), .A2(G22), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G166), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1971), .ZN(new_n688));
  NOR2_X1   g263(.A1(G6), .A2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G305), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(G16), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  MUX2_X1   g268(.A(G23), .B(new_n568), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  NOR3_X1   g271(.A1(new_n688), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT34), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n470), .A2(G131), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT84), .ZN(new_n701));
  MUX2_X1   g276(.A(G95), .B(G107), .S(G2105), .Z(new_n702));
  AOI22_X1  g277(.A1(G119), .A2(new_n486), .B1(new_n702), .B2(G2104), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT85), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n697), .A2(new_n698), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n685), .A2(new_n699), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT36), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G33), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n475), .A2(G127), .ZN(new_n714));
  NAND2_X1  g289(.A1(G115), .A2(G2104), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n474), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n465), .A2(G103), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT25), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n716), .B(new_n718), .C1(G139), .C2(new_n470), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT88), .Z(new_n720));
  AOI21_X1  g295(.A(new_n713), .B1(new_n720), .B2(G29), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2072), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT31), .B(G11), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n712), .B1(new_n724), .B2(G28), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT91), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(G28), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n725), .B2(KEYINPUT91), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n723), .B1(new_n726), .B2(new_n728), .C1(new_n625), .C2(new_n712), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G34), .ZN(new_n731));
  MUX2_X1   g306(.A(new_n731), .B(G160), .S(G29), .Z(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n712), .A2(G32), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n486), .A2(G129), .ZN(new_n736));
  INV_X1    g311(.A(G141), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n471), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT26), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n465), .A2(G105), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n735), .B1(new_n744), .B2(new_n712), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  OAI22_X1  g321(.A1(new_n745), .A2(new_n746), .B1(new_n733), .B2(new_n732), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g323(.A1(G27), .A2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G164), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AND4_X1   g327(.A1(new_n722), .A2(new_n734), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G16), .A2(G21), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G168), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT90), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1966), .ZN(new_n757));
  NOR2_X1   g332(.A1(G5), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G171), .B2(G16), .ZN(new_n759));
  INV_X1    g334(.A(G1961), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n753), .A2(KEYINPUT92), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT95), .B(KEYINPUT23), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n681), .A2(G20), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1956), .ZN(new_n767));
  NOR2_X1   g342(.A1(G4), .A2(G16), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n609), .B2(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G1348), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n712), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  MUX2_X1   g347(.A(G104), .B(G116), .S(G2105), .Z(new_n773));
  AOI22_X1  g348(.A1(G128), .A2(new_n486), .B1(new_n773), .B2(G2104), .ZN(new_n774));
  INV_X1    g349(.A(G140), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n471), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G29), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(KEYINPUT87), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(KEYINPUT87), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n767), .A2(new_n770), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n712), .A2(G35), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT93), .Z(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n488), .B2(G29), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2090), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G19), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n549), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1341), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n769), .A2(G1348), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n783), .A2(new_n790), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n762), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n753), .A2(new_n757), .A3(new_n761), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n711), .A2(new_n799), .ZN(G150));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n801));
  XNOR2_X1  g376(.A(G150), .B(new_n801), .ZN(G311));
  NAND2_X1  g377(.A1(new_n519), .A2(G55), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT97), .B(G93), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n803), .B1(new_n522), .B2(new_n804), .C1(new_n535), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G860), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT37), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n548), .B(new_n806), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n600), .A2(new_n610), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT98), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n812), .B2(KEYINPUT39), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n808), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT99), .ZN(G145));
  AOI22_X1  g393(.A1(G130), .A2(new_n486), .B1(new_n470), .B2(G142), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n820), .A2(new_n474), .A3(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n474), .B2(G118), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n617), .B(new_n824), .Z(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(new_n704), .Z(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT101), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n504), .B(new_n776), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n743), .ZN(new_n829));
  MUX2_X1   g404(.A(new_n720), .B(new_n719), .S(new_n829), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n827), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(G160), .B(new_n625), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G162), .ZN(new_n833));
  AOI21_X1  g408(.A(G37), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(KEYINPUT103), .Z(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n827), .B2(new_n830), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n830), .B(KEYINPUT102), .ZN(new_n837));
  INV_X1    g412(.A(new_n826), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g416(.A1(new_n806), .A2(G868), .ZN(new_n842));
  NAND2_X1  g417(.A1(G299), .A2(new_n600), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n606), .A2(new_n609), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT41), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n846), .A3(new_n844), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(new_n844), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT41), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n847), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n809), .B(new_n613), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n851), .B2(new_n854), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT42), .ZN(new_n857));
  OR2_X1    g432(.A1(G166), .A2(KEYINPUT105), .ZN(new_n858));
  NAND2_X1  g433(.A1(G166), .A2(KEYINPUT105), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n690), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(G305), .A3(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(G290), .B(new_n568), .Z(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n861), .A3(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n857), .B(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n842), .B1(new_n869), .B2(G868), .ZN(G295));
  AOI21_X1  g445(.A(new_n842), .B1(new_n869), .B2(G868), .ZN(G331));
  NAND3_X1  g446(.A1(new_n539), .A2(G286), .A3(new_n540), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G286), .B1(new_n539), .B2(new_n540), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n809), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(G171), .A2(G168), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n548), .A2(new_n806), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n548), .A2(new_n806), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n872), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n875), .A2(new_n879), .A3(new_n845), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n879), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n853), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n882), .B2(new_n868), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n866), .A2(new_n867), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n875), .A2(new_n879), .B1(new_n848), .B2(new_n852), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT43), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n853), .A2(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n875), .A2(new_n879), .A3(new_n845), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n868), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n882), .A2(KEYINPUT106), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n889), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n897), .B2(new_n884), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n887), .B1(new_n898), .B2(KEYINPUT43), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT107), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n883), .A2(new_n906), .A3(new_n886), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n900), .B1(new_n898), .B2(new_n903), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n894), .A2(new_n895), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT106), .B1(new_n888), .B2(new_n889), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n884), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n903), .A3(new_n883), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT44), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n916), .A2(new_n908), .A3(KEYINPUT108), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n901), .B1(new_n911), .B2(new_n917), .ZN(G397));
  INV_X1    g493(.A(G8), .ZN(new_n919));
  NOR2_X1   g494(.A1(G166), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT111), .ZN(new_n922));
  AOI21_X1  g497(.A(G1384), .B1(new_n501), .B2(new_n503), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT45), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n504), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT110), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(KEYINPUT45), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G40), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n473), .A2(new_n478), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n922), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1971), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n927), .A2(KEYINPUT110), .A3(new_n928), .ZN(new_n937));
  INV_X1    g512(.A(new_n930), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n924), .B1(new_n923), .B2(KEYINPUT45), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(KEYINPUT111), .A3(new_n933), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n943));
  XNOR2_X1  g518(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n934), .B1(new_n923), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n927), .B2(KEYINPUT50), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n923), .A2(KEYINPUT113), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n950), .A2(G2090), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n942), .A2(new_n943), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n952), .A2(G8), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n942), .A2(new_n951), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT114), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n921), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n957));
  INV_X1    g532(.A(G1981), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n577), .A2(new_n958), .A3(new_n578), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n577), .B2(new_n578), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n961), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n959), .A3(KEYINPUT49), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n919), .B1(new_n923), .B2(new_n933), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n570), .A2(new_n967), .A3(new_n571), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n566), .B(G1976), .C1(new_n567), .C2(new_n535), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n965), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n965), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n965), .B2(new_n970), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT52), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(KEYINPUT117), .B(KEYINPUT52), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT121), .B(G2084), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n950), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n927), .A2(new_n928), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n933), .A3(new_n930), .ZN(new_n984));
  INV_X1    g559(.A(G1966), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(G286), .A2(new_n919), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n980), .A2(KEYINPUT63), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n956), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n955), .A2(G8), .A3(new_n921), .A4(new_n952), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT115), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n953), .A2(new_n993), .A3(new_n921), .A4(new_n955), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n987), .A2(new_n988), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n980), .A2(new_n998), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT120), .B(new_n972), .C1(new_n978), .C2(new_n979), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n923), .A2(new_n948), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n933), .C1(new_n923), .C2(new_n944), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(KEYINPUT119), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(KEYINPUT119), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n789), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n919), .B1(new_n942), .B2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n999), .A2(new_n1000), .B1(new_n921), .B2(new_n1006), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n997), .B(new_n1007), .C1(new_n992), .C2(new_n994), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n996), .B1(new_n1008), .B2(KEYINPUT63), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n984), .A2(new_n1010), .A3(G2078), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n760), .B2(new_n950), .ZN(new_n1012));
  AOI21_X1  g587(.A(G2078), .B1(new_n935), .B2(new_n941), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT53), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G171), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n982), .A2(G168), .A3(new_n986), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT51), .ZN(new_n1019));
  AOI21_X1  g594(.A(G168), .B1(new_n982), .B2(new_n986), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  OAI211_X1 g596(.A(G8), .B(new_n1017), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1019), .A2(new_n1022), .A3(KEYINPUT62), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT62), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1016), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n606), .A2(KEYINPUT57), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n560), .B2(new_n561), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT56), .B(G2072), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n940), .A2(new_n933), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1956), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1002), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1029), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1348), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n950), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n923), .A2(new_n933), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G2067), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n600), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1031), .A2(new_n1033), .A3(new_n1029), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1034), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n609), .B(new_n1038), .C1(new_n950), .C2(new_n1035), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT60), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n600), .A2(KEYINPUT60), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1036), .A2(new_n1039), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n549), .A2(KEYINPUT122), .ZN(new_n1047));
  INV_X1    g622(.A(G1996), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n940), .A2(new_n1048), .A3(new_n933), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT58), .B(G1341), .Z(new_n1050));
  NAND2_X1  g625(.A1(new_n1037), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1047), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g629(.A(KEYINPUT59), .B(new_n1047), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1044), .B(new_n1046), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1031), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n1034), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1029), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(KEYINPUT61), .A3(new_n1041), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1042), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(G301), .B(new_n1012), .C1(new_n1013), .C2(KEYINPUT53), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1015), .A2(KEYINPUT54), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n931), .A2(new_n922), .A3(new_n934), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT111), .B1(new_n940), .B2(new_n933), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n751), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1010), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(KEYINPUT123), .A3(G301), .A4(new_n1012), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT54), .B1(new_n1077), .B2(new_n1015), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1025), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1007), .B1(new_n992), .B2(new_n994), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n992), .A2(new_n994), .A3(new_n980), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n1083));
  INV_X1    g658(.A(new_n966), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1084), .A2(G1976), .A3(G288), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n965), .B1(new_n1085), .B2(new_n960), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT118), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1009), .A2(new_n1081), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n983), .A2(new_n934), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(new_n1048), .A3(new_n744), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1092), .A2(KEYINPUT109), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(KEYINPUT109), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n776), .B(new_n781), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1048), .B2(new_n744), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1093), .A2(new_n1094), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1091), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n704), .B(new_n707), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G290), .B(G1986), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1090), .A2(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n701), .A2(new_n1097), .A3(new_n703), .A4(new_n707), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n776), .A2(G2067), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1091), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1091), .A2(new_n1048), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT46), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(KEYINPUT124), .B2(KEYINPUT46), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1095), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1091), .B1(new_n743), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT47), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1098), .A2(G1986), .A3(G290), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT125), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT48), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1106), .B(new_n1116), .C1(new_n1100), .C2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT126), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1103), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g697(.A1(G227), .A2(G401), .A3(new_n462), .ZN(new_n1124));
  NOR3_X1   g698(.A1(new_n840), .A2(G229), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g699(.A1(new_n1125), .A2(new_n899), .ZN(G225));
  INV_X1    g700(.A(G225), .ZN(G308));
endmodule


