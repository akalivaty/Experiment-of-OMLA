

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XOR2_X1 U324 ( .A(G176GAT), .B(G64GAT), .Z(n416) );
  XNOR2_X2 U325 ( .A(n472), .B(n471), .ZN(n530) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n473) );
  NOR2_X2 U327 ( .A1(n547), .A2(n475), .ZN(n571) );
  XNOR2_X1 U328 ( .A(n324), .B(n344), .ZN(n325) );
  NOR2_X1 U329 ( .A1(n408), .A2(n407), .ZN(n531) );
  XNOR2_X1 U330 ( .A(n470), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U331 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U332 ( .A(n433), .B(n432), .ZN(n577) );
  XNOR2_X1 U333 ( .A(n477), .B(KEYINPUT121), .ZN(n478) );
  XNOR2_X1 U334 ( .A(n326), .B(n325), .ZN(n327) );
  NOR2_X2 U335 ( .A1(n533), .A2(n480), .ZN(n567) );
  XOR2_X2 U336 ( .A(n577), .B(n462), .Z(n562) );
  XNOR2_X1 U337 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n458) );
  XNOR2_X1 U338 ( .A(n459), .B(n458), .ZN(n461) );
  INV_X1 U339 ( .A(KEYINPUT22), .ZN(n366) );
  INV_X1 U340 ( .A(KEYINPUT102), .ZN(n412) );
  XNOR2_X1 U341 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U342 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U343 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U344 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U345 ( .A(n415), .B(n414), .ZN(n517) );
  XOR2_X1 U346 ( .A(n310), .B(n353), .Z(n522) );
  XNOR2_X1 U347 ( .A(KEYINPUT122), .B(G169GAT), .ZN(n481) );
  XNOR2_X1 U348 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U349 ( .A(n482), .B(n481), .ZN(G1348GAT) );
  XNOR2_X1 U350 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(G176GAT), .B(KEYINPUT87), .Z(n293) );
  XNOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT66), .ZN(n292) );
  XNOR2_X1 U353 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U354 ( .A(G190GAT), .B(G134GAT), .Z(n295) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U356 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U357 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U358 ( .A(G183GAT), .B(KEYINPUT86), .ZN(n296) );
  XNOR2_X1 U359 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U360 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U361 ( .A(G113GAT), .B(KEYINPUT0), .Z(n395) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G71GAT), .Z(n427) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G127GAT), .Z(n330) );
  XOR2_X1 U364 ( .A(n427), .B(n330), .Z(n301) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U366 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U367 ( .A(n395), .B(n302), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U370 ( .A(KEYINPUT18), .B(KEYINPUT85), .Z(n308) );
  XNOR2_X1 U371 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n307) );
  XNOR2_X1 U372 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(n309), .ZN(n353) );
  XOR2_X1 U374 ( .A(KEYINPUT75), .B(KEYINPUT78), .Z(n312) );
  XNOR2_X1 U375 ( .A(KEYINPUT76), .B(KEYINPUT9), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n328) );
  XOR2_X1 U377 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n314) );
  NAND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U380 ( .A(n315), .B(KEYINPUT11), .Z(n321) );
  XOR2_X1 U381 ( .A(G29GAT), .B(G43GAT), .Z(n317) );
  XNOR2_X1 U382 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n316) );
  XNOR2_X1 U383 ( .A(n317), .B(n316), .ZN(n437) );
  XOR2_X1 U384 ( .A(KEYINPUT72), .B(G85GAT), .Z(n319) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(G106GAT), .ZN(n318) );
  XNOR2_X1 U386 ( .A(n319), .B(n318), .ZN(n431) );
  XNOR2_X1 U387 ( .A(n437), .B(n431), .ZN(n320) );
  XOR2_X1 U388 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U389 ( .A(G50GAT), .B(G162GAT), .Z(n359) );
  XOR2_X1 U390 ( .A(G134GAT), .B(KEYINPUT77), .Z(n394) );
  XNOR2_X1 U391 ( .A(n359), .B(n394), .ZN(n324) );
  XOR2_X1 U392 ( .A(G92GAT), .B(G218GAT), .Z(n323) );
  XNOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U394 ( .A(n323), .B(n322), .ZN(n344) );
  XOR2_X1 U395 ( .A(n328), .B(n327), .Z(n557) );
  XNOR2_X1 U396 ( .A(n557), .B(KEYINPUT79), .ZN(n487) );
  XNOR2_X1 U397 ( .A(KEYINPUT36), .B(n487), .ZN(n585) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(G211GAT), .ZN(n329) );
  XOR2_X1 U399 ( .A(G8GAT), .B(G183GAT), .Z(n347) );
  XNOR2_X1 U400 ( .A(n329), .B(n347), .ZN(n343) );
  XOR2_X1 U401 ( .A(G57GAT), .B(KEYINPUT13), .Z(n424) );
  XOR2_X1 U402 ( .A(n424), .B(n330), .Z(n332) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U404 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U405 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n334) );
  XNOR2_X1 U406 ( .A(KEYINPUT15), .B(KEYINPUT80), .ZN(n333) );
  XNOR2_X1 U407 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U408 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G1GAT), .Z(n436) );
  XOR2_X1 U410 ( .A(KEYINPUT12), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U411 ( .A(G155GAT), .B(G78GAT), .ZN(n337) );
  XNOR2_X1 U412 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U413 ( .A(n436), .B(n339), .ZN(n340) );
  XNOR2_X1 U414 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U415 ( .A(n343), .B(n342), .Z(n581) );
  XOR2_X1 U416 ( .A(KEYINPUT98), .B(n344), .Z(n346) );
  NAND2_X1 U417 ( .A1(G226GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U418 ( .A(n346), .B(n345), .ZN(n348) );
  XOR2_X1 U419 ( .A(n348), .B(n347), .Z(n352) );
  XOR2_X1 U420 ( .A(G204GAT), .B(G211GAT), .Z(n350) );
  XNOR2_X1 U421 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n365), .B(n416), .ZN(n351) );
  XNOR2_X1 U424 ( .A(n352), .B(n351), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n354), .B(n353), .ZN(n519) );
  NAND2_X1 U426 ( .A1(n522), .A2(n519), .ZN(n355) );
  XNOR2_X1 U427 ( .A(KEYINPUT100), .B(n355), .ZN(n375) );
  XOR2_X1 U428 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n357) );
  XNOR2_X1 U429 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n356) );
  XNOR2_X1 U430 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U431 ( .A(G106GAT), .B(G218GAT), .Z(n358) );
  XNOR2_X1 U432 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U433 ( .A(G148GAT), .B(G78GAT), .Z(n417) );
  XNOR2_X1 U434 ( .A(n360), .B(n417), .ZN(n361) );
  XOR2_X1 U435 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U436 ( .A1(G228GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n365), .B(KEYINPUT23), .ZN(n367) );
  XOR2_X1 U439 ( .A(KEYINPUT2), .B(G155GAT), .Z(n371) );
  XNOR2_X1 U440 ( .A(G141GAT), .B(KEYINPUT90), .ZN(n370) );
  XNOR2_X1 U441 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U442 ( .A(KEYINPUT91), .B(KEYINPUT3), .Z(n372) );
  XOR2_X1 U443 ( .A(n373), .B(n372), .Z(n393) );
  XOR2_X1 U444 ( .A(n374), .B(n393), .Z(n476) );
  NAND2_X1 U445 ( .A1(n375), .A2(n476), .ZN(n376) );
  XOR2_X1 U446 ( .A(KEYINPUT25), .B(n376), .Z(n380) );
  NOR2_X1 U447 ( .A1(n476), .A2(n522), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n377), .B(KEYINPUT26), .ZN(n570) );
  XOR2_X1 U449 ( .A(n519), .B(KEYINPUT99), .Z(n378) );
  XOR2_X1 U450 ( .A(KEYINPUT27), .B(n378), .Z(n408) );
  INV_X1 U451 ( .A(n408), .ZN(n379) );
  NAND2_X1 U452 ( .A1(n570), .A2(n379), .ZN(n549) );
  NAND2_X1 U453 ( .A1(n380), .A2(n549), .ZN(n406) );
  XOR2_X1 U454 ( .A(G57GAT), .B(KEYINPUT97), .Z(n382) );
  XNOR2_X1 U455 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n381) );
  XNOR2_X1 U456 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U457 ( .A(G148GAT), .B(G162GAT), .Z(n384) );
  XNOR2_X1 U458 ( .A(G127GAT), .B(G120GAT), .ZN(n383) );
  XNOR2_X1 U459 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U460 ( .A(n386), .B(n385), .ZN(n405) );
  XOR2_X1 U461 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n388) );
  XNOR2_X1 U462 ( .A(KEYINPUT93), .B(KEYINPUT96), .ZN(n387) );
  XNOR2_X1 U463 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U464 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n390) );
  XNOR2_X1 U465 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n389) );
  XNOR2_X1 U466 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U467 ( .A(n392), .B(n391), .ZN(n403) );
  INV_X1 U468 ( .A(n393), .ZN(n399) );
  XOR2_X1 U469 ( .A(G85GAT), .B(n394), .Z(n397) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(n395), .ZN(n396) );
  XNOR2_X1 U471 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n399), .B(n398), .ZN(n401) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U474 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U475 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U476 ( .A(n405), .B(n404), .Z(n457) );
  NAND2_X1 U477 ( .A1(n406), .A2(n457), .ZN(n410) );
  XOR2_X1 U478 ( .A(n476), .B(KEYINPUT28), .Z(n525) );
  OR2_X1 U479 ( .A1(n457), .A2(n525), .ZN(n407) );
  INV_X1 U480 ( .A(n522), .ZN(n533) );
  NAND2_X1 U481 ( .A1(n531), .A2(n533), .ZN(n409) );
  NAND2_X1 U482 ( .A1(n410), .A2(n409), .ZN(n490) );
  NAND2_X1 U483 ( .A1(n581), .A2(n490), .ZN(n411) );
  NOR2_X1 U484 ( .A1(n585), .A2(n411), .ZN(n415) );
  XNOR2_X1 U485 ( .A(KEYINPUT37), .B(KEYINPUT101), .ZN(n413) );
  XOR2_X1 U486 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U489 ( .A(KEYINPUT71), .B(KEYINPUT73), .Z(n421) );
  XNOR2_X1 U490 ( .A(KEYINPUT70), .B(KEYINPUT32), .ZN(n420) );
  XNOR2_X1 U491 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U492 ( .A(n423), .B(n422), .Z(n429) );
  XNOR2_X1 U493 ( .A(G204GAT), .B(G92GAT), .ZN(n425) );
  XNOR2_X1 U494 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U497 ( .A(n430), .B(KEYINPUT33), .Z(n433) );
  XNOR2_X1 U498 ( .A(n431), .B(KEYINPUT31), .ZN(n432) );
  XOR2_X1 U499 ( .A(G197GAT), .B(G15GAT), .Z(n435) );
  XNOR2_X1 U500 ( .A(G169GAT), .B(G113GAT), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n450) );
  XOR2_X1 U502 ( .A(n436), .B(G36GAT), .Z(n439) );
  XNOR2_X1 U503 ( .A(n437), .B(G50GAT), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U505 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n441) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U507 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U508 ( .A(n443), .B(n442), .Z(n448) );
  XOR2_X1 U509 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n445) );
  XNOR2_X1 U510 ( .A(G141GAT), .B(G8GAT), .ZN(n444) );
  XNOR2_X1 U511 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U512 ( .A(n446), .B(KEYINPUT67), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U514 ( .A(n450), .B(n449), .ZN(n550) );
  NAND2_X1 U515 ( .A1(n577), .A2(n550), .ZN(n492) );
  NOR2_X1 U516 ( .A1(n517), .A2(n492), .ZN(n451) );
  XOR2_X1 U517 ( .A(KEYINPUT38), .B(n451), .Z(n452) );
  XNOR2_X1 U518 ( .A(KEYINPUT103), .B(n452), .ZN(n503) );
  NAND2_X1 U519 ( .A1(n522), .A2(n503), .ZN(n456) );
  XOR2_X1 U520 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n454) );
  XNOR2_X1 U521 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n453) );
  INV_X1 U522 ( .A(n457), .ZN(n547) );
  NOR2_X1 U523 ( .A1(n585), .A2(n581), .ZN(n459) );
  INV_X1 U524 ( .A(n550), .ZN(n572) );
  AND2_X1 U525 ( .A1(n577), .A2(n572), .ZN(n460) );
  NAND2_X1 U526 ( .A1(n461), .A2(n460), .ZN(n469) );
  INV_X1 U527 ( .A(n581), .ZN(n568) );
  XNOR2_X1 U528 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n462) );
  AND2_X1 U529 ( .A1(n550), .A2(n562), .ZN(n463) );
  XNOR2_X1 U530 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  NOR2_X1 U531 ( .A1(n568), .A2(n464), .ZN(n466) );
  INV_X1 U532 ( .A(n557), .ZN(n465) );
  NAND2_X1 U533 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U534 ( .A(n467), .B(KEYINPUT47), .Z(n468) );
  AND2_X1 U535 ( .A1(n469), .A2(n468), .ZN(n472) );
  INV_X1 U536 ( .A(KEYINPUT64), .ZN(n470) );
  NAND2_X1 U537 ( .A1(n530), .A2(n519), .ZN(n474) );
  AND2_X1 U538 ( .A1(n571), .A2(n476), .ZN(n479) );
  INV_X1 U539 ( .A(KEYINPUT55), .ZN(n477) );
  NAND2_X1 U540 ( .A1(n550), .A2(n567), .ZN(n482) );
  INV_X1 U541 ( .A(G190GAT), .ZN(n486) );
  INV_X1 U542 ( .A(n487), .ZN(n541) );
  NAND2_X1 U543 ( .A1(n567), .A2(n541), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1351GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n489) );
  NAND2_X1 U548 ( .A1(n568), .A2(n487), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n491), .A2(n490), .ZN(n505) );
  NOR2_X1 U551 ( .A1(n492), .A2(n505), .ZN(n498) );
  NAND2_X1 U552 ( .A1(n498), .A2(n547), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT34), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n519), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .Z(n497) );
  NAND2_X1 U558 ( .A1(n498), .A2(n522), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n525), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U562 ( .A1(n547), .A2(n503), .ZN(n501) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n519), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n503), .A2(n525), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n572), .A2(n562), .ZN(n516) );
  NOR2_X1 U571 ( .A1(n516), .A2(n505), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n547), .A2(n511), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n519), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n508), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n522), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U580 ( .A1(n511), .A2(n525), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(n515) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT108), .Z(n514) );
  XNOR2_X1 U583 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n547), .A2(n526), .ZN(n518) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  XOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT109), .Z(n521) );
  NAND2_X1 U588 ( .A1(n526), .A2(n519), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n522), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(KEYINPUT110), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n550), .A2(n542), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U602 ( .A1(n542), .A2(n562), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n539) );
  NAND2_X1 U606 ( .A1(n542), .A2(n568), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT116), .Z(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n547), .A2(n530), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n550), .A2(n558), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n553) );
  NAND2_X1 U619 ( .A1(n558), .A2(n562), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n568), .A2(n558), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n567), .A2(n562), .ZN(n564) );
  XOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT57), .Z(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n584) );
  NOR2_X1 U637 ( .A1(n584), .A2(n572), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n584), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

