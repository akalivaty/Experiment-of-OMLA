

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730;

  XNOR2_X1 U368 ( .A(n575), .B(KEYINPUT38), .ZN(n648) );
  BUF_X1 U369 ( .A(G107), .Z(n347) );
  XNOR2_X1 U370 ( .A(n501), .B(KEYINPUT16), .ZN(n410) );
  INV_X2 U371 ( .A(G953), .ZN(n711) );
  NAND2_X1 U372 ( .A1(n346), .A2(n454), .ZN(n420) );
  NAND2_X1 U373 ( .A1(n452), .A2(n453), .ZN(n346) );
  AND2_X4 U374 ( .A1(n371), .A2(n348), .ZN(n698) );
  NAND2_X2 U375 ( .A1(n609), .A2(n608), .ZN(n348) );
  XOR2_X1 U376 ( .A(n351), .B(n467), .Z(n349) );
  NOR2_X2 U377 ( .A1(G902), .A2(n691), .ZN(n490) );
  NOR2_X1 U378 ( .A1(n702), .A2(n718), .ZN(n682) );
  XNOR2_X2 U379 ( .A(n588), .B(KEYINPUT41), .ZN(n673) );
  NOR2_X2 U380 ( .A1(n524), .A2(n558), .ZN(n498) );
  XNOR2_X2 U381 ( .A(n462), .B(KEYINPUT0), .ZN(n361) );
  NAND2_X1 U382 ( .A1(n359), .A2(n430), .ZN(n718) );
  NOR2_X1 U383 ( .A1(n583), .A2(n559), .ZN(n563) );
  INV_X1 U384 ( .A(n634), .ZN(n378) );
  NOR2_X1 U385 ( .A1(n571), .A2(n529), .ZN(n530) );
  INV_X1 U386 ( .A(KEYINPUT76), .ZN(n429) );
  NAND2_X1 U387 ( .A1(n682), .A2(KEYINPUT2), .ZN(n371) );
  AND2_X1 U388 ( .A1(n364), .A2(n362), .ZN(n549) );
  XNOR2_X1 U389 ( .A(n718), .B(n429), .ZN(n358) );
  NOR2_X1 U390 ( .A1(n531), .A2(n547), .ZN(n391) );
  XNOR2_X1 U391 ( .A(n589), .B(KEYINPUT42), .ZN(n360) );
  OR2_X1 U392 ( .A1(n524), .A2(n582), .ZN(n669) );
  NOR2_X1 U393 ( .A1(n558), .A2(n377), .ZN(n376) );
  XNOR2_X1 U394 ( .A(n478), .B(n477), .ZN(n660) );
  NOR2_X1 U395 ( .A1(n554), .A2(n553), .ZN(n576) );
  OR2_X1 U396 ( .A1(n694), .A2(G902), .ZN(n408) );
  XOR2_X1 U397 ( .A(n607), .B(KEYINPUT65), .Z(n608) );
  INV_X1 U398 ( .A(n647), .ZN(n377) );
  XNOR2_X1 U399 ( .A(n451), .B(KEYINPUT71), .ZN(n413) );
  XOR2_X1 U400 ( .A(G146), .B(G125), .Z(n463) );
  XNOR2_X1 U401 ( .A(G119), .B(G113), .ZN(n412) );
  XNOR2_X1 U402 ( .A(n603), .B(KEYINPUT48), .ZN(n359) );
  XNOR2_X1 U403 ( .A(n535), .B(KEYINPUT103), .ZN(n587) );
  NAND2_X1 U404 ( .A1(n567), .A2(n571), .ZN(n535) );
  XOR2_X1 U405 ( .A(KEYINPUT66), .B(G101), .Z(n491) );
  XNOR2_X1 U406 ( .A(n439), .B(n503), .ZN(n717) );
  XNOR2_X1 U407 ( .A(n485), .B(n440), .ZN(n439) );
  XNOR2_X1 U408 ( .A(n441), .B(G137), .ZN(n440) );
  INV_X1 U409 ( .A(G131), .ZN(n441) );
  INV_X1 U410 ( .A(n582), .ZN(n664) );
  INV_X1 U411 ( .A(G469), .ZN(n489) );
  NOR2_X1 U412 ( .A1(n699), .A2(G902), .ZN(n478) );
  INV_X1 U413 ( .A(KEYINPUT25), .ZN(n475) );
  XNOR2_X1 U414 ( .A(n491), .B(n710), .ZN(n481) );
  XNOR2_X1 U415 ( .A(n717), .B(n486), .ZN(n495) );
  INV_X1 U416 ( .A(G146), .ZN(n486) );
  XNOR2_X1 U417 ( .A(n370), .B(KEYINPUT86), .ZN(n545) );
  NAND2_X1 U418 ( .A1(n728), .A2(n626), .ZN(n370) );
  NAND2_X1 U419 ( .A1(n533), .A2(n532), .ZN(n366) );
  NAND2_X1 U420 ( .A1(n392), .A2(n391), .ZN(n533) );
  XNOR2_X1 U421 ( .A(n384), .B(n447), .ZN(n450) );
  XNOR2_X1 U422 ( .A(n463), .B(KEYINPUT79), .ZN(n447) );
  XNOR2_X1 U423 ( .A(n425), .B(n446), .ZN(n384) );
  OR2_X1 U424 ( .A1(G237), .A2(G902), .ZN(n456) );
  XNOR2_X1 U425 ( .A(n389), .B(n388), .ZN(n583) );
  INV_X1 U426 ( .A(KEYINPUT68), .ZN(n388) );
  NOR2_X1 U427 ( .A1(n556), .A2(n557), .ZN(n389) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n512) );
  XNOR2_X1 U429 ( .A(KEYINPUT5), .B(G116), .ZN(n492) );
  INV_X1 U430 ( .A(n643), .ZN(n431) );
  INV_X1 U431 ( .A(KEYINPUT107), .ZN(n380) );
  AND2_X1 U432 ( .A1(n529), .A2(n519), .ZN(n520) );
  NOR2_X1 U433 ( .A1(n361), .A2(n427), .ZN(n426) );
  INV_X1 U434 ( .A(n660), .ZN(n557) );
  INV_X1 U435 ( .A(n565), .ZN(n397) );
  XNOR2_X1 U436 ( .A(n472), .B(n716), .ZN(n699) );
  INV_X1 U437 ( .A(KEYINPUT123), .ZN(n443) );
  XNOR2_X1 U438 ( .A(n481), .B(n393), .ZN(n483) );
  XNOR2_X1 U439 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n600) );
  INV_X1 U441 ( .A(KEYINPUT47), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n369), .B(n367), .ZN(n425) );
  XNOR2_X1 U443 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n369) );
  NOR2_X1 U444 ( .A1(n368), .A2(G953), .ZN(n367) );
  INV_X1 U445 ( .A(G224), .ZN(n368) );
  NOR2_X1 U446 ( .A1(n661), .A2(n576), .ZN(n555) );
  XNOR2_X1 U447 ( .A(n484), .B(G134), .ZN(n503) );
  XOR2_X1 U448 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n514) );
  XOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .Z(n606) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n457) );
  INV_X1 U451 ( .A(n576), .ZN(n433) );
  NAND2_X1 U452 ( .A1(n587), .A2(n428), .ZN(n427) );
  INV_X1 U453 ( .A(n661), .ZN(n428) );
  XNOR2_X1 U454 ( .A(n363), .B(KEYINPUT72), .ZN(n362) );
  INV_X1 U455 ( .A(n503), .ZN(n504) );
  XNOR2_X1 U456 ( .A(n482), .B(n394), .ZN(n393) );
  INV_X1 U457 ( .A(G140), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n450), .B(n449), .ZN(n419) );
  INV_X1 U459 ( .A(KEYINPUT30), .ZN(n436) );
  XNOR2_X1 U460 ( .A(n505), .B(n409), .ZN(n567) );
  XNOR2_X1 U461 ( .A(G478), .B(KEYINPUT100), .ZN(n409) );
  NOR2_X1 U462 ( .A1(G902), .A2(n696), .ZN(n505) );
  XNOR2_X1 U463 ( .A(n383), .B(KEYINPUT19), .ZN(n595) );
  XNOR2_X1 U464 ( .A(n584), .B(KEYINPUT28), .ZN(n586) );
  NOR2_X1 U465 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U466 ( .A(n518), .B(n407), .ZN(n406) );
  INV_X1 U467 ( .A(G475), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n437), .B(n495), .ZN(n617) );
  XNOR2_X1 U469 ( .A(n493), .B(n494), .ZN(n438) );
  NOR2_X1 U470 ( .A1(G953), .A2(n719), .ZN(n720) );
  OR2_X1 U471 ( .A1(G953), .A2(n702), .ZN(n707) );
  XNOR2_X1 U472 ( .A(n405), .B(n403), .ZN(n696) );
  XNOR2_X1 U473 ( .A(n404), .B(n501), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n375), .B(n504), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n500), .B(n350), .ZN(n404) );
  XNOR2_X1 U476 ( .A(n560), .B(n379), .ZN(n562) );
  XNOR2_X1 U477 ( .A(n561), .B(n380), .ZN(n379) );
  XNOR2_X1 U478 ( .A(n390), .B(KEYINPUT36), .ZN(n564) );
  XNOR2_X1 U479 ( .A(n445), .B(n415), .ZN(n414) );
  INV_X1 U480 ( .A(KEYINPUT82), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n525), .B(KEYINPUT31), .ZN(n526) );
  NOR2_X1 U482 ( .A1(n397), .A2(n557), .ZN(n396) );
  XNOR2_X1 U483 ( .A(n444), .B(n442), .ZN(n700) );
  XNOR2_X1 U484 ( .A(n699), .B(n443), .ZN(n442) );
  INV_X1 U485 ( .A(KEYINPUT60), .ZN(n399) );
  XNOR2_X1 U486 ( .A(n689), .B(n395), .ZN(n692) );
  INV_X1 U487 ( .A(KEYINPUT56), .ZN(n386) );
  XNOR2_X1 U488 ( .A(n688), .B(n385), .ZN(G75) );
  XNOR2_X1 U489 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n385) );
  NOR2_X1 U490 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U491 ( .A(n360), .B(n729), .ZN(G39) );
  XOR2_X1 U492 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n350) );
  XOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT77), .Z(n351) );
  AND2_X1 U494 ( .A1(G210), .A2(n456), .ZN(n352) );
  AND2_X1 U495 ( .A1(n582), .A2(n543), .ZN(n353) );
  AND2_X1 U496 ( .A1(G953), .A2(G902), .ZN(n354) );
  XOR2_X1 U497 ( .A(n694), .B(n693), .Z(n355) );
  XOR2_X1 U498 ( .A(n617), .B(KEYINPUT62), .Z(n356) );
  NOR2_X1 U499 ( .A1(G952), .A2(n711), .ZN(n701) );
  INV_X1 U500 ( .A(n701), .ZN(n422) );
  XNOR2_X2 U501 ( .A(n410), .B(n357), .ZN(n708) );
  XNOR2_X1 U502 ( .A(n438), .B(n357), .ZN(n437) );
  XNOR2_X2 U503 ( .A(n413), .B(n412), .ZN(n357) );
  NAND2_X1 U504 ( .A1(n358), .A2(n606), .ZN(n605) );
  NOR2_X2 U505 ( .A1(n360), .A2(n730), .ZN(n374) );
  NOR2_X1 U506 ( .A1(n361), .A2(n669), .ZN(n527) );
  XNOR2_X1 U507 ( .A(n361), .B(KEYINPUT90), .ZN(n522) );
  NAND2_X1 U508 ( .A1(n372), .A2(n373), .ZN(n363) );
  NOR2_X1 U509 ( .A1(n548), .A2(n365), .ZN(n364) );
  NAND2_X1 U510 ( .A1(n366), .A2(n618), .ZN(n365) );
  NAND2_X1 U511 ( .A1(n540), .A2(n557), .ZN(n618) );
  NAND2_X1 U512 ( .A1(n698), .A2(G475), .ZN(n402) );
  NAND2_X1 U513 ( .A1(n698), .A2(G472), .ZN(n424) );
  XNOR2_X1 U514 ( .A(n424), .B(n356), .ZN(n423) );
  XNOR2_X1 U515 ( .A(n402), .B(n355), .ZN(n401) );
  AND2_X1 U516 ( .A1(n727), .A2(n547), .ZN(n372) );
  NAND2_X1 U517 ( .A1(n401), .A2(n422), .ZN(n400) );
  NAND2_X1 U518 ( .A1(n423), .A2(n422), .ZN(n421) );
  NOR2_X1 U519 ( .A1(n727), .A2(KEYINPUT85), .ZN(n544) );
  XNOR2_X2 U520 ( .A(n416), .B(n414), .ZN(n727) );
  NOR2_X1 U521 ( .A1(n547), .A2(n546), .ZN(n548) );
  INV_X1 U522 ( .A(n545), .ZN(n373) );
  NAND2_X1 U523 ( .A1(n708), .A2(n481), .ZN(n454) );
  XNOR2_X2 U524 ( .A(n496), .B(n497), .ZN(n582) );
  INV_X1 U525 ( .A(n727), .ZN(n392) );
  XOR2_X2 U526 ( .A(KEYINPUT4), .B(KEYINPUT67), .Z(n485) );
  XNOR2_X1 U527 ( .A(n374), .B(KEYINPUT46), .ZN(n590) );
  NOR2_X1 U528 ( .A1(n645), .A2(n431), .ZN(n430) );
  INV_X1 U529 ( .A(n567), .ZN(n529) );
  NOR2_X2 U530 ( .A1(n652), .A2(n650), .ZN(n588) );
  NAND2_X1 U531 ( .A1(n502), .A2(G217), .ZN(n375) );
  NAND2_X1 U532 ( .A1(n378), .A2(n376), .ZN(n559) );
  NAND2_X1 U533 ( .A1(n631), .A2(n597), .ZN(n382) );
  XNOR2_X1 U534 ( .A(n349), .B(n468), .ZN(n471) );
  NAND2_X1 U535 ( .A1(n611), .A2(n473), .ZN(n418) );
  XNOR2_X2 U536 ( .A(n420), .B(n419), .ZN(n611) );
  NAND2_X1 U537 ( .A1(n566), .A2(n647), .ZN(n383) );
  XNOR2_X2 U538 ( .A(n549), .B(KEYINPUT45), .ZN(n702) );
  XNOR2_X1 U539 ( .A(n426), .B(n536), .ZN(n543) );
  XNOR2_X1 U540 ( .A(n387), .B(n386), .ZN(G51) );
  NAND2_X1 U541 ( .A1(n616), .A2(n422), .ZN(n387) );
  NAND2_X1 U542 ( .A1(n458), .A2(n354), .ZN(n550) );
  XNOR2_X1 U543 ( .A(n530), .B(KEYINPUT101), .ZN(n580) );
  NAND2_X1 U544 ( .A1(n563), .A2(n566), .ZN(n390) );
  XNOR2_X1 U545 ( .A(n691), .B(n690), .ZN(n395) );
  NAND2_X1 U546 ( .A1(n353), .A2(n396), .ZN(n626) );
  XNOR2_X2 U547 ( .A(n398), .B(KEYINPUT32), .ZN(n728) );
  NAND2_X1 U548 ( .A1(n543), .A2(n542), .ZN(n398) );
  XNOR2_X1 U549 ( .A(n400), .B(n399), .ZN(G60) );
  XNOR2_X2 U550 ( .A(n411), .B(G122), .ZN(n501) );
  XNOR2_X2 U551 ( .A(n408), .B(n406), .ZN(n571) );
  XNOR2_X2 U552 ( .A(G116), .B(G107), .ZN(n411) );
  NAND2_X1 U553 ( .A1(n521), .A2(n520), .ZN(n416) );
  AND2_X1 U554 ( .A1(n417), .A2(n592), .ZN(n531) );
  NAND2_X1 U555 ( .A1(n637), .A2(n620), .ZN(n417) );
  XNOR2_X2 U556 ( .A(n418), .B(n352), .ZN(n566) );
  XNOR2_X1 U557 ( .A(n421), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U558 ( .A(n527), .B(n526), .ZN(n637) );
  NAND2_X1 U559 ( .A1(n434), .A2(n432), .ZN(n579) );
  AND2_X1 U560 ( .A1(n648), .A2(n433), .ZN(n432) );
  INV_X1 U561 ( .A(n577), .ZN(n434) );
  NAND2_X1 U562 ( .A1(n435), .A2(n570), .ZN(n577) );
  XNOR2_X1 U563 ( .A(n569), .B(n436), .ZN(n435) );
  NAND2_X1 U564 ( .A1(n698), .A2(G217), .ZN(n444) );
  XNOR2_X1 U565 ( .A(n615), .B(n614), .ZN(n616) );
  OR2_X2 U566 ( .A1(n702), .A2(n605), .ZN(n609) );
  XNOR2_X1 U567 ( .A(n579), .B(n578), .ZN(n604) );
  INV_X1 U568 ( .A(n571), .ZN(n519) );
  XNOR2_X1 U569 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n445) );
  INV_X1 U570 ( .A(KEYINPUT93), .ZN(n525) );
  XNOR2_X1 U571 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U572 ( .A(KEYINPUT73), .B(KEYINPUT39), .ZN(n578) );
  XOR2_X1 U573 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n446) );
  XNOR2_X2 U574 ( .A(G143), .B(G128), .ZN(n484) );
  INV_X1 U575 ( .A(n484), .ZN(n448) );
  XOR2_X1 U576 ( .A(n448), .B(n485), .Z(n449) );
  XNOR2_X1 U577 ( .A(G110), .B(G104), .ZN(n710) );
  INV_X1 U578 ( .A(n481), .ZN(n453) );
  XNOR2_X2 U579 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n451) );
  INV_X1 U580 ( .A(n708), .ZN(n452) );
  INV_X1 U581 ( .A(n606), .ZN(n473) );
  NAND2_X1 U582 ( .A1(G214), .A2(n456), .ZN(n647) );
  XNOR2_X1 U583 ( .A(n457), .B(KEYINPUT14), .ZN(n458) );
  NAND2_X1 U584 ( .A1(G952), .A2(n458), .ZN(n680) );
  NOR2_X1 U585 ( .A1(G953), .A2(n680), .ZN(n554) );
  NOR2_X1 U586 ( .A1(G898), .A2(n550), .ZN(n459) );
  NOR2_X1 U587 ( .A1(n554), .A2(n459), .ZN(n460) );
  XNOR2_X1 U588 ( .A(KEYINPUT89), .B(n460), .ZN(n461) );
  NAND2_X1 U589 ( .A1(n595), .A2(n461), .ZN(n462) );
  XNOR2_X1 U590 ( .A(n463), .B(G140), .ZN(n464) );
  XNOR2_X1 U591 ( .A(n464), .B(KEYINPUT10), .ZN(n716) );
  XOR2_X1 U592 ( .A(G110), .B(G119), .Z(n466) );
  XNOR2_X1 U593 ( .A(G128), .B(G137), .ZN(n465) );
  XNOR2_X1 U594 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U595 ( .A(KEYINPUT23), .B(KEYINPUT91), .ZN(n467) );
  NAND2_X1 U596 ( .A1(G234), .A2(n711), .ZN(n469) );
  XOR2_X1 U597 ( .A(KEYINPUT8), .B(n469), .Z(n502) );
  NAND2_X1 U598 ( .A1(G221), .A2(n502), .ZN(n470) );
  XNOR2_X1 U599 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U600 ( .A1(n473), .A2(G234), .ZN(n474) );
  XNOR2_X1 U601 ( .A(n474), .B(KEYINPUT20), .ZN(n479) );
  NAND2_X1 U602 ( .A1(n479), .A2(G217), .ZN(n476) );
  NAND2_X1 U603 ( .A1(G221), .A2(n479), .ZN(n480) );
  XNOR2_X1 U604 ( .A(KEYINPUT21), .B(n480), .ZN(n661) );
  NOR2_X1 U605 ( .A1(n660), .A2(n661), .ZN(n658) );
  NAND2_X1 U606 ( .A1(G227), .A2(n711), .ZN(n482) );
  XOR2_X1 U607 ( .A(n483), .B(KEYINPUT78), .Z(n488) );
  XNOR2_X1 U608 ( .A(n495), .B(n347), .ZN(n487) );
  XNOR2_X1 U609 ( .A(n488), .B(n487), .ZN(n691) );
  XNOR2_X2 U610 ( .A(n490), .B(n489), .ZN(n585) );
  XNOR2_X2 U611 ( .A(n585), .B(KEYINPUT1), .ZN(n657) );
  NAND2_X1 U612 ( .A1(n658), .A2(n657), .ZN(n524) );
  XNOR2_X1 U613 ( .A(G472), .B(KEYINPUT92), .ZN(n497) );
  XNOR2_X1 U614 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U615 ( .A1(n512), .A2(G210), .ZN(n494) );
  NOR2_X1 U616 ( .A1(n617), .A2(G902), .ZN(n496) );
  XNOR2_X1 U617 ( .A(n664), .B(KEYINPUT6), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n498), .B(KEYINPUT33), .ZN(n646) );
  NOR2_X1 U619 ( .A1(n522), .A2(n646), .ZN(n499) );
  XNOR2_X1 U620 ( .A(n499), .B(KEYINPUT34), .ZN(n521) );
  XOR2_X1 U621 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n500) );
  XOR2_X1 U622 ( .A(G104), .B(G113), .Z(n507) );
  XNOR2_X1 U623 ( .A(G131), .B(G143), .ZN(n506) );
  XNOR2_X1 U624 ( .A(n507), .B(n506), .ZN(n511) );
  XOR2_X1 U625 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n509) );
  XNOR2_X1 U626 ( .A(G122), .B(KEYINPUT12), .ZN(n508) );
  XNOR2_X1 U627 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U628 ( .A(n511), .B(n510), .ZN(n516) );
  NAND2_X1 U629 ( .A1(G214), .A2(n512), .ZN(n513) );
  XNOR2_X1 U630 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U631 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U632 ( .A(n716), .B(n517), .ZN(n694) );
  XNOR2_X1 U633 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n518) );
  INV_X1 U634 ( .A(KEYINPUT44), .ZN(n547) );
  NAND2_X1 U635 ( .A1(n585), .A2(n658), .ZN(n568) );
  NOR2_X1 U636 ( .A1(n568), .A2(n522), .ZN(n523) );
  NAND2_X1 U637 ( .A1(n582), .A2(n523), .ZN(n620) );
  NAND2_X1 U638 ( .A1(n571), .A2(n529), .ZN(n528) );
  XNOR2_X1 U639 ( .A(n528), .B(KEYINPUT102), .ZN(n638) );
  NAND2_X1 U640 ( .A1(n638), .A2(n580), .ZN(n592) );
  OR2_X1 U641 ( .A1(n531), .A2(KEYINPUT85), .ZN(n532) );
  XNOR2_X1 U642 ( .A(KEYINPUT22), .B(KEYINPUT74), .ZN(n534) );
  XNOR2_X1 U643 ( .A(n534), .B(KEYINPUT64), .ZN(n536) );
  AND2_X1 U644 ( .A1(n543), .A2(n558), .ZN(n537) );
  XNOR2_X1 U645 ( .A(KEYINPUT83), .B(n537), .ZN(n538) );
  NOR2_X1 U646 ( .A1(n397), .A2(n538), .ZN(n539) );
  XNOR2_X1 U647 ( .A(n539), .B(KEYINPUT84), .ZN(n540) );
  INV_X1 U648 ( .A(n657), .ZN(n565) );
  NOR2_X1 U649 ( .A1(n557), .A2(n565), .ZN(n541) );
  AND2_X1 U650 ( .A1(n558), .A2(n541), .ZN(n542) );
  NOR2_X1 U651 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U652 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n561) );
  XOR2_X1 U653 ( .A(n550), .B(KEYINPUT105), .Z(n551) );
  NOR2_X1 U654 ( .A1(G900), .A2(n551), .ZN(n552) );
  XNOR2_X1 U655 ( .A(n552), .B(KEYINPUT106), .ZN(n553) );
  XNOR2_X1 U656 ( .A(n555), .B(KEYINPUT69), .ZN(n556) );
  XNOR2_X1 U657 ( .A(KEYINPUT104), .B(n580), .ZN(n634) );
  NAND2_X1 U658 ( .A1(n563), .A2(n565), .ZN(n560) );
  NOR2_X1 U659 ( .A1(n566), .A2(n562), .ZN(n645) );
  NOR2_X1 U660 ( .A1(n565), .A2(n564), .ZN(n640) );
  INV_X1 U661 ( .A(n566), .ZN(n575) );
  NOR2_X1 U662 ( .A1(n576), .A2(n567), .ZN(n573) );
  INV_X1 U663 ( .A(n568), .ZN(n570) );
  NAND2_X1 U664 ( .A1(n647), .A2(n664), .ZN(n569) );
  NOR2_X1 U665 ( .A1(n571), .A2(n577), .ZN(n572) );
  NAND2_X1 U666 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U667 ( .A1(n575), .A2(n574), .ZN(n630) );
  NOR2_X1 U668 ( .A1(n640), .A2(n630), .ZN(n591) );
  NOR2_X1 U669 ( .A1(n604), .A2(n580), .ZN(n581) );
  XNOR2_X1 U670 ( .A(n581), .B(KEYINPUT40), .ZN(n730) );
  NAND2_X1 U671 ( .A1(n586), .A2(n585), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n648), .A2(n647), .ZN(n652) );
  INV_X1 U673 ( .A(n587), .ZN(n650) );
  NOR2_X1 U674 ( .A1(n593), .A2(n673), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n591), .A2(n590), .ZN(n602) );
  INV_X1 U676 ( .A(n592), .ZN(n653) );
  NOR2_X1 U677 ( .A1(n653), .A2(KEYINPUT75), .ZN(n597) );
  INV_X1 U678 ( .A(n593), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X2 U680 ( .A(n596), .B(KEYINPUT81), .ZN(n631) );
  AND2_X1 U681 ( .A1(n653), .A2(KEYINPUT75), .ZN(n598) );
  NAND2_X1 U682 ( .A1(n598), .A2(n631), .ZN(n599) );
  NAND2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X2 U684 ( .A1(n602), .A2(n601), .ZN(n603) );
  OR2_X1 U685 ( .A1(n604), .A2(n638), .ZN(n643) );
  NAND2_X1 U686 ( .A1(KEYINPUT2), .A2(n606), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n698), .A2(G210), .ZN(n615) );
  XOR2_X1 U688 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n613) );
  XNOR2_X1 U689 ( .A(n611), .B(KEYINPUT55), .ZN(n612) );
  XNOR2_X1 U690 ( .A(G101), .B(n618), .ZN(G3) );
  NOR2_X1 U691 ( .A1(n634), .A2(n620), .ZN(n619) );
  XOR2_X1 U692 ( .A(G104), .B(n619), .Z(G6) );
  NOR2_X1 U693 ( .A1(n638), .A2(n620), .ZN(n625) );
  XOR2_X1 U694 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n622) );
  XNOR2_X1 U695 ( .A(n347), .B(KEYINPUT26), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U697 ( .A(KEYINPUT27), .B(n623), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n625), .B(n624), .ZN(G9) );
  XNOR2_X1 U699 ( .A(G110), .B(n626), .ZN(G12) );
  XOR2_X1 U700 ( .A(G128), .B(KEYINPUT29), .Z(n629) );
  INV_X1 U701 ( .A(n638), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n631), .A2(n627), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(G30) );
  XOR2_X1 U704 ( .A(G143), .B(n630), .Z(G45) );
  XOR2_X1 U705 ( .A(G146), .B(KEYINPUT111), .Z(n633) );
  NAND2_X1 U706 ( .A1(n631), .A2(n378), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n633), .B(n632), .ZN(G48) );
  NOR2_X1 U708 ( .A1(n634), .A2(n637), .ZN(n635) );
  XOR2_X1 U709 ( .A(KEYINPUT112), .B(n635), .Z(n636) );
  XNOR2_X1 U710 ( .A(G113), .B(n636), .ZN(G15) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U712 ( .A(G116), .B(n639), .Z(G18) );
  XOR2_X1 U713 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n642) );
  XNOR2_X1 U714 ( .A(G125), .B(n640), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(G27) );
  XNOR2_X1 U716 ( .A(G134), .B(KEYINPUT114), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(G36) );
  XOR2_X1 U718 ( .A(G140), .B(n645), .Z(G42) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT119), .B(n651), .Z(n655) );
  NOR2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n646), .A2(n656), .ZN(n677) );
  XOR2_X1 U725 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n672) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT50), .B(n659), .Z(n668) );
  XOR2_X1 U728 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n663) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U732 ( .A(KEYINPUT116), .B(n666), .ZN(n667) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U735 ( .A(n672), .B(n671), .ZN(n674) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U737 ( .A(n675), .B(KEYINPUT118), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U739 ( .A(n678), .B(KEYINPUT52), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U741 ( .A(KEYINPUT120), .B(n681), .Z(n684) );
  XNOR2_X1 U742 ( .A(KEYINPUT2), .B(n682), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n673), .A2(n646), .ZN(n685) );
  NAND2_X1 U745 ( .A1(n711), .A2(n687), .ZN(n688) );
  XOR2_X1 U746 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n690) );
  NAND2_X1 U747 ( .A1(n698), .A2(G469), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n701), .A2(n692), .ZN(G54) );
  INV_X1 U749 ( .A(KEYINPUT59), .ZN(n693) );
  NAND2_X1 U750 ( .A1(G478), .A2(n698), .ZN(n695) );
  XNOR2_X1 U751 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U752 ( .A1(n701), .A2(n697), .ZN(G63) );
  NOR2_X1 U753 ( .A1(n701), .A2(n700), .ZN(G66) );
  NAND2_X1 U754 ( .A1(G224), .A2(G953), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n703), .B(KEYINPUT124), .ZN(n704) );
  XNOR2_X1 U756 ( .A(KEYINPUT61), .B(n704), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n705), .A2(G898), .ZN(n706) );
  NAND2_X1 U758 ( .A1(n707), .A2(n706), .ZN(n715) );
  XOR2_X1 U759 ( .A(n708), .B(G101), .Z(n709) );
  XNOR2_X1 U760 ( .A(n710), .B(n709), .ZN(n713) );
  NOR2_X1 U761 ( .A1(G898), .A2(n711), .ZN(n712) );
  NOR2_X1 U762 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n715), .B(n714), .ZN(G69) );
  XOR2_X1 U764 ( .A(n717), .B(n716), .Z(n721) );
  XOR2_X1 U765 ( .A(n721), .B(n718), .Z(n719) );
  XNOR2_X1 U766 ( .A(n720), .B(KEYINPUT125), .ZN(n726) );
  XNOR2_X1 U767 ( .A(n721), .B(G227), .ZN(n722) );
  XNOR2_X1 U768 ( .A(n722), .B(KEYINPUT126), .ZN(n723) );
  NAND2_X1 U769 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U770 ( .A1(G953), .A2(n724), .ZN(n725) );
  NAND2_X1 U771 ( .A1(n726), .A2(n725), .ZN(G72) );
  XNOR2_X1 U772 ( .A(G122), .B(n727), .ZN(G24) );
  XNOR2_X1 U773 ( .A(n728), .B(G119), .ZN(G21) );
  XNOR2_X1 U774 ( .A(G137), .B(KEYINPUT127), .ZN(n729) );
  XOR2_X1 U775 ( .A(G131), .B(n730), .Z(G33) );
endmodule

