//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT65), .B(G244), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G77), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n215), .B(new_n216), .C1(new_n202), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT66), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n210), .B(new_n213), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n220), .B1(new_n219), .B2(new_n218), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n209), .B(new_n228), .C1(new_n222), .C2(new_n212), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n229), .A2(KEYINPUT0), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n233), .A2(G20), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n229), .A2(KEYINPUT0), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n230), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT64), .Z(new_n239));
  NOR2_X1   g0039(.A1(new_n226), .A2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G250), .B(G257), .Z(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G87), .B(G97), .Z(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  NAND2_X1  g0057(.A1(G33), .A2(G283), .ZN(new_n258));
  INV_X1    g0058(.A(G20), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n258), .B(new_n259), .C1(G33), .C2(new_n221), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n234), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n260), .B(new_n262), .C1(new_n259), .C2(G116), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT20), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT79), .ZN(new_n268));
  INV_X1    g0068(.A(new_n262), .ZN(new_n269));
  INV_X1    g0069(.A(G13), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n270), .A2(new_n259), .A3(G1), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n271), .A2(new_n262), .A3(KEYINPUT79), .ZN(new_n274));
  OAI211_X1 g0074(.A(G116), .B(new_n267), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G116), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n265), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n212), .A2(G1698), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(new_n284), .C1(G257), .C2(G1698), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT70), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n281), .A2(new_n289), .A3(new_n282), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G303), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n235), .B1(new_n280), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT5), .A2(G41), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT5), .A2(G41), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n266), .B(G45), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n300), .A2(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G270), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n297), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n278), .A2(new_n305), .A3(G169), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT21), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n305), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G179), .A3(new_n278), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n278), .A2(new_n305), .A3(KEYINPUT21), .A4(G169), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n305), .A2(G200), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n305), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n312), .B1(new_n278), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n291), .A2(new_n259), .A3(G87), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT22), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n259), .A2(G33), .A3(G116), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n211), .A2(G20), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT23), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n283), .A2(KEYINPUT22), .A3(new_n259), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n324), .A2(new_n208), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n319), .A2(new_n320), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT93), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT24), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n323), .B1(new_n324), .B2(new_n208), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n318), .B2(new_n317), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n328), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n331), .A2(new_n320), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n262), .A3(new_n334), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n262), .B(KEYINPUT71), .Z(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(new_n267), .A3(new_n272), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G107), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n321), .A2(G1), .A3(new_n270), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT25), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n222), .A2(G1698), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n283), .B(new_n343), .C1(G250), .C2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G294), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n280), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n295), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G264), .B2(new_n303), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n302), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n314), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(G200), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n342), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n350), .A2(G179), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n342), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(KEYINPUT94), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT94), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n342), .B2(new_n358), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n355), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT95), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT95), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n355), .B(new_n365), .C1(new_n360), .C2(new_n362), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n316), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n203), .A2(G20), .ZN(new_n368));
  INV_X1    g0168(.A(G150), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G20), .A2(G33), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT72), .B(KEYINPUT8), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G58), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n206), .A2(KEYINPUT8), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT73), .B1(new_n373), .B2(G58), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT74), .B1(new_n280), .B2(G20), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(new_n259), .A3(G33), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n368), .B1(new_n369), .B2(new_n371), .C1(new_n378), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n262), .B(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n271), .A2(new_n202), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n384), .A2(new_n271), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n266), .A2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(G50), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT9), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n291), .ZN(new_n395));
  INV_X1    g0195(.A(G1698), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(G222), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G223), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n396), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n296), .C1(G77), .C2(new_n291), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n301), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT69), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n404), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n405), .A2(new_n295), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G226), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n400), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G200), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n387), .A2(KEYINPUT9), .A3(new_n388), .A4(new_n391), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n409), .A2(new_n314), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n394), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT10), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n273), .A2(new_n274), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n266), .B2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G68), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n270), .A2(G1), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n259), .A2(G68), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT12), .ZN(new_n421));
  INV_X1    g0221(.A(G77), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n382), .A2(new_n422), .B1(new_n202), .B2(new_n371), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n384), .B1(new_n423), .B2(new_n419), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n417), .A2(new_n421), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n217), .A2(new_n396), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n291), .B(new_n429), .C1(G232), .C2(new_n396), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G97), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n296), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n407), .A2(G238), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(new_n403), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n402), .B1(new_n432), .B2(new_n296), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT13), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n434), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT14), .B1(new_n441), .B2(new_n357), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(G179), .A3(new_n439), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n444), .A3(G169), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT82), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n436), .A2(G190), .A3(new_n439), .ZN(new_n448));
  INV_X1    g0248(.A(new_n428), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G200), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n436), .B2(new_n439), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n447), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n452), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT82), .A3(new_n448), .A4(new_n449), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n428), .A2(new_n446), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n409), .A2(new_n357), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n392), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT76), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n409), .A2(G179), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT76), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n392), .A2(new_n461), .A3(new_n457), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT77), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n459), .A2(KEYINPUT77), .A3(new_n460), .A4(new_n462), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n414), .A2(new_n456), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT85), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT18), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n283), .B1(G223), .B2(G1698), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n396), .A2(G226), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n472), .A2(new_n473), .B1(new_n280), .B2(new_n208), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n296), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n407), .A2(G232), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n403), .ZN(new_n477));
  INV_X1    g0277(.A(G179), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(G169), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(KEYINPUT84), .A3(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n378), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n389), .A3(new_n390), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n378), .A2(new_n271), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G68), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n206), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(G20), .B1(new_n491), .B2(new_n201), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n370), .A2(G159), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT7), .ZN(new_n496));
  NOR4_X1   g0296(.A1(new_n286), .A2(new_n287), .A3(new_n496), .A4(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n288), .A2(new_n290), .A3(new_n259), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n495), .B1(new_n499), .B2(new_n490), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT16), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n496), .B1(new_n283), .B2(G20), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n286), .A2(new_n287), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(KEYINPUT7), .A3(new_n259), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n494), .B1(new_n506), .B2(G68), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n269), .B1(new_n507), .B2(KEYINPUT16), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT83), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n502), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n489), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n468), .B(new_n471), .C1(new_n485), .C2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n479), .A2(KEYINPUT84), .A3(new_n480), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT84), .B1(new_n479), .B2(new_n480), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n489), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n502), .A2(new_n511), .A3(new_n508), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n511), .B1(new_n502), .B2(new_n508), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n517), .A2(new_n469), .A3(new_n521), .A4(new_n470), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n477), .A2(new_n451), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G190), .B2(new_n477), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n525), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT17), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n510), .A2(new_n512), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(KEYINPUT17), .A3(new_n518), .A4(new_n525), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT86), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n528), .B2(new_n530), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n523), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G238), .A2(G1698), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n291), .B(new_n535), .C1(new_n207), .C2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(new_n296), .C1(G107), .C2(new_n291), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n407), .A2(new_n214), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n403), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G179), .ZN(new_n540));
  XOR2_X1   g0340(.A(new_n540), .B(KEYINPUT80), .Z(new_n541));
  NAND2_X1  g0341(.A1(new_n416), .A2(G77), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n271), .A2(new_n422), .ZN(new_n543));
  INV_X1    g0343(.A(new_n375), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n206), .A2(KEYINPUT8), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n370), .A2(KEYINPUT78), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n370), .A2(KEYINPUT78), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g0349(.A(KEYINPUT15), .B(G87), .ZN(new_n550));
  OAI221_X1 g0350(.A(new_n549), .B1(new_n259), .B2(new_n422), .C1(new_n382), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n262), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n542), .A2(new_n543), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(new_n357), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n555), .A2(KEYINPUT81), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(KEYINPUT81), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n541), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n553), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n539), .A2(G200), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n314), .C2(new_n539), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n534), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n467), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n283), .A2(new_n564), .A3(G244), .A4(new_n396), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G244), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n396), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n291), .B(new_n568), .C1(G250), .C2(new_n396), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n569), .B2(KEYINPUT4), .ZN(new_n570));
  INV_X1    g0370(.A(new_n258), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n296), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n303), .A2(G257), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n302), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT88), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n572), .A2(KEYINPUT88), .A3(new_n302), .A4(new_n573), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(G200), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n337), .A2(new_n221), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n370), .A2(G77), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT6), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n581), .A2(new_n221), .A3(G107), .ZN(new_n582));
  XNOR2_X1  g0382(.A(G97), .B(G107), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI221_X1 g0384(.A(new_n580), .B1(new_n259), .B2(new_n584), .C1(new_n499), .C2(new_n211), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n579), .B1(new_n585), .B2(new_n262), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n271), .A2(new_n221), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT87), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n574), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G190), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n578), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n574), .A2(new_n357), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n572), .A2(new_n478), .A3(new_n302), .A4(new_n573), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n590), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT89), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT92), .ZN(new_n601));
  INV_X1    g0401(.A(new_n550), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n272), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n379), .A2(new_n381), .A3(G97), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n259), .B1(new_n431), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n208), .A2(new_n221), .A3(new_n211), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n283), .A2(new_n259), .A3(G68), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n269), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n603), .B(new_n610), .C1(new_n338), .C2(G87), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G116), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n283), .A2(G244), .A3(G1698), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n283), .A2(G238), .A3(new_n396), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT91), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n612), .B(new_n613), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n296), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n266), .A2(G45), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(new_n301), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n295), .A2(G250), .A3(new_n620), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n623), .B(KEYINPUT90), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n619), .A2(G190), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n621), .B(new_n624), .C1(new_n618), .C2(new_n296), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n611), .B(new_n626), .C1(new_n627), .C2(new_n451), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n619), .A2(new_n478), .A3(new_n622), .A4(new_n625), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n610), .A2(new_n603), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n337), .B2(new_n550), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n629), .B(new_n631), .C1(new_n627), .C2(G169), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n597), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n600), .A2(new_n601), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n600), .A2(new_n634), .A3(new_n635), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT92), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n367), .A2(new_n563), .A3(new_n636), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(KEYINPUT96), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n628), .A2(new_n632), .A3(KEYINPUT96), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n641), .A2(new_n594), .A3(new_n597), .A4(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT97), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n312), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT97), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n645), .A2(new_n647), .B1(new_n342), .B2(new_n358), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n643), .A2(new_n648), .A3(new_n354), .ZN(new_n649));
  INV_X1    g0449(.A(new_n632), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n590), .A2(new_n596), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(new_n632), .A3(new_n628), .A4(new_n595), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(KEYINPUT98), .A3(new_n595), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT98), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n597), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n641), .A2(new_n654), .A3(new_n642), .A4(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n563), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n465), .A2(new_n466), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n446), .A2(new_n428), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n453), .A2(new_n455), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n558), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n532), .A2(new_n533), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n521), .A2(KEYINPUT18), .A3(new_n481), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT18), .B1(new_n521), .B2(new_n481), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n660), .B1(new_n672), .B2(new_n414), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n659), .A2(new_n673), .ZN(G369));
  NAND2_X1  g0474(.A1(new_n364), .A2(new_n366), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n270), .A2(G20), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n418), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT100), .Z(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n342), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n683), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n359), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n683), .A2(new_n278), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n645), .A2(new_n647), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n316), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n312), .A2(new_n683), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n675), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n359), .A2(new_n683), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(G399));
  NOR2_X1   g0500(.A1(new_n228), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n607), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n232), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(new_n658), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n643), .A2(new_n648), .A3(new_n354), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n683), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n312), .B1(new_n360), .B2(new_n362), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n641), .A2(new_n642), .ZN(new_n714));
  INV_X1    g0514(.A(new_n598), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n355), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n650), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(new_n686), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n710), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n367), .A2(new_n638), .A3(new_n636), .A4(new_n686), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n627), .A2(G179), .A3(new_n309), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n572), .A2(new_n302), .A3(new_n349), .A4(new_n573), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n350), .A2(new_n478), .A3(new_n305), .ZN(new_n728));
  OR3_X1    g0528(.A1(new_n592), .A2(new_n627), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(new_n683), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n722), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n712), .B(new_n721), .C1(G330), .C2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n706), .B1(new_n735), .B2(G1), .ZN(G364));
  OR2_X1    g0536(.A1(new_n690), .A2(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n676), .A2(G45), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n702), .A2(G1), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n737), .A2(new_n691), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT101), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n228), .A2(new_n283), .ZN(new_n742));
  INV_X1    g0542(.A(G45), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n233), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n742), .B(new_n744), .C1(new_n253), .C2(new_n743), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n291), .A2(new_n227), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n745), .B1(G116), .B2(new_n227), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT102), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n234), .B1(G20), .B2(new_n357), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n739), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n752), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n259), .A2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n451), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G283), .A2(new_n760), .B1(new_n763), .B2(G329), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n478), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n757), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n259), .B1(new_n761), .B2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n291), .B(new_n768), .C1(G294), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n259), .A2(new_n314), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n766), .ZN(new_n773));
  INV_X1    g0573(.A(G322), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n478), .A2(new_n451), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n757), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n772), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n775), .B(new_n781), .C1(G326), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(new_n758), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n771), .B(new_n784), .C1(new_n292), .C2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT103), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n769), .A2(new_n221), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n291), .B1(new_n211), .B2(new_n759), .ZN(new_n789));
  INV_X1    g0589(.A(new_n773), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n788), .B(new_n789), .C1(G58), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n785), .A2(new_n208), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n782), .A2(new_n202), .B1(new_n767), .B2(new_n422), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT32), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n762), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n763), .A2(KEYINPUT32), .A3(G159), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n792), .B(new_n793), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n791), .B(new_n798), .C1(new_n490), .C2(new_n777), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n787), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n753), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n755), .B1(new_n690), .B2(new_n756), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n741), .A2(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n734), .A2(G330), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n558), .A2(new_n561), .B1(new_n553), .B2(new_n683), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n553), .A2(new_n683), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n555), .B(KEYINPUT81), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n807), .B2(new_n541), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n686), .C1(new_n649), .C2(new_n658), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT104), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n804), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n709), .A2(new_n809), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n813), .A2(new_n815), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n816), .A2(new_n739), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n739), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n785), .A2(new_n202), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n759), .A2(new_n490), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n769), .A2(new_n206), .ZN(new_n822));
  OR4_X1    g0622(.A1(new_n504), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n777), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G143), .A2(new_n790), .B1(new_n824), .B2(G150), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n783), .A2(G137), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(new_n795), .C2(new_n767), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n828), .B2(new_n827), .C1(new_n830), .C2(new_n762), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n759), .A2(new_n208), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n211), .A2(new_n785), .B1(new_n773), .B2(new_n345), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G311), .B2(new_n763), .ZN(new_n834));
  INV_X1    g0634(.A(G283), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n782), .A2(new_n292), .B1(new_n777), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n767), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(G116), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n291), .A2(new_n788), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n831), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n753), .A2(new_n750), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n841), .A2(new_n753), .B1(new_n422), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n819), .B(new_n843), .C1(new_n809), .C2(new_n751), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n818), .A2(new_n844), .ZN(G384));
  INV_X1    g0645(.A(KEYINPUT40), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n733), .B(KEYINPUT110), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n722), .A2(new_n732), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n428), .A2(new_n683), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n456), .B(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n850), .A2(new_n809), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n507), .A2(KEYINPUT16), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n507), .A2(KEYINPUT16), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n384), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n518), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n681), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n514), .A2(new_n522), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n666), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n857), .B1(new_n481), .B2(new_n858), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(new_n526), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n521), .A2(new_n858), .ZN(new_n866));
  XOR2_X1   g0666(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n526), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n517), .A2(new_n521), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n853), .B1(new_n861), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n864), .B2(new_n863), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(KEYINPUT38), .C1(new_n534), .C2(new_n859), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n846), .B1(new_n852), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT108), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n528), .B(new_n530), .C1(new_n668), .C2(new_n669), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT107), .ZN(new_n881));
  INV_X1    g0681(.A(new_n866), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n521), .A2(new_n481), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(new_n866), .A3(new_n526), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n870), .A2(new_n871), .B1(new_n886), .B2(new_n867), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n879), .B1(new_n888), .B2(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n528), .A2(new_n530), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n882), .B1(new_n670), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT107), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n886), .A2(new_n867), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n874), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(KEYINPUT108), .A3(new_n853), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n889), .A2(new_n876), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n898), .A2(KEYINPUT40), .A3(new_n848), .A4(new_n851), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n878), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n563), .A2(new_n848), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(G330), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT109), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n446), .A2(new_n428), .A3(new_n686), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT106), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n876), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n906), .B(new_n907), .C1(new_n898), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n671), .A2(new_n858), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n558), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n686), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n810), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n850), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n911), .B1(new_n915), .B2(new_n877), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n904), .B1(new_n909), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n906), .ZN(new_n918));
  INV_X1    g0718(.A(new_n907), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n896), .A2(KEYINPUT108), .A3(new_n853), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT108), .B1(new_n896), .B2(new_n853), .ZN(new_n921));
  INV_X1    g0721(.A(new_n876), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n918), .B(new_n919), .C1(new_n923), .C2(KEYINPUT39), .ZN(new_n924));
  INV_X1    g0724(.A(new_n916), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(KEYINPUT109), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n903), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n563), .B1(new_n721), .B2(new_n712), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n673), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n266), .B2(new_n676), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT35), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n259), .B(new_n234), .C1(new_n584), .C2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(G116), .C1(new_n933), .C2(new_n584), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  OAI21_X1  g0736(.A(G77), .B1(new_n206), .B2(new_n490), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n232), .A2(new_n937), .B1(G50), .B2(new_n490), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(G1), .A3(new_n270), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT111), .ZN(G367));
  INV_X1    g0741(.A(new_n693), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n715), .B1(new_n591), .B2(new_n686), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n651), .A2(new_n595), .A3(new_n683), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n675), .A2(new_n694), .ZN(new_n948));
  INV_X1    g0748(.A(new_n943), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n948), .A2(KEYINPUT42), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT42), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n360), .A2(new_n362), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n594), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(new_n597), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n950), .A2(new_n951), .B1(new_n683), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n686), .A2(new_n611), .ZN(new_n956));
  MUX2_X1   g0756(.A(new_n714), .B(new_n650), .S(new_n956), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n955), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n955), .A2(new_n959), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n947), .B(new_n961), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n962), .B(KEYINPUT112), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n947), .B1(new_n967), .B2(new_n961), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n701), .B(KEYINPUT41), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n698), .B1(new_n943), .B2(new_n944), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT45), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT44), .B1(new_n699), .B2(new_n945), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n699), .A2(KEYINPUT44), .A3(new_n945), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(new_n942), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n695), .A2(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n695), .A2(KEYINPUT113), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n687), .C2(new_n694), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n692), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n735), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n976), .A2(new_n942), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n977), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n971), .B1(new_n985), .B2(new_n735), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n738), .A2(G1), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n969), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT117), .ZN(new_n989));
  INV_X1    g0789(.A(new_n742), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n754), .B1(new_n227), .B2(new_n550), .C1(new_n247), .C2(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n785), .A2(new_n206), .B1(new_n759), .B2(new_n422), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G50), .B2(new_n837), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT116), .B(G137), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n773), .A2(new_n369), .B1(new_n762), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G159), .B2(new_n824), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n783), .A2(G143), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n770), .A2(G68), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n998), .A2(new_n291), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n993), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n785), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT46), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n785), .B2(new_n276), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(new_n345), .C2(new_n777), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT115), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n782), .A2(new_n765), .B1(new_n762), .B2(new_n778), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n283), .B(new_n1008), .C1(G97), .C2(new_n760), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n767), .A2(new_n835), .B1(new_n769), .B2(new_n211), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT114), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n773), .A2(new_n292), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1000), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT47), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n739), .B1(new_n1016), .B2(new_n753), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n991), .B(new_n1017), .C1(new_n957), .C2(new_n756), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n988), .A2(new_n989), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n989), .B1(new_n988), .B2(new_n1018), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(G387));
  NOR2_X1   g0822(.A1(new_n687), .A2(new_n756), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n742), .B1(new_n244), .B2(new_n743), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n703), .B2(new_n747), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n546), .A2(new_n202), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G116), .B(new_n607), .C1(new_n1027), .C2(KEYINPUT50), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1028), .B(new_n743), .C1(KEYINPUT50), .C2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n490), .A2(new_n422), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n228), .A2(new_n211), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n753), .B(new_n752), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n763), .A2(G326), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G311), .A2(new_n824), .B1(new_n790), .B2(G317), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n292), .B2(new_n767), .C1(new_n774), .C2(new_n782), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n835), .B2(new_n769), .C1(new_n345), .C2(new_n785), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n283), .B(new_n1034), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n1039), .B2(new_n1038), .C1(new_n276), .C2(new_n759), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n283), .B1(new_n762), .B2(new_n369), .C1(new_n221), .C2(new_n759), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1001), .A2(G77), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n773), .B2(new_n202), .C1(new_n795), .C2(new_n782), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n602), .C2(new_n770), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n490), .B2(new_n767), .C1(new_n378), .C2(new_n777), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n801), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1023), .A2(new_n739), .A3(new_n1033), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n981), .B2(new_n987), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n701), .B1(new_n981), .B2(new_n735), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n983), .B2(new_n1050), .ZN(G393));
  NAND2_X1  g0851(.A1(new_n977), .A2(new_n984), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n982), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(new_n701), .A3(new_n985), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n977), .A2(new_n987), .A3(new_n984), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n754), .B1(new_n221), .B2(new_n227), .C1(new_n256), .C2(new_n990), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n546), .A2(new_n837), .B1(new_n824), .B2(G50), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT118), .Z(new_n1058));
  OAI22_X1  g0858(.A1(new_n782), .A2(new_n369), .B1(new_n773), .B2(new_n795), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n283), .B1(new_n759), .B2(new_n208), .C1(new_n490), .C2(new_n785), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G77), .B2(new_n770), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n763), .A2(G143), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n785), .A2(new_n835), .B1(new_n762), .B2(new_n774), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT119), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n291), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .C1(new_n211), .C2(new_n759), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT120), .Z(new_n1069));
  OAI22_X1  g0869(.A1(new_n782), .A2(new_n778), .B1(new_n773), .B2(new_n765), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n824), .A2(G303), .B1(new_n770), .B2(G116), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n767), .A2(new_n345), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1064), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n739), .B1(new_n1075), .B2(new_n753), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1056), .B(new_n1076), .C1(new_n945), .C2(new_n756), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1055), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1054), .A2(new_n1078), .ZN(G390));
  NAND2_X1  g0879(.A1(new_n719), .A2(new_n686), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n809), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n913), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n850), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n898), .A3(new_n906), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n809), .A2(G330), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n734), .A2(new_n850), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n907), .B1(new_n898), .B2(new_n908), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n915), .A2(new_n906), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1084), .B(new_n1086), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT121), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1084), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n848), .A2(new_n850), .A3(new_n1085), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n563), .A2(G330), .A3(new_n848), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n929), .A2(new_n1097), .A3(new_n673), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1082), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n848), .A2(new_n1085), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1086), .C1(new_n1100), .C2(new_n850), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n850), .B1(new_n734), .B2(new_n1085), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n914), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1098), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1096), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n919), .B1(new_n923), .B2(KEYINPUT39), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1088), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1108), .A2(new_n1091), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1090), .A2(KEYINPUT121), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n1104), .A4(new_n1095), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(new_n701), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1092), .A2(new_n987), .A3(new_n1095), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n821), .B(new_n792), .C1(G116), .C2(new_n790), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n837), .A2(G97), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n782), .A2(new_n835), .B1(new_n762), .B2(new_n345), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G107), .B2(new_n824), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n291), .B1(G77), .B2(new_n770), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G132), .A2(new_n790), .B1(new_n763), .B2(G125), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n202), .B2(new_n759), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n395), .B(new_n1122), .C1(G159), .C2(new_n770), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1125), .A2(new_n767), .B1(new_n777), .B2(new_n994), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT122), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n785), .A2(new_n369), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n782), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1120), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1133), .A2(new_n753), .B1(new_n378), .B2(new_n842), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n819), .B(new_n1134), .C1(new_n1087), .C2(new_n751), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1113), .A2(new_n1114), .A3(new_n1135), .ZN(G378));
  NAND2_X1  g0936(.A1(new_n414), .A2(new_n463), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT55), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n392), .A2(new_n858), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT56), .Z(new_n1141));
  OR2_X1    g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n878), .A2(new_n899), .A3(G330), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n917), .A2(new_n926), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n917), .B2(new_n926), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1145), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n904), .B(new_n916), .C1(new_n1087), .C2(new_n918), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT109), .B1(new_n924), .B2(new_n925), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1144), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n917), .A2(new_n926), .A3(new_n1145), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1148), .A2(new_n987), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n842), .A2(new_n202), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n773), .A2(new_n1131), .B1(new_n769), .B2(new_n369), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1001), .A2(new_n1124), .B1(new_n837), .B2(G137), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n830), .B2(new_n777), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G125), .C2(new_n783), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT59), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G41), .B1(new_n763), .B2(G124), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G33), .B1(new_n760), .B2(G159), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G116), .A2(new_n783), .B1(new_n824), .B2(G97), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n206), .B2(new_n759), .C1(new_n835), .C2(new_n762), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G107), .A2(new_n790), .B1(new_n837), .B2(new_n602), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1168), .A2(new_n294), .A3(new_n998), .A4(new_n1043), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1167), .A2(new_n283), .A3(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT58), .Z(new_n1171));
  OAI21_X1  g0971(.A(new_n202), .B1(new_n286), .B2(G41), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1165), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT123), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n739), .B1(new_n1174), .B2(new_n753), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1157), .B(new_n1175), .C1(new_n1144), .C2(new_n751), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1156), .A2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1153), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1098), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1111), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1148), .A2(new_n1182), .A3(KEYINPUT57), .A4(new_n1155), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n701), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1177), .B1(new_n1183), .B2(new_n1185), .ZN(G375));
  OR2_X1    g0986(.A1(new_n850), .A2(new_n751), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n785), .A2(new_n795), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n782), .A2(new_n830), .B1(new_n773), .B2(new_n994), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n824), .C2(new_n1124), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n283), .B1(new_n762), .B2(new_n1131), .C1(new_n206), .C2(new_n759), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G50), .B2(new_n770), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n369), .C2(new_n767), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n782), .A2(new_n345), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n221), .A2(new_n785), .B1(new_n773), .B2(new_n835), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G303), .B2(new_n763), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n422), .A2(new_n759), .B1(new_n767), .B2(new_n211), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G116), .B2(new_n824), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n770), .A2(new_n602), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1196), .A2(new_n1198), .A3(new_n395), .A4(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1193), .B1(new_n1194), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1201), .A2(new_n753), .B1(new_n490), .B2(new_n842), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1187), .A2(new_n819), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n987), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1101), .A2(new_n1103), .A3(new_n1098), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n970), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1207), .B2(new_n1104), .ZN(G381));
  INV_X1    g1008(.A(G375), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1114), .A2(new_n1135), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1212), .A2(G384), .A3(G381), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1021), .A3(new_n1214), .ZN(G407));
  OAI211_X1 g1015(.A(G407), .B(G213), .C1(G343), .C2(new_n1212), .ZN(G409));
  OAI211_X1 g1016(.A(G378), .B(new_n1177), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1148), .A2(new_n1182), .A3(new_n970), .A4(new_n1155), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n1156), .A3(new_n1176), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1211), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n682), .A2(G213), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1105), .B(new_n701), .C1(new_n1206), .C2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1206), .A2(new_n1224), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT124), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(new_n1228), .A3(G384), .A4(new_n1205), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1205), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1230));
  INV_X1    g1030(.A(G384), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT124), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1222), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(G2897), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1234), .B(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT61), .B1(new_n1223), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1234), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1221), .A2(new_n1222), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT62), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1235), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1243), .A3(new_n1239), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1238), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G390), .A2(new_n988), .A3(new_n1018), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(KEYINPUT126), .ZN(new_n1249));
  XOR2_X1   g1049(.A(G393), .B(G396), .Z(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(KEYINPUT126), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1247), .A2(new_n1249), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1248), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G390), .B1(new_n988), .B2(new_n1018), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1250), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1245), .A2(new_n1258), .ZN(new_n1259));
  AND4_X1   g1059(.A1(KEYINPUT63), .A2(new_n1221), .A3(new_n1222), .A4(new_n1239), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT63), .B1(new_n1242), .B2(new_n1239), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1223), .A2(KEYINPUT125), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1242), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1237), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1262), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1259), .A2(new_n1268), .ZN(G405));
  NAND2_X1  g1069(.A1(new_n1217), .A2(KEYINPUT127), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1239), .B1(new_n1209), .B2(G378), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G375), .A2(new_n1211), .A3(new_n1234), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1271), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1258), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1257), .B1(new_n1277), .B2(new_n1273), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(G402));
endmodule


