//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(KEYINPUT66), .B1(G567), .B2(new_n455), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n460), .B1(KEYINPUT66), .B2(new_n459), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n469), .A2(new_n470), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n464), .A2(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G137), .B1(G101), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n475), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n474), .A2(new_n464), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT69), .B(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n481), .A2(G126), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n490), .A2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT70), .B1(new_n499), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(new_n497), .A3(KEYINPUT5), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n506), .A2(new_n514), .ZN(G166));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  INV_X1    g091(.A(new_n498), .ZN(new_n517));
  NAND2_X1  g092(.A1(G63), .A2(G651), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n501), .B1(KEYINPUT5), .B2(new_n497), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n499), .A2(KEYINPUT70), .A3(G543), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n517), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(G51), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n522), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n500), .A2(new_n502), .ZN(new_n532));
  AND4_X1   g107(.A1(G89), .A2(new_n532), .A3(new_n517), .A4(new_n511), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n516), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n503), .A2(G89), .A3(new_n511), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n527), .A2(new_n530), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT71), .A4(new_n522), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(G168));
  XNOR2_X1  g113(.A(KEYINPUT73), .B(G90), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n503), .A2(new_n511), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n509), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n503), .B2(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT72), .B1(new_n544), .B2(new_n505), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  AOI211_X1 g122(.A(new_n547), .B(new_n498), .C1(new_n500), .C2(new_n502), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n546), .B(G651), .C1(new_n548), .C2(new_n543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n542), .B1(new_n545), .B2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n503), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n505), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n503), .A2(G81), .A3(new_n511), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n509), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XNOR2_X1  g134(.A(KEYINPUT74), .B(KEYINPUT8), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n509), .A2(new_n565), .A3(G53), .ZN(new_n566));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n532), .A2(G91), .A3(new_n517), .A4(new_n511), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n505), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  OAI21_X1  g150(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n509), .A2(G49), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n512), .ZN(G288));
  NAND2_X1  g154(.A1(new_n503), .A2(G61), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(new_n581), .B1(G73), .B2(G543), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n503), .A2(KEYINPUT76), .A3(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n505), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n509), .A2(G48), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n512), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n505), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n503), .A2(G85), .A3(new_n511), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT77), .B(G47), .Z(new_n593));
  NAND2_X1  g168(.A1(new_n509), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n592), .A2(KEYINPUT78), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(KEYINPUT78), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n532), .A2(G92), .A3(new_n517), .A4(new_n511), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n503), .A2(KEYINPUT10), .A3(G92), .A4(new_n511), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n509), .A2(G54), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT79), .B(G66), .Z(new_n605));
  AOI22_X1  g180(.A1(new_n503), .A2(new_n605), .B1(G79), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n606), .B2(new_n505), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT80), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G321));
  XNOR2_X1  g185(.A(G321), .B(KEYINPUT81), .ZN(G284));
  NOR2_X1   g186(.A1(G299), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g188(.A(new_n612), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n557), .ZN(G323));
  XOR2_X1   g194(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n620));
  XNOR2_X1  g195(.A(G323), .B(new_n620), .ZN(G282));
  OR2_X1    g196(.A1(new_n465), .A2(new_n466), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n476), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n475), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n481), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n464), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(KEYINPUT85), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(KEYINPUT85), .B2(new_n652), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n659), .C1(new_n654), .C2(new_n655), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n652), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n670), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n672), .A2(new_n673), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n670), .A2(new_n680), .A3(new_n674), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n670), .A2(new_n680), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n678), .A2(new_n679), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G229));
  XNOR2_X1  g264(.A(KEYINPUT98), .B(KEYINPUT31), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G11), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT30), .B(G28), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n481), .A2(G129), .ZN(new_n695));
  NAND3_X1  g270(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT26), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n475), .A2(G141), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n476), .A2(G105), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(new_n692), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n692), .B2(G32), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n694), .B1(new_n692), .B2(new_n633), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G164), .A2(new_n692), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n692), .A2(G27), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT99), .Z(new_n709));
  NOR3_X1   g284(.A1(new_n707), .A2(G2078), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G19), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n557), .B2(new_n712), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1341), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n692), .A2(G26), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n475), .A2(G140), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n481), .A2(G128), .ZN(new_n719));
  OR2_X1    g294(.A1(G104), .A2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n717), .B1(new_n723), .B2(new_n692), .ZN(new_n724));
  INV_X1    g299(.A(G2067), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(G2078), .B1(new_n707), .B2(new_n709), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n711), .A2(new_n715), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n712), .A2(G20), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT23), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n565), .B1(new_n509), .B2(G53), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n570), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n532), .A2(G65), .A3(new_n517), .ZN(new_n734));
  NAND2_X1  g309(.A1(G78), .A2(G543), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n505), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(new_n712), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1956), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n692), .B1(new_n740), .B2(G34), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(G34), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT96), .Z(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n478), .B2(new_n692), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n728), .A2(new_n739), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n692), .A2(G35), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT100), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n485), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT102), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n704), .A2(new_n705), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n475), .A2(G139), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n622), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n763), .B(new_n764), .C1(new_n464), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT94), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  NOR2_X1   g343(.A1(G29), .A2(G33), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT92), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n768), .A2(G2072), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(G2072), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n756), .B2(new_n755), .ZN(new_n773));
  AND4_X1   g348(.A1(new_n758), .A2(new_n760), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G21), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G168), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n712), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n712), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n780), .B1(G1961), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G1961), .B2(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n712), .A2(G4), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n609), .B2(new_n712), .ZN(new_n787));
  INV_X1    g362(.A(G1348), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n750), .A2(new_n774), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G22), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n791), .A2(KEYINPUT91), .A3(G16), .ZN(new_n792));
  OAI21_X1  g367(.A(KEYINPUT91), .B1(new_n791), .B2(G16), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(G166), .C2(new_n712), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  MUX2_X1   g370(.A(G23), .B(G288), .S(G16), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT33), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G1976), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(G1976), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n712), .A2(G6), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n588), .B2(new_n712), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT90), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT32), .B(G1981), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n800), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n800), .A2(new_n805), .A3(new_n809), .A4(new_n806), .ZN(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G24), .ZN(new_n811));
  XNOR2_X1  g386(.A(G290), .B(KEYINPUT89), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1986), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n692), .A2(G25), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n475), .A2(G131), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n481), .A2(G119), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n464), .A2(G107), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT88), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n815), .B1(new_n825), .B2(new_n692), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G1991), .Z(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n814), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n808), .A2(new_n810), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n808), .A2(new_n833), .A3(new_n810), .A4(new_n830), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n790), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(G311));
  INV_X1    g412(.A(new_n835), .ZN(G150));
  NAND2_X1  g413(.A1(new_n609), .A2(G559), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n532), .A2(G67), .A3(new_n517), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G651), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n532), .A2(G93), .A3(new_n517), .A4(new_n511), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n509), .A2(G55), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n847), .A3(KEYINPUT105), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n555), .B(new_n554), .C1(new_n849), .C2(new_n505), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n505), .B1(new_n840), .B2(new_n841), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(new_n846), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n848), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n852), .A2(new_n846), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n557), .A2(KEYINPUT105), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n839), .B(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  OAI21_X1  g438(.A(G860), .B1(new_n852), .B2(new_n846), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  NAND2_X1  g441(.A1(new_n767), .A2(KEYINPUT106), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n702), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n481), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n464), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(G142), .B2(new_n475), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n624), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n868), .B(new_n874), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n490), .A2(new_n495), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n723), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n825), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n868), .B(new_n874), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n478), .B(new_n633), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n485), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n880), .A2(new_n888), .A3(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g466(.A1(new_n855), .A2(G868), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G166), .A2(G288), .ZN(new_n894));
  INV_X1    g469(.A(new_n512), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n895), .A2(G87), .B1(G49), .B2(new_n509), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(new_n576), .C1(new_n506), .C2(new_n514), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G290), .ZN(new_n900));
  NAND2_X1  g475(.A1(G305), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n588), .A2(G290), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n899), .A3(new_n902), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(KEYINPUT108), .B2(KEYINPUT42), .ZN(new_n907));
  NAND2_X1  g482(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n907), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n854), .A2(new_n856), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n617), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n737), .B1(new_n603), .B2(new_n607), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  INV_X1    g489(.A(new_n604), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n503), .A2(new_n605), .ZN(new_n916));
  NAND2_X1  g491(.A1(G79), .A2(G543), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n918), .B2(G651), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n601), .A2(new_n602), .ZN(new_n920));
  NAND3_X1  g495(.A1(G299), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n608), .A2(KEYINPUT107), .A3(G299), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n913), .A2(new_n927), .A3(new_n921), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n912), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n910), .A2(new_n925), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n907), .B(new_n908), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n925), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G868), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n893), .B1(new_n936), .B2(new_n937), .ZN(G295));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n939), .B(new_n893), .C1(new_n936), .C2(new_n937), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n932), .B2(new_n935), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT109), .B1(new_n941), .B2(new_n892), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(G331));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n901), .A2(new_n899), .A3(new_n902), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(new_n903), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n534), .A2(new_n947), .A3(new_n537), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n534), .B2(new_n537), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n948), .A2(new_n949), .A3(G171), .ZN(new_n950));
  AND3_X1   g525(.A1(G171), .A2(G168), .A3(KEYINPUT110), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n911), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n924), .ZN(new_n953));
  NAND2_X1  g528(.A1(G168), .A2(KEYINPUT110), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n534), .A2(new_n947), .A3(new_n537), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(G301), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(G171), .A2(G168), .A3(KEYINPUT110), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n857), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n952), .A2(new_n953), .A3(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n950), .A2(new_n911), .A3(new_n951), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n956), .A2(new_n957), .B1(new_n856), .B2(new_n854), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(KEYINPUT111), .B(new_n959), .C1(new_n962), .C2(new_n929), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n952), .A2(new_n958), .A3(new_n953), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n946), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n913), .A2(new_n921), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT41), .B(new_n967), .C1(new_n960), .C2(new_n961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n946), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n952), .A2(new_n958), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n953), .B1(new_n970), .B2(KEYINPUT41), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n887), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n959), .A2(KEYINPUT111), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n929), .B1(new_n958), .B2(new_n952), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n946), .B(new_n965), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n979), .A2(new_n887), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n965), .B1(new_n977), .B2(new_n978), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT43), .B1(new_n981), .B2(new_n906), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n976), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT112), .B(KEYINPUT43), .C1(new_n966), .C2(new_n972), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n975), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n982), .B(new_n887), .C1(new_n971), .C2(new_n969), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n887), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT43), .B1(new_n987), .B2(new_n966), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT44), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n944), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n988), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n976), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n975), .A2(new_n983), .A3(new_n984), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(KEYINPUT113), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(G397));
  NAND4_X1  g570(.A1(new_n473), .A2(KEYINPUT114), .A3(G40), .A4(new_n477), .ZN(new_n996));
  OAI211_X1 g571(.A(G40), .B(new_n477), .C1(new_n471), .C2(new_n472), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n490), .B2(new_n495), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n588), .B2(new_n1006), .ZN(new_n1007));
  NOR4_X1   g582(.A1(new_n584), .A2(KEYINPUT118), .A3(G1981), .A4(new_n587), .ZN(new_n1008));
  OAI22_X1  g583(.A1(new_n1007), .A2(new_n1008), .B1(new_n1006), .B2(new_n588), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1003), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(new_n1004), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT55), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1001), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n996), .A2(new_n999), .B1(KEYINPUT50), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1001), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n756), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1971), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT116), .B(new_n1023), .C1(G164), .C2(G1384), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1001), .A2(KEYINPUT45), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n997), .B(KEYINPUT114), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1022), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1016), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1017), .B1(new_n996), .B2(new_n999), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT117), .B(G1976), .Z(new_n1033));
  AND2_X1   g608(.A1(G288), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G288), .A2(new_n1036), .ZN(new_n1037));
  NOR4_X1   g612(.A1(new_n1032), .A2(new_n1035), .A3(new_n1016), .A4(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1002), .B(G8), .C1(new_n1036), .C2(G288), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(KEYINPUT52), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1012), .A2(new_n1015), .A3(new_n1031), .A4(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1042));
  XOR2_X1   g617(.A(new_n1042), .B(KEYINPUT120), .Z(new_n1043));
  NOR2_X1   g618(.A1(G288), .A2(G1976), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1012), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1003), .B(KEYINPUT119), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1020), .B(KEYINPUT121), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1049), .A2(new_n1018), .A3(new_n756), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1024), .A2(new_n1027), .A3(new_n1026), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1971), .B1(new_n1051), .B2(new_n1000), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1014), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1031), .A2(new_n1015), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1012), .A4(new_n1040), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1001), .B(new_n1023), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1000), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n777), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1018), .A2(new_n748), .A3(new_n1020), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(G8), .A3(G168), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1048), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1012), .A2(new_n1040), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1031), .A2(new_n1015), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1062), .A2(new_n1048), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1055), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1047), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1061), .B2(G286), .ZN(new_n1069));
  AOI21_X1  g644(.A(G168), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT51), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(G8), .C1(new_n1061), .C2(G286), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT62), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1071), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1056), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1028), .A2(new_n1029), .A3(G2078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(KEYINPUT53), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1081));
  INV_X1    g656(.A(G1961), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT53), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1080), .B(new_n1083), .C1(new_n1058), .C2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .A4(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1002), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1028), .A2(new_n1029), .A3(G1996), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n557), .B(new_n1089), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1081), .A2(new_n788), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1032), .A2(new_n725), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n608), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1093), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n850), .B1(new_n1099), .B2(new_n1091), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT123), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1094), .B(new_n1098), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1095), .B(new_n1097), .C1(new_n603), .C2(new_n607), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1097), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1348), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n608), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1096), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n737), .B(KEYINPUT57), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1051), .A2(new_n1000), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1956), .B1(new_n1049), .B2(new_n1018), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1049), .A2(new_n1018), .ZN(new_n1115));
  INV_X1    g690(.A(G1956), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1111), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1119), .A3(new_n1109), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT61), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1103), .A2(new_n1108), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1109), .B(KEYINPUT122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n1120), .A3(KEYINPUT61), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1124), .A2(new_n1120), .A3(KEYINPUT124), .A4(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1107), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1122), .A2(new_n1129), .B1(new_n1120), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(G171), .B(KEYINPUT54), .Z(new_n1132));
  AND2_X1   g707(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1133));
  INV_X1    g708(.A(new_n469), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n477), .A2(G40), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1085), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1132), .B1(new_n1057), .B2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1086), .A2(new_n1132), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1078), .A3(new_n1074), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1068), .B(new_n1088), .C1(new_n1131), .C2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1001), .A2(KEYINPUT45), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1000), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n824), .B(new_n827), .ZN(new_n1147));
  INV_X1    g722(.A(G1996), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n702), .B(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n722), .B(new_n725), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1986), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n900), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n900), .A2(new_n1155), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT115), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1146), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1143), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT48), .B1(new_n1158), .B2(new_n1146), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1158), .A2(KEYINPUT48), .A3(new_n1146), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1161), .B(new_n1162), .C1(new_n1146), .C2(new_n1153), .ZN(new_n1163));
  INV_X1    g738(.A(new_n702), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1146), .B1(new_n1164), .B2(new_n1151), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT46), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1145), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT47), .Z(new_n1170));
  NOR2_X1   g745(.A1(new_n824), .A2(new_n828), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(KEYINPUT126), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1152), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n1173), .A2(new_n1175), .B1(G2067), .B2(new_n722), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1163), .B(new_n1170), .C1(new_n1146), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1160), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(new_n650), .ZN(new_n1180));
  NOR4_X1   g754(.A1(G229), .A2(new_n462), .A3(new_n1180), .A4(G227), .ZN(new_n1181));
  NAND3_X1  g755(.A1(new_n1181), .A2(new_n890), .A3(new_n991), .ZN(G225));
  INV_X1    g756(.A(G225), .ZN(G308));
endmodule


