//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT72), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT72), .ZN(new_n192));
  OAI21_X1  g006(.A(G140), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(G125), .A2(G140), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n188), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT72), .B(G125), .ZN(new_n197));
  INV_X1    g011(.A(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n188), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n187), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT73), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n191), .A2(KEYINPUT72), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n189), .A2(G125), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT16), .B1(new_n205), .B2(new_n194), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n204), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n188), .A3(new_n198), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(G146), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n201), .A2(new_n202), .A3(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(KEYINPUT73), .B(new_n187), .C1(new_n196), .C2(new_n200), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(G128), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT66), .A2(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT23), .B1(new_n217), .B2(G119), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(G119), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n215), .B2(G119), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT24), .B(G110), .Z(new_n223));
  AOI22_X1  g037(.A1(new_n221), .A2(G110), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n210), .A2(new_n211), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT74), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n209), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n200), .B1(new_n228), .B2(KEYINPUT16), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT74), .A3(G146), .ZN(new_n230));
  OAI22_X1  g044(.A1(new_n221), .A2(G110), .B1(new_n222), .B2(new_n223), .ZN(new_n231));
  XNOR2_X1  g045(.A(G125), .B(G140), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n187), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n227), .A2(new_n230), .A3(new_n231), .A4(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n225), .A2(KEYINPUT75), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT75), .B1(new_n225), .B2(new_n234), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G137), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n238), .A2(G221), .A3(G234), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n237), .B(new_n239), .Z(new_n240));
  NOR3_X1   g054(.A1(new_n235), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n225), .A2(new_n234), .A3(new_n240), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT25), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n225), .A2(new_n234), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n225), .A2(KEYINPUT75), .A3(new_n234), .ZN(new_n249));
  INV_X1    g063(.A(new_n240), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n252), .A3(new_n243), .A4(new_n242), .ZN(new_n253));
  INV_X1    g067(.A(G217), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(G234), .B2(new_n243), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n245), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(G902), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n251), .A2(new_n242), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n259), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n256), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n187), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT0), .A3(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT11), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(G137), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G131), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n282), .A3(new_n279), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n272), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G119), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G116), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G119), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT2), .B(G113), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n289), .A2(new_n293), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n266), .A2(KEYINPUT1), .A3(new_n217), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT1), .B1(new_n264), .B2(G146), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n263), .A2(KEYINPUT65), .A3(KEYINPUT1), .ZN(new_n303));
  OR2_X1    g117(.A1(KEYINPUT66), .A2(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n212), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n266), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(KEYINPUT67), .A3(new_n266), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n299), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT64), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n279), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n273), .B2(G137), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n279), .A2(new_n312), .ZN(new_n315));
  OAI21_X1  g129(.A(G131), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n283), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n298), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT69), .ZN(new_n319));
  INV_X1    g133(.A(new_n284), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n311), .B2(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n297), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n298), .B(new_n323), .C1(new_n311), .C2(new_n317), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n319), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT28), .ZN(new_n326));
  INV_X1    g140(.A(new_n299), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n306), .A2(KEYINPUT67), .A3(new_n266), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT67), .B1(new_n306), .B2(new_n266), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n317), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT28), .B1(new_n332), .B2(new_n298), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G237), .A2(G953), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G210), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT27), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(G101), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n326), .A2(new_n335), .A3(KEYINPUT29), .A4(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n340), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n286), .A2(new_n288), .A3(new_n291), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n291), .B1(new_n286), .B2(new_n288), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n295), .B1(new_n345), .B2(new_n293), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n321), .A2(KEYINPUT30), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(new_n348), .A3(new_n320), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n319), .A2(new_n324), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n342), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n333), .B(new_n342), .C1(new_n325), .C2(KEYINPUT28), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n341), .B(new_n243), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n319), .A2(new_n324), .A3(new_n340), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT31), .B1(new_n350), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n348), .B1(new_n332), .B2(new_n320), .ZN(new_n359));
  AOI211_X1 g173(.A(KEYINPUT30), .B(new_n284), .C1(new_n330), .C2(new_n331), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n297), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n324), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n323), .B1(new_n332), .B2(new_n298), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n361), .A2(new_n364), .A3(new_n340), .A4(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n333), .B1(new_n325), .B2(KEYINPUT28), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n358), .B(new_n366), .C1(new_n367), .C2(new_n340), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n369), .A2(G472), .A3(G902), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n356), .A2(G472), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G472), .A2(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n358), .A2(new_n366), .ZN(new_n373));
  INV_X1    g187(.A(new_n333), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n340), .B1(new_n326), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n372), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n369), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n262), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n304), .A2(G143), .A3(new_n212), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n264), .A2(G128), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n273), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n273), .B1(new_n380), .B2(new_n381), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n384), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT90), .A3(new_n382), .ZN(new_n387));
  INV_X1    g201(.A(G122), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n287), .A2(G122), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n389), .B2(KEYINPUT14), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n391), .B(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n389), .A2(new_n390), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n392), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n382), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT13), .B1(new_n264), .B2(G128), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n264), .A2(KEYINPUT13), .A3(G128), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n264), .A2(KEYINPUT13), .A3(G128), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT88), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n405), .A3(new_n380), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G134), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT89), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n215), .A2(G143), .B1(new_n404), .B2(KEYINPUT88), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n273), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n382), .A2(new_n396), .A3(new_n398), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT89), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n395), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT9), .B(G234), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n415), .A2(new_n254), .A3(G953), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n412), .B1(new_n410), .B2(new_n411), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n399), .A2(new_n407), .A3(KEYINPUT89), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n395), .A3(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n243), .ZN(new_n424));
  INV_X1    g238(.A(G478), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT15), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n424), .B(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  INV_X1    g242(.A(G104), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(G143), .B1(new_n336), .B2(G214), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n436));
  INV_X1    g250(.A(new_n434), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n432), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n436), .A2(new_n282), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n435), .A2(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n233), .B1(new_n228), .B2(new_n187), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT82), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n443), .B(new_n233), .C1(new_n228), .C2(new_n187), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n210), .A2(new_n211), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT17), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n435), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n437), .A2(new_n282), .A3(new_n432), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n435), .A2(new_n449), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT85), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n435), .A2(new_n449), .A3(new_n452), .A4(new_n447), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n431), .B(new_n445), .C1(new_n446), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n445), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT19), .B(new_n195), .C1(new_n197), .C2(new_n198), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT19), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n232), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n187), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT83), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n457), .A2(new_n462), .A3(new_n187), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n464), .A2(KEYINPUT84), .A3(new_n227), .A4(new_n230), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n435), .A2(new_n449), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT74), .B1(new_n229), .B2(G146), .ZN(new_n468));
  AND4_X1   g282(.A1(KEYINPUT74), .A2(new_n206), .A3(G146), .A4(new_n208), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT84), .B1(new_n470), .B2(new_n464), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n456), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n455), .B1(new_n472), .B2(new_n431), .ZN(new_n473));
  NOR2_X1   g287(.A1(G475), .A2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT20), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n478));
  INV_X1    g292(.A(new_n464), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n227), .A2(new_n230), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n466), .A3(new_n465), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n430), .B1(new_n482), .B2(new_n456), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n477), .B(new_n474), .C1(new_n483), .C2(new_n455), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n446), .A2(new_n454), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(new_n431), .C1(new_n487), .C2(new_n445), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n445), .B1(new_n446), .B2(new_n454), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT86), .B1(new_n489), .B2(new_n430), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n455), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G475), .B1(new_n491), .B2(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n492), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n427), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  AND2_X1   g313(.A1(KEYINPUT77), .A2(G101), .ZN(new_n500));
  NOR2_X1   g314(.A1(KEYINPUT77), .A2(G101), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT3), .B1(new_n429), .B2(G107), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n429), .A2(G107), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT3), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n392), .A3(G104), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n508));
  XNOR2_X1  g322(.A(G104), .B(G107), .ZN(new_n509));
  INV_X1    g323(.A(G101), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n392), .A2(G104), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n504), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT78), .A3(G101), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT10), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n330), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n270), .B1(G128), .B2(new_n300), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n299), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n516), .B1(new_n520), .B2(new_n515), .ZN(new_n521));
  INV_X1    g335(.A(new_n272), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT4), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n503), .A2(new_n506), .A3(new_n504), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G101), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n525), .B2(new_n507), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT4), .B1(new_n524), .B2(G101), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n281), .A2(new_n283), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT79), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT79), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n281), .A2(new_n283), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n518), .A2(new_n521), .A3(new_n528), .A4(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT80), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G140), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n238), .A2(G227), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n327), .B(new_n515), .C1(new_n328), .C2(new_n329), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n520), .A2(new_n515), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT12), .B1(new_n543), .B2(new_n529), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n545));
  INV_X1    g359(.A(new_n529), .ZN(new_n546));
  AOI211_X1 g360(.A(new_n545), .B(new_n546), .C1(new_n541), .C2(new_n542), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n535), .B1(new_n534), .B2(new_n539), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n540), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n330), .A2(new_n517), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n528), .A2(new_n521), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n529), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n539), .B1(new_n553), .B2(new_n534), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n499), .B(new_n243), .C1(new_n550), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n499), .A2(new_n243), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n534), .B1(new_n544), .B2(new_n547), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n534), .A2(new_n539), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n557), .A2(new_n538), .B1(new_n558), .B2(new_n553), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n556), .B1(new_n559), .B2(G469), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G214), .B1(G237), .B2(G902), .ZN(new_n562));
  XNOR2_X1  g376(.A(G110), .B(G122), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n297), .B1(new_n526), .B2(new_n527), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G113), .B1(new_n286), .B2(KEYINPUT5), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n290), .A2(new_n292), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(KEYINPUT5), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n569), .A2(new_n295), .A3(new_n515), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n564), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT5), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n290), .B2(new_n292), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n296), .B1(new_n573), .B2(new_n567), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n565), .B(new_n563), .C1(new_n515), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(KEYINPUT6), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n564), .C1(new_n566), .C2(new_n570), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n522), .A2(new_n207), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n311), .B2(new_n207), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(G224), .A3(new_n238), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n238), .A2(G224), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n582), .B(new_n579), .C1(new_n311), .C2(new_n207), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n576), .A2(new_n578), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(KEYINPUT7), .A3(new_n582), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(KEYINPUT7), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n579), .B(new_n586), .C1(new_n311), .C2(new_n207), .ZN(new_n587));
  INV_X1    g401(.A(new_n515), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n289), .A2(new_n572), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n296), .B1(new_n589), .B2(new_n567), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n563), .B(KEYINPUT8), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n591), .B(new_n592), .C1(new_n574), .C2(new_n588), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n585), .A2(new_n575), .A3(new_n587), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n584), .A2(new_n243), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(G210), .B1(G237), .B2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n587), .A2(new_n575), .A3(new_n593), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n599), .B2(new_n585), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n584), .A3(new_n596), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND4_X1   g416(.A1(new_n498), .A2(new_n561), .A3(new_n562), .A4(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G952), .ZN(new_n604));
  AOI211_X1 g418(.A(G953), .B(new_n604), .C1(G234), .C2(G237), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT21), .B(G898), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT91), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n243), .B(new_n238), .C1(G234), .C2(G237), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n378), .A2(new_n497), .A3(new_n603), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT92), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n502), .ZN(G3));
  NAND4_X1  g428(.A1(new_n600), .A2(KEYINPUT93), .A3(new_n584), .A4(new_n596), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n615), .A2(new_n562), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT93), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n598), .A2(new_n617), .A3(new_n601), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n616), .A2(new_n618), .A3(new_n611), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT96), .B(G478), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n424), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n425), .A2(G902), .ZN(new_n622));
  INV_X1    g436(.A(new_n422), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n416), .B1(new_n421), .B2(new_n395), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT33), .B1(new_n624), .B2(KEYINPUT94), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n418), .B(new_n422), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n622), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(KEYINPUT95), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT95), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n423), .B(KEYINPUT33), .C1(KEYINPUT94), .C2(new_n624), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n630), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n636), .B2(new_n622), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n621), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n619), .A2(new_n495), .A3(new_n496), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT97), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n492), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT87), .B1(new_n485), .B2(new_n492), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n643), .A2(new_n644), .A3(new_n638), .A4(new_n619), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n256), .A2(new_n260), .A3(new_n261), .ZN(new_n647));
  INV_X1    g461(.A(new_n498), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n555), .B2(new_n560), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n368), .A2(new_n243), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G472), .ZN(new_n651));
  AND4_X1   g465(.A1(new_n376), .A2(new_n647), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT98), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NAND2_X1  g470(.A1(new_n616), .A2(new_n618), .ZN(new_n657));
  INV_X1    g471(.A(new_n427), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n657), .A2(new_n493), .A3(new_n610), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n651), .A2(new_n376), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n248), .B(new_n249), .C1(KEYINPUT36), .C2(new_n250), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n250), .A2(KEYINPUT36), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n235), .B2(new_n236), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n664), .A2(new_n257), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n256), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n497), .A3(new_n603), .A4(new_n611), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  NAND2_X1  g487(.A1(new_n356), .A2(G472), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n368), .A2(new_n370), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n377), .A3(new_n675), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n561), .A2(new_n498), .A3(new_n668), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n605), .B1(new_n609), .B2(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n493), .A2(new_n658), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n616), .A2(new_n618), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n676), .A2(new_n677), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n679), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n649), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT40), .Z(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n602), .B(new_n687), .Z(new_n688));
  NAND3_X1  g502(.A1(new_n669), .A2(new_n427), .A3(new_n562), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n340), .B1(new_n364), .B2(new_n322), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n350), .A2(new_n357), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n243), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G472), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n675), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT32), .B1(new_n368), .B2(new_n372), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n688), .A2(new_n689), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n686), .A2(new_n643), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  INV_X1    g513(.A(new_n679), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n495), .A2(new_n638), .A3(new_n496), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n561), .A2(new_n668), .A3(new_n498), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n377), .B2(new_n371), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n704), .A3(new_n681), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n534), .A2(new_n539), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n520), .A2(new_n515), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n311), .B2(new_n515), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n545), .B1(new_n710), .B2(new_n546), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n543), .A2(KEYINPUT12), .A3(new_n529), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n708), .A2(KEYINPUT80), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n554), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(G902), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT100), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n555), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT100), .B(G469), .C1(new_n715), .C2(G902), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n648), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n676), .A3(new_n647), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n707), .B1(new_n646), .B2(new_n722), .ZN(new_n723));
  AOI211_X1 g537(.A(KEYINPUT101), .B(new_n721), .C1(new_n640), .C2(new_n645), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT102), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n725), .B(new_n727), .ZN(G15));
  NAND3_X1  g542(.A1(new_n659), .A2(new_n378), .A3(new_n720), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  AND2_X1   g544(.A1(new_n720), .A2(new_n681), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n669), .B1(new_n371), .B2(new_n377), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n611), .A3(new_n497), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  NAND3_X1  g548(.A1(new_n616), .A2(new_n618), .A3(new_n427), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n495), .A3(new_n496), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n340), .B1(new_n326), .B2(new_n335), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n372), .B1(new_n373), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT104), .B(G472), .Z(new_n742));
  NAND2_X1  g556(.A1(new_n650), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT103), .B(new_n372), .C1(new_n373), .C2(new_n738), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n647), .A2(new_n741), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n737), .A2(new_n745), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n610), .B(new_n648), .C1(new_n718), .C2(new_n719), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT105), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n745), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n641), .A2(new_n735), .A3(new_n642), .ZN(new_n750));
  AND4_X1   g564(.A1(KEYINPUT105), .A2(new_n749), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n388), .ZN(G24));
  NAND2_X1  g567(.A1(new_n720), .A2(new_n681), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n741), .A2(new_n743), .A3(new_n668), .A4(new_n744), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n754), .A2(new_n701), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n191), .ZN(G27));
  OR2_X1    g571(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n371), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n598), .A2(new_n498), .A3(new_n562), .A4(new_n601), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n708), .A2(KEYINPUT80), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n711), .A2(new_n712), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n714), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n554), .ZN(new_n765));
  AOI21_X1  g579(.A(G902), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n556), .B1(new_n766), .B2(new_n499), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  INV_X1    g582(.A(new_n557), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n539), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n558), .A2(new_n553), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n557), .A2(KEYINPUT106), .A3(new_n538), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(G469), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n761), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT42), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n702), .A2(new_n760), .A3(new_n775), .A4(new_n647), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n676), .A2(new_n647), .A3(new_n774), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n777), .B1(new_n778), .B2(new_n701), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  NAND4_X1  g595(.A1(new_n676), .A2(new_n680), .A3(new_n647), .A4(new_n774), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n378), .A2(KEYINPUT108), .A3(new_n680), .A4(new_n774), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NOR2_X1   g601(.A1(new_n559), .A2(KEYINPUT45), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n499), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n770), .A2(KEYINPUT45), .A3(new_n771), .A4(new_n772), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n556), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n555), .B1(new_n791), .B2(KEYINPUT46), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n498), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  INV_X1    g609(.A(new_n684), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n562), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n602), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT43), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n495), .A2(new_n496), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n638), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(new_n807), .A3(new_n663), .A4(new_n668), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n802), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n799), .B(new_n810), .C1(new_n809), .C2(new_n808), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT110), .B(G137), .Z(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G39));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n794), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(KEYINPUT47), .B(new_n498), .C1(new_n792), .C2(new_n793), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n676), .A2(new_n647), .A3(new_n802), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n702), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT111), .B(G140), .Z(new_n820));
  XNOR2_X1  g634(.A(new_n819), .B(new_n820), .ZN(G42));
  OAI211_X1 g635(.A(new_n729), .B(new_n733), .C1(new_n748), .C2(new_n751), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n725), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n679), .A2(new_n648), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n256), .A2(new_n667), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n368), .A2(new_n370), .B1(new_n692), .B2(G472), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n825), .B1(new_n377), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n767), .A2(new_n773), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n643), .A2(new_n827), .A3(new_n736), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n676), .A2(new_n677), .A3(new_n681), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n829), .B(new_n682), .C1(new_n701), .C2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT114), .B1(new_n831), .B2(new_n756), .ZN(new_n832));
  INV_X1    g646(.A(new_n825), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n828), .B(new_n833), .C1(new_n695), .C2(new_n694), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n657), .A2(new_n493), .A3(new_n658), .A4(new_n679), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n750), .A2(new_n835), .B1(new_n704), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n701), .A2(new_n755), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n731), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .A4(new_n705), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n632), .A2(KEYINPUT95), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n636), .A2(new_n634), .A3(new_n622), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n845), .A2(new_n846), .B1(new_n424), .B2(new_n620), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n643), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n805), .A2(new_n658), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n610), .B(new_n800), .C1(new_n598), .C2(new_n601), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n849), .A3(new_n652), .A4(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n851), .A2(new_n612), .A3(new_n671), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n776), .A2(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n802), .A2(new_n427), .A3(new_n493), .A4(new_n679), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n839), .A2(new_n774), .B1(new_n854), .B2(new_n704), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n832), .A2(KEYINPUT52), .A3(new_n841), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n823), .A2(new_n844), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n832), .B2(new_n841), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n831), .A2(new_n756), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n843), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n823), .A4(new_n856), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n865), .A3(KEYINPUT54), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n844), .A2(new_n857), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n641), .A2(new_n847), .A3(new_n642), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n644), .B1(new_n868), .B2(new_n619), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n639), .A2(KEYINPUT97), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n722), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT101), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n646), .A2(new_n707), .A3(new_n722), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n732), .A2(new_n497), .A3(new_n611), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n729), .B1(new_n875), .B2(new_n754), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n746), .A2(new_n747), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT105), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n746), .A2(KEYINPUT105), .A3(new_n747), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n856), .A2(new_n874), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n864), .B1(new_n867), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n864), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n725), .B2(new_n822), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n874), .A2(KEYINPUT115), .A3(new_n881), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n863), .A2(new_n885), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n647), .A2(new_n605), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n720), .A3(new_n696), .A4(new_n801), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n643), .A2(new_n638), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n720), .A2(new_n801), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n804), .A3(new_n807), .A4(new_n605), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n755), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n804), .A2(new_n807), .A3(new_n605), .A4(new_n749), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n688), .A2(new_n800), .A3(new_n720), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT50), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n900), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(KEYINPUT117), .A3(new_n801), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n900), .B2(new_n802), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n718), .A2(new_n719), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n648), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n815), .A2(new_n816), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n907), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n905), .A2(KEYINPUT51), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n804), .A2(new_n807), .A3(new_n605), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT48), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n760), .A2(new_n647), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n915), .A2(new_n916), .A3(new_n918), .A4(new_n897), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT48), .B1(new_n898), .B2(new_n917), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n868), .ZN(new_n922));
  OAI211_X1 g736(.A(G952), .B(new_n238), .C1(new_n893), .C2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n906), .B2(new_n731), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n921), .A2(KEYINPUT119), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT119), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n914), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n911), .B(KEYINPUT118), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n907), .B(new_n909), .C1(new_n817), .C2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT51), .B1(new_n905), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n866), .A2(new_n891), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n604), .A2(new_n238), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR4_X1    g748(.A1(new_n262), .A2(new_n803), .A3(new_n648), .A4(new_n800), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT112), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT49), .ZN(new_n937));
  OAI22_X1  g751(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n910), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n936), .B2(new_n935), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT113), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n910), .A2(new_n937), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n940), .A2(new_n696), .A3(new_n688), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT120), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n934), .A2(new_n945), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(G75));
  NOR2_X1   g761(.A1(new_n238), .A2(G952), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n243), .B1(new_n883), .B2(new_n889), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT56), .B1(new_n950), .B2(G210), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n576), .A2(new_n578), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n581), .A2(new_n583), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n584), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT55), .Z(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  NOR4_X1   g771(.A1(new_n860), .A2(new_n884), .A3(new_n862), .A4(new_n864), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n725), .A2(new_n822), .A3(new_n886), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT115), .B1(new_n874), .B2(new_n881), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI22_X1  g775(.A1(new_n958), .A2(new_n961), .B1(new_n858), .B2(new_n864), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT121), .B1(new_n962), .B2(new_n243), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n883), .A2(new_n889), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n965), .A3(G902), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n597), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n956), .A2(KEYINPUT122), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n956), .A2(KEYINPUT122), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT56), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n957), .B1(new_n967), .B2(new_n970), .ZN(G51));
  INV_X1    g785(.A(new_n890), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(new_n891), .ZN(new_n974));
  XOR2_X1   g788(.A(KEYINPUT123), .B(KEYINPUT57), .Z(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(new_n556), .ZN(new_n976));
  OAI22_X1  g790(.A1(new_n974), .A2(new_n976), .B1(new_n554), .B2(new_n550), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n963), .A2(new_n790), .A3(new_n966), .A4(new_n789), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n948), .B1(new_n977), .B2(new_n978), .ZN(G54));
  AND2_X1   g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n963), .A2(new_n966), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n473), .ZN(new_n982));
  INV_X1    g796(.A(new_n473), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n963), .A2(new_n983), .A3(new_n966), .A4(new_n980), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n982), .A2(new_n949), .A3(new_n984), .ZN(G60));
  XNOR2_X1  g799(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n425), .A2(new_n243), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n866), .B2(new_n891), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n949), .B1(new_n990), .B2(new_n636), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT125), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n973), .A2(new_n891), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n636), .A2(new_n988), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g810(.A(KEYINPUT125), .B(new_n994), .C1(new_n973), .C2(new_n891), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n991), .A2(new_n996), .A3(new_n997), .ZN(G63));
  XNOR2_X1  g812(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G217), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT60), .Z(new_n1002));
  NAND2_X1  g816(.A1(new_n964), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n251), .A2(new_n242), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n949), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n664), .A2(new_n666), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1000), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n948), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1010), .B(new_n999), .C1(new_n1007), .C2(new_n1003), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(G66));
  AOI21_X1  g826(.A(new_n238), .B1(new_n607), .B2(G224), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n823), .A2(new_n852), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1013), .B1(new_n1014), .B2(new_n238), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n952), .B1(G898), .B2(new_n238), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1015), .B(new_n1016), .Z(G69));
  NOR2_X1   g831(.A1(new_n359), .A2(new_n360), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n457), .A2(new_n459), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n811), .A2(new_n819), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n799), .A2(new_n750), .A3(new_n918), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n840), .A2(new_n682), .A3(new_n705), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1022), .A2(new_n853), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n238), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n678), .A2(G953), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1020), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1023), .A2(new_n698), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT62), .Z(new_n1032));
  NOR2_X1   g846(.A1(new_n685), .A2(new_n802), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n848), .A2(new_n849), .A3(new_n378), .A4(new_n1033), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1032), .A2(new_n811), .A3(new_n819), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1020), .A2(G953), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(G227), .A2(G900), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(G953), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1030), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(KEYINPUT127), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1044), .A2(G953), .A3(new_n1038), .A4(new_n1020), .ZN(new_n1045));
  AND2_X1   g859(.A1(new_n1040), .A2(new_n1045), .ZN(G72));
  NAND2_X1  g860(.A1(new_n859), .A2(new_n865), .ZN(new_n1047));
  NAND2_X1  g861(.A1(G472), .A2(G902), .ZN(new_n1048));
  XOR2_X1   g862(.A(new_n1048), .B(KEYINPUT63), .Z(new_n1049));
  INV_X1    g863(.A(new_n352), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1049), .B1(new_n1050), .B2(new_n691), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n949), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1049), .B1(new_n1035), .B2(new_n1014), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1053), .B1(new_n351), .B2(new_n350), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1049), .B1(new_n1055), .B2(new_n1014), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1056), .A2(new_n342), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1052), .B1(new_n1058), .B2(new_n352), .ZN(G57));
endmodule


