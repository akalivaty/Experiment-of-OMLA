//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  XOR2_X1   g000(.A(G110), .B(G140), .Z(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT10), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(G143), .B2(new_n193), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n196), .A3(new_n198), .A4(G128), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n207), .A2(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n204), .A2(G107), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n192), .B1(new_n203), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT76), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n201), .A2(new_n202), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT76), .A3(new_n192), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT65), .A2(G128), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT65), .A2(G128), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n197), .B1(new_n226), .B2(new_n199), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n202), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n211), .A2(new_n214), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n211), .B2(new_n214), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT10), .B(new_n228), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n205), .A2(new_n208), .A3(new_n210), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT75), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n211), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n197), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n197), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n234), .B(G101), .C1(KEYINPUT75), .C2(new_n236), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n238), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n233), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(KEYINPUT64), .A3(KEYINPUT11), .A4(G134), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(G137), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(new_n251), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n252), .A2(new_n253), .B1(new_n248), .B2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G131), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n258), .A2(new_n259), .A3(new_n249), .A4(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n223), .A2(new_n246), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n223), .B2(new_n246), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n191), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT79), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT79), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n191), .C1(new_n263), .C2(new_n264), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n221), .B1(new_n228), .B2(new_n219), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n261), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n223), .A2(new_n246), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n272), .B(new_n190), .C1(new_n261), .C2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G469), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT69), .B(G902), .Z(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n272), .B(new_n283), .C1(new_n261), .C2(new_n273), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n270), .B(KEYINPUT12), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT78), .B1(new_n285), .B2(new_n263), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n286), .A3(new_n191), .ZN(new_n287));
  OR3_X1    g101(.A1(new_n263), .A2(new_n264), .A3(new_n191), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(G469), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(KEYINPUT9), .B(G234), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G221), .B1(new_n292), .B2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G475), .A2(G902), .ZN(new_n296));
  XNOR2_X1  g110(.A(G113), .B(G122), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n204), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G125), .B(G140), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G146), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n193), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(G143), .A3(G214), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(G143), .B1(new_n305), .B2(G214), .ZN(new_n308));
  OAI21_X1  g122(.A(G131), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT18), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(G214), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n195), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(new_n306), .C1(new_n310), .C2(new_n259), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n314), .A2(KEYINPUT86), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(KEYINPUT86), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n311), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n259), .A3(new_n306), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n301), .A2(KEYINPUT19), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT19), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n300), .A2(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n320), .A2(new_n322), .A3(G146), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT72), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n327), .A3(new_n331), .A4(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n193), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n319), .A2(new_n323), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n299), .B1(new_n317), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n315), .A2(new_n316), .ZN(new_n336));
  INV_X1    g150(.A(new_n311), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT17), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n309), .A2(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT72), .B1(new_n325), .B2(KEYINPUT16), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n193), .B(new_n332), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n332), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G146), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n309), .A2(new_n339), .A3(new_n318), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n340), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n338), .A2(new_n298), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT87), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n335), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n335), .B2(new_n348), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT20), .B(new_n296), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n335), .ZN(new_n353));
  INV_X1    g167(.A(new_n348), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n296), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n298), .B1(new_n338), .B2(new_n347), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n280), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G475), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n352), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT65), .A2(G128), .ZN(new_n362));
  NOR2_X1   g176(.A1(KEYINPUT65), .A2(G128), .ZN(new_n363));
  OAI21_X1  g177(.A(G143), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n195), .A2(G128), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT13), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n368), .A3(G134), .ZN(new_n369));
  XOR2_X1   g183(.A(G116), .B(G122), .Z(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  XNOR2_X1  g185(.A(G116), .B(G122), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n207), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n364), .B(new_n365), .C1(new_n367), .C2(new_n248), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G116), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT14), .A3(G122), .ZN(new_n378));
  OAI211_X1 g192(.A(G107), .B(new_n378), .C1(new_n370), .C2(KEYINPUT14), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n364), .A2(new_n248), .A3(new_n365), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n248), .B1(new_n364), .B2(new_n365), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n379), .B(new_n373), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT88), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT88), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n376), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G217), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n292), .A2(new_n388), .A3(G953), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(new_n389), .A3(new_n386), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n278), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G478), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT15), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n393), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G952), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G953), .ZN(new_n399));
  INV_X1    g213(.A(G234), .ZN(new_n400));
  INV_X1    g214(.A(G237), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n277), .B(G953), .C1(new_n400), .C2(new_n401), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT21), .B(G898), .Z(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n405), .B(KEYINPUT89), .Z(new_n406));
  AND3_X1   g220(.A1(new_n361), .A2(new_n397), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n194), .A2(new_n196), .A3(G128), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n224), .A3(new_n225), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n198), .A2(new_n410), .B1(new_n412), .B2(new_n197), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G125), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(G125), .B2(new_n243), .ZN(new_n415));
  INV_X1    g229(.A(G224), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G953), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(G110), .B(G122), .Z(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n377), .A2(G119), .ZN(new_n422));
  INV_X1    g236(.A(G119), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT66), .B1(new_n423), .B2(G116), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT66), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n377), .A3(G119), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n422), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT2), .B(G113), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n427), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n238), .A3(new_n244), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT5), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n432), .B(new_n422), .C1(new_n426), .C2(new_n424), .ZN(new_n433));
  INV_X1    g247(.A(G113), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n422), .B2(new_n432), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT80), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n427), .A2(new_n429), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n427), .A2(KEYINPUT5), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n435), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n231), .A2(new_n232), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n421), .B(new_n431), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n215), .A2(KEYINPUT77), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n230), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n448), .A2(new_n438), .A3(new_n437), .A4(new_n441), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n449), .A2(KEYINPUT82), .A3(new_n421), .A4(new_n431), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n431), .B1(new_n442), .B2(new_n443), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(KEYINPUT81), .A3(new_n431), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n421), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT6), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n449), .A2(KEYINPUT81), .A3(new_n431), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT81), .B1(new_n449), .B2(new_n431), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n420), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n419), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n415), .B1(new_n464), .B2(new_n417), .ZN(new_n465));
  INV_X1    g279(.A(new_n417), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT7), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n415), .A2(new_n464), .A3(KEYINPUT7), .A4(new_n466), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n468), .A2(new_n469), .B1(new_n446), .B2(new_n450), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n433), .B(KEYINPUT83), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n438), .B1(new_n471), .B2(new_n436), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n219), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n420), .B(KEYINPUT8), .Z(new_n474));
  OAI211_X1 g288(.A(new_n473), .B(new_n474), .C1(new_n219), .C2(new_n442), .ZN(new_n475));
  AOI21_X1  g289(.A(G902), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n409), .B1(new_n463), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n446), .A2(new_n450), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n461), .B1(new_n460), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n418), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n408), .A3(new_n476), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT85), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n487));
  INV_X1    g301(.A(new_n485), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n487), .B(new_n488), .C1(new_n478), .C2(new_n483), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n295), .B(new_n407), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n255), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n248), .A2(G137), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n260), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n413), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n257), .A2(new_n260), .B1(new_n240), .B2(new_n242), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT30), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n261), .A2(new_n243), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n228), .A2(new_n260), .A3(new_n495), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n430), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n427), .B(new_n428), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n506), .A3(new_n502), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n508));
  NAND2_X1  g322(.A1(new_n305), .A2(G210), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G101), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n497), .A2(new_n498), .A3(new_n430), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n504), .B2(new_n430), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT31), .A3(new_n513), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n430), .B1(new_n497), .B2(new_n498), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n520), .B1(new_n521), .B2(new_n507), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n497), .A2(new_n498), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT28), .B1(new_n523), .B2(new_n506), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT68), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n506), .B1(new_n500), .B2(new_n502), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT28), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n516), .A2(new_n519), .B1(new_n530), .B2(new_n512), .ZN(new_n531));
  NOR2_X1   g345(.A1(G472), .A2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT32), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n507), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT68), .B1(new_n535), .B2(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n507), .A2(new_n520), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n527), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n538), .B2(KEYINPUT68), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT31), .B1(new_n518), .B2(new_n513), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n506), .B1(new_n499), .B2(new_n503), .ZN(new_n541));
  NOR4_X1   g355(.A1(new_n541), .A2(new_n515), .A3(new_n517), .A4(new_n512), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n539), .A2(new_n513), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n532), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n505), .A2(new_n507), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n512), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n547), .B(new_n549), .C1(new_n530), .C2(new_n512), .ZN(new_n550));
  INV_X1    g364(.A(new_n538), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n512), .A2(new_n547), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n277), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT70), .B1(new_n554), .B2(G472), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  AOI211_X1 g371(.A(new_n556), .B(new_n557), .C1(new_n550), .C2(new_n553), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n546), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n226), .A2(KEYINPUT71), .A3(G119), .ZN(new_n561));
  OAI21_X1  g375(.A(G119), .B1(new_n362), .B2(new_n363), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n423), .A2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT71), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT23), .B(G119), .C1(new_n362), .C2(new_n363), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n423), .B2(G128), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n563), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G110), .ZN(new_n572));
  INV_X1    g386(.A(new_n343), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n567), .B(new_n572), .C1(new_n573), .C2(new_n333), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(G110), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n566), .B1(new_n561), .B2(new_n565), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n345), .B(new_n303), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT22), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G137), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT73), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n574), .A2(new_n577), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n574), .B2(new_n577), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n581), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n560), .B(KEYINPUT25), .C1(new_n589), .C2(new_n277), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n574), .A2(new_n577), .A3(new_n584), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n588), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n277), .B1(new_n594), .B2(new_n582), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n591), .B1(new_n595), .B2(KEYINPUT74), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n388), .B1(new_n278), .B2(G234), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n590), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n589), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n559), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n482), .A2(new_n408), .A3(new_n476), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n408), .B1(new_n482), .B2(new_n476), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n485), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n487), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n484), .A2(KEYINPUT85), .A3(new_n485), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(KEYINPUT90), .A3(new_n295), .A4(new_n407), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n492), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT91), .B(G101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  NOR2_X1   g429(.A1(new_n531), .A2(new_n277), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n557), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n531), .A2(new_n533), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n620), .A2(new_n294), .A3(new_n602), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n478), .A2(KEYINPUT92), .A3(new_n483), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n607), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n622), .A2(new_n485), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n393), .A2(new_n394), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n391), .A2(new_n627), .A3(new_n392), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n391), .A2(new_n627), .A3(KEYINPUT33), .A4(new_n392), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n277), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n626), .B1(new_n632), .B2(G478), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n361), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT94), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT94), .B1(new_n633), .B2(new_n361), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(new_n406), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n621), .A2(new_n625), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT34), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n204), .ZN(G6));
  AND2_X1   g455(.A1(new_n352), .A2(new_n360), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n406), .B(KEYINPUT95), .Z(new_n643));
  OAI21_X1  g457(.A(new_n296), .B1(new_n350), .B2(new_n351), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n356), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n642), .A2(new_n396), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT96), .Z(new_n647));
  NAND3_X1  g461(.A1(new_n621), .A2(new_n625), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n588), .A2(KEYINPUT36), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n587), .B(new_n652), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n600), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n598), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n619), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n651), .B1(new_n619), .B2(new_n655), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n492), .A2(new_n612), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G12));
  AND4_X1   g476(.A1(new_n559), .A2(new_n293), .A3(new_n290), .A4(new_n655), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n402), .B1(new_n403), .B2(G900), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT99), .Z(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n642), .A2(new_n396), .A3(new_n645), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT100), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n663), .A2(new_n625), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XNOR2_X1  g484(.A(new_n665), .B(KEYINPUT102), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n295), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n295), .A2(KEYINPUT40), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT38), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n606), .A2(new_n607), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n484), .A2(KEYINPUT101), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n484), .A2(KEYINPUT101), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(KEYINPUT38), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n655), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n361), .A2(new_n397), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n548), .A2(new_n513), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n535), .A2(new_n513), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(G902), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n557), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n534), .B2(new_n545), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n677), .A2(new_n687), .A3(new_n485), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  AOI21_X1  g511(.A(new_n488), .B1(new_n679), .B2(KEYINPUT92), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n633), .A2(new_n361), .A3(new_n665), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n698), .A2(new_n699), .A3(new_n624), .A4(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n622), .A3(new_n485), .A4(new_n624), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT103), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n663), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  INV_X1    g519(.A(new_n279), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n276), .B1(new_n275), .B2(new_n278), .ZN(new_n707));
  INV_X1    g521(.A(new_n293), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n638), .A2(new_n605), .A3(new_n625), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  INV_X1    g526(.A(new_n709), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n622), .A2(new_n485), .A3(new_n624), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n605), .A3(new_n647), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AND2_X1   g531(.A1(new_n559), .A2(new_n655), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n407), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n625), .A2(new_n688), .A3(new_n709), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n598), .A2(KEYINPUT104), .A3(new_n601), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT104), .B1(new_n598), .B2(new_n601), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n540), .A2(new_n542), .B1(new_n551), .B2(new_n513), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n532), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n616), .B2(new_n557), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(new_n643), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n721), .B1(new_n722), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n730), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n714), .A2(new_n689), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT105), .A4(new_n709), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  AOI21_X1  g550(.A(new_n728), .B1(new_n598), .B2(new_n654), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n625), .A2(new_n737), .A3(new_n700), .A4(new_n709), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n602), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n598), .A2(KEYINPUT104), .A3(new_n601), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n534), .A2(KEYINPUT106), .A3(new_n545), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT106), .B1(new_n534), .B2(new_n545), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n555), .A2(new_n558), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n633), .ZN(new_n749));
  INV_X1    g563(.A(new_n361), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n666), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n478), .A2(new_n485), .A3(new_n483), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n294), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n748), .A2(new_n753), .A3(KEYINPUT107), .A4(KEYINPUT42), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n533), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n544), .B1(new_n543), .B2(new_n532), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n534), .A2(KEYINPUT106), .A3(new_n545), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n555), .A2(new_n558), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n725), .B(KEYINPUT42), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n752), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n293), .A3(new_n290), .A4(new_n700), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n755), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n294), .A2(new_n752), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n605), .A2(new_n700), .A3(new_n768), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n754), .A2(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n259), .ZN(G33));
  NOR3_X1   g585(.A1(new_n604), .A2(new_n294), .A3(new_n752), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n668), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  NAND2_X1  g588(.A1(new_n287), .A2(new_n288), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT45), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(G469), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(KEYINPUT108), .A3(G469), .A4(new_n778), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n282), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n281), .B1(new_n781), .B2(new_n782), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n706), .B1(new_n788), .B2(KEYINPUT46), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT109), .B1(new_n788), .B2(KEYINPUT46), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n293), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n750), .A2(new_n633), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n749), .A2(new_n361), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n795), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n620), .A3(new_n655), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(new_n808), .A3(new_n805), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n752), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n804), .A2(new_n805), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n793), .A2(new_n810), .A3(new_n672), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n792), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n791), .A2(new_n293), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n559), .A2(new_n603), .A3(new_n752), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n816), .A2(new_n700), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  AND2_X1   g636(.A1(new_n683), .A2(new_n686), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT49), .B1(new_n706), .B2(new_n707), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n706), .A2(new_n707), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n488), .B(new_n801), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n823), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n293), .A3(new_n694), .A4(new_n725), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  INV_X1    g644(.A(new_n819), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n791), .A2(new_n293), .B1(KEYINPUT112), .B2(new_n814), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT115), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n816), .A2(new_n834), .A3(new_n819), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n825), .A2(new_n708), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n402), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n803), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n725), .A2(new_n729), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n839), .A2(new_n840), .A3(new_n752), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n709), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n823), .A2(new_n488), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n839), .A2(new_n713), .A3(new_n752), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n737), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n713), .A2(new_n602), .A3(new_n752), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n838), .A3(new_n694), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n750), .A3(new_n749), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n849), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n830), .B1(new_n842), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n636), .A2(new_n637), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n850), .A2(new_n748), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n862));
  OAI221_X1 g676(.A(new_n399), .B1(new_n859), .B2(new_n853), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n836), .B1(new_n831), .B2(new_n832), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n830), .B1(new_n864), .B2(new_n841), .ZN(new_n865));
  INV_X1    g679(.A(new_n851), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n866), .B(new_n854), .C1(new_n847), .C2(new_n848), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n863), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n843), .A2(new_n715), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n857), .A2(new_n858), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n856), .B1(new_n837), .B2(new_n841), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n868), .B(new_n869), .C1(new_n871), .C2(KEYINPUT51), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(new_n773), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n642), .A2(new_n645), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n559), .A2(new_n397), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n634), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n877), .B1(new_n878), .B2(new_n728), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n655), .A2(new_n879), .A3(new_n666), .A4(new_n768), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n770), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n621), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n634), .B(new_n643), .C1(new_n486), .C2(new_n489), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT113), .ZN(new_n884));
  INV_X1    g698(.A(new_n643), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n609), .B2(new_n610), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT113), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n634), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n882), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n642), .A2(new_n357), .A3(new_n396), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n710), .B1(new_n891), .B2(new_n882), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n716), .A2(new_n719), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n492), .B(new_n612), .C1(new_n605), .C2(new_n658), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(new_n735), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n881), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n694), .A2(new_n655), .A3(new_n665), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n733), .A2(new_n295), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n704), .A2(new_n669), .A3(new_n738), .A4(new_n899), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT52), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(KEYINPUT53), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT52), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n900), .A2(new_n905), .A3(KEYINPUT52), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n881), .A2(new_n894), .A3(new_n896), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n874), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n904), .B1(new_n910), .B2(new_n901), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n900), .A2(new_n905), .A3(KEYINPUT52), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n906), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n883), .A2(KEYINPUT113), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n887), .B1(new_n886), .B2(new_n634), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n621), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n709), .A2(new_n485), .A3(new_n624), .A4(new_n622), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n636), .A2(new_n406), .A3(new_n637), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n604), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n886), .A2(new_n890), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n621), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n716), .A2(new_n719), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n895), .A2(new_n735), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n915), .A2(new_n927), .A3(KEYINPUT53), .A4(new_n881), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n913), .A2(new_n928), .A3(new_n874), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n912), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n870), .A2(new_n873), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n398), .A2(new_n188), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT117), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n829), .B1(new_n931), .B2(new_n933), .ZN(G75));
  AOI21_X1  g748(.A(new_n278), .B1(new_n913), .B2(new_n928), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(new_n409), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n480), .A2(new_n481), .A3(new_n418), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n463), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n936), .A2(new_n939), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n398), .A2(G953), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT118), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(G51));
  INV_X1    g759(.A(KEYINPUT119), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n281), .B(KEYINPUT57), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n913), .A2(new_n928), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT54), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n913), .A2(new_n928), .A3(new_n874), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n275), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n935), .A2(new_n781), .A3(new_n782), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n874), .B1(new_n913), .B2(new_n928), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n947), .B1(new_n929), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(KEYINPUT119), .A3(new_n275), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n943), .ZN(G54));
  NAND3_X1  g774(.A1(new_n935), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n350), .A2(new_n351), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n963), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n943), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n964), .A2(KEYINPUT120), .A3(new_n943), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G60));
  NAND2_X1  g784(.A1(new_n630), .A2(new_n631), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT59), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n929), .B2(new_n956), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(KEYINPUT121), .B(new_n975), .C1(new_n929), .C2(new_n956), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT53), .B1(new_n897), .B2(new_n915), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n910), .A2(new_n904), .A3(new_n901), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT54), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n974), .B1(new_n983), .B2(new_n951), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n943), .B1(new_n984), .B2(new_n971), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT122), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n974), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n912), .B2(new_n929), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n944), .B1(new_n988), .B2(new_n972), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(new_n990), .A3(new_n978), .A4(new_n979), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n986), .A2(new_n991), .ZN(G63));
  XNOR2_X1  g806(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n388), .A2(new_n280), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n949), .A2(new_n653), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n949), .A2(new_n995), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n943), .B(new_n996), .C1(new_n997), .C2(new_n599), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT123), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT61), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(KEYINPUT61), .B1(new_n998), .B2(new_n999), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(G66));
  INV_X1    g817(.A(new_n404), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n1004), .B2(new_n416), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n927), .B2(G953), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n457), .B(new_n462), .C1(G898), .C2(new_n188), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G69));
  AND2_X1   g822(.A1(new_n669), .A2(new_n738), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1009), .A2(new_n704), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(KEYINPUT62), .A3(new_n696), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1012));
  INV_X1    g826(.A(new_n696), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1009), .A2(new_n704), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n772), .B(new_n672), .C1(new_n634), .C2(new_n890), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1016), .A2(new_n812), .A3(new_n821), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n188), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n320), .A2(new_n322), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n504), .B(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(KEYINPUT125), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n821), .A2(new_n812), .A3(new_n1010), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n770), .A2(new_n875), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n793), .A2(new_n672), .A3(new_n733), .A4(new_n748), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1024), .A2(new_n188), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1021), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G900), .A2(G953), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT125), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1019), .A2(new_n1031), .A3(new_n1021), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1023), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT126), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OR2_X1    g850(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1033), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1036), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  AND4_X1   g854(.A1(new_n927), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1041));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  OAI211_X1 g858(.A(new_n518), .B(new_n512), .C1(new_n1041), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n927), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1043), .B1(new_n1018), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(new_n690), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n944), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1044), .B1(new_n549), .B2(new_n514), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT127), .Z(new_n1051));
  OAI21_X1  g865(.A(new_n1051), .B1(new_n981), .B2(new_n982), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n1045), .A2(new_n1049), .A3(new_n1052), .ZN(G57));
endmodule


