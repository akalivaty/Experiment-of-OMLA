//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  OR2_X1    g031(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  AOI21_X1  g033(.A(G2105), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G137), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n459), .A2(new_n462), .A3(G137), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n461), .A2(KEYINPUT66), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n457), .A2(new_n458), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n464), .B1(new_n457), .B2(new_n458), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NAND2_X1  g053(.A1(G112), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G100), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT68), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n459), .A2(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n459), .A2(KEYINPUT67), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n478), .B(new_n483), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT69), .ZN(G162));
  NAND2_X1  g064(.A1(new_n459), .A2(G138), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n457), .B2(new_n458), .ZN(new_n494));
  AND2_X1   g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n457), .B2(new_n458), .ZN(new_n498));
  AND2_X1   g073(.A1(G102), .A2(G2104), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n464), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n492), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n504));
  OAI211_X1 g079(.A(KEYINPUT72), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT70), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT70), .A2(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT5), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT72), .B1(new_n510), .B2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT73), .A3(G62), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n503), .B2(new_n504), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(new_n505), .A3(new_n508), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(G75), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n513), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n517), .A2(new_n505), .A3(new_n508), .A4(new_n525), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT74), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  AOI211_X1 g109(.A(new_n534), .B(new_n531), .C1(new_n523), .C2(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  AND2_X1   g112(.A1(new_n505), .A2(new_n508), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n538), .A2(G63), .A3(G651), .A4(new_n517), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n527), .A2(G51), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT75), .B(G89), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n539), .B(new_n543), .C1(new_n529), .C2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n527), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n529), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n517), .A2(G64), .A3(new_n505), .A4(new_n508), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n549), .A2(new_n553), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n518), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n527), .A2(G43), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n560), .C1(new_n529), .C2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n538), .A2(G81), .A3(new_n517), .A4(new_n525), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n559), .B1(new_n564), .B2(new_n560), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n558), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  NAND3_X1  g148(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  AND4_X1   g150(.A1(new_n517), .A2(new_n505), .A3(new_n508), .A4(new_n525), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G91), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n517), .A2(G65), .A3(new_n505), .A4(new_n508), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n575), .B(new_n577), .C1(new_n580), .C2(new_n550), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  NAND2_X1  g157(.A1(new_n527), .A2(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n529), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n550), .B1(new_n518), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G288));
  NAND4_X1  g164(.A1(new_n517), .A2(G61), .A3(new_n505), .A4(new_n508), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(KEYINPUT77), .B1(new_n592), .B2(G651), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  AOI211_X1 g169(.A(new_n594), .B(new_n550), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n529), .ZN(new_n600));
  NOR3_X1   g175(.A1(new_n593), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n527), .A2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n576), .A2(G85), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n550), .ZN(G290));
  NAND4_X1  g181(.A1(new_n517), .A2(G66), .A3(new_n505), .A4(new_n508), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n527), .A2(G54), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n512), .A2(G92), .A3(new_n525), .A4(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n612), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n529), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n610), .A2(new_n611), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  MUX2_X1   g192(.A(new_n617), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g193(.A(new_n617), .B(G301), .S(G868), .Z(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g196(.A(new_n620), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(new_n617), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NOR2_X1   g200(.A1(new_n566), .A2(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n617), .A2(G559), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n626), .B1(G868), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n459), .A2(G2104), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2100), .ZN(new_n635));
  MUX2_X1   g210(.A(G99), .B(G111), .S(G2105), .Z(new_n636));
  AOI22_X1  g211(.A1(G123), .A2(new_n477), .B1(new_n636), .B2(G2104), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n486), .B2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n635), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2427), .ZN(new_n646));
  INV_X1    g221(.A(G2430), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2084), .B(G2090), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(KEYINPUT17), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n663), .B2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT80), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n666), .A2(new_n659), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n660), .A2(new_n659), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n665), .B(new_n668), .C1(new_n663), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n640), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT81), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n674), .A2(new_n676), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n683), .A2(new_n679), .A3(new_n677), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n684), .C1(new_n679), .C2(new_n683), .ZN(new_n685));
  XOR2_X1   g260(.A(G1981), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT82), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n687), .B(new_n691), .ZN(G229));
  NAND2_X1  g267(.A1(G162), .A2(G29), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G29), .B2(G35), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT29), .ZN(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G32), .ZN(new_n699));
  INV_X1    g274(.A(new_n486), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(G141), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT93), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n477), .A2(G129), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND3_X1  g281(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n699), .B1(new_n708), .B2(new_n698), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G27), .A2(G29), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G164), .B2(G29), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT94), .B(G2078), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n709), .A2(new_n711), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n712), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G21), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G168), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G1966), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n714), .A2(new_n715), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n698), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n639), .B2(new_n698), .ZN(new_n729));
  NOR4_X1   g304(.A1(new_n718), .A2(new_n724), .A3(new_n725), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n697), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n695), .A2(new_n696), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n719), .A2(G19), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT86), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n567), .B2(new_n719), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1341), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n698), .A2(G33), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(new_n464), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT89), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n700), .A2(G139), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n742));
  NAND3_X1  g317(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT90), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n737), .B1(new_n746), .B2(new_n698), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2072), .ZN(new_n748));
  NOR4_X1   g323(.A1(new_n731), .A2(new_n732), .A3(new_n736), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT95), .B(KEYINPUT23), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n719), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n698), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  MUX2_X1   g333(.A(G104), .B(G116), .S(G2105), .Z(new_n759));
  AOI22_X1  g334(.A1(G128), .A2(new_n477), .B1(new_n759), .B2(G2104), .ZN(new_n760));
  INV_X1    g335(.A(G140), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n486), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT87), .Z(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(new_n763), .B2(new_n698), .ZN(new_n764));
  INV_X1    g339(.A(G2067), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G171), .A2(new_n719), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G5), .B2(new_n719), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n766), .B1(G1961), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(KEYINPUT24), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(KEYINPUT24), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(KEYINPUT91), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(KEYINPUT91), .B2(new_n773), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n475), .B2(new_n698), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2084), .ZN(new_n778));
  NOR2_X1   g353(.A1(G4), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n623), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1348), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n768), .A2(new_n782), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n770), .A2(new_n778), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n749), .A2(new_n756), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n749), .A2(KEYINPUT97), .A3(new_n756), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G6), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n601), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT84), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT32), .B(G1981), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n719), .A2(G23), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n588), .B2(new_n719), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n794), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n719), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n719), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT85), .B(G1971), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n800), .A2(new_n804), .A3(KEYINPUT34), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT34), .B1(new_n800), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g381(.A1(G25), .A2(G29), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n700), .A2(G131), .ZN(new_n808));
  MUX2_X1   g383(.A(G95), .B(G107), .S(G2105), .Z(new_n809));
  AOI22_X1  g384(.A1(G119), .A2(new_n477), .B1(new_n809), .B2(G2104), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(G29), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NAND2_X1  g390(.A1(G290), .A2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1986), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n719), .A2(G24), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT83), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n816), .B2(new_n819), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n815), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n805), .A2(new_n806), .A3(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n789), .A2(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n789), .A2(new_n826), .ZN(G150));
  NAND4_X1  g403(.A1(new_n517), .A2(G67), .A3(new_n505), .A4(new_n508), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n829), .A2(KEYINPUT98), .A3(new_n830), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(G651), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n576), .A2(G93), .B1(G55), .B2(new_n527), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT99), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n566), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n560), .B1(new_n529), .B2(new_n561), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT76), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n562), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n558), .A2(new_n844), .B1(new_n835), .B2(new_n836), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n617), .A2(new_n624), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n850), .B2(KEYINPUT39), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n840), .B1(new_n851), .B2(new_n853), .ZN(G145));
  XNOR2_X1  g429(.A(G162), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n639), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n763), .A2(G164), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n762), .B(KEYINPUT87), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n501), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n708), .ZN(new_n861));
  INV_X1    g436(.A(new_n708), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n862), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n746), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n745), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n867), .A3(new_n863), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n811), .B(new_n631), .ZN(new_n870));
  MUX2_X1   g445(.A(G106), .B(G118), .S(G2105), .Z(new_n871));
  AOI22_X1  g446(.A1(G130), .A2(new_n477), .B1(new_n871), .B2(G2104), .ZN(new_n872));
  INV_X1    g447(.A(G142), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n486), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT100), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n869), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n866), .A2(KEYINPUT100), .A3(new_n868), .A4(new_n875), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n856), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(G37), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n856), .A3(new_n879), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(KEYINPUT101), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(KEYINPUT101), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g461(.A1(new_n837), .A2(G868), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n524), .A2(new_n532), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n534), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n524), .A2(KEYINPUT74), .A3(new_n532), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(G305), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n601), .B1(new_n533), .B2(new_n535), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n585), .B2(new_n587), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n576), .A2(G87), .ZN(new_n895));
  OAI21_X1  g470(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT105), .A4(new_n583), .ZN(new_n897));
  AND3_X1   g472(.A1(G290), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G290), .B1(new_n894), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n891), .A2(new_n892), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n891), .B2(new_n892), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT42), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT107), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT106), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n891), .A2(new_n892), .ZN(new_n906));
  INV_X1    g481(.A(new_n900), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n891), .A2(new_n892), .A3(new_n900), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n904), .B1(KEYINPUT42), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n846), .B(new_n627), .Z(new_n914));
  AOI21_X1  g489(.A(new_n550), .B1(new_n578), .B2(new_n579), .ZN(new_n915));
  INV_X1    g490(.A(G91), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n529), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT9), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n574), .B(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n613), .A2(new_n616), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n617), .A2(G299), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT103), .A4(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT41), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n914), .A2(KEYINPUT104), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT102), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n933), .B1(new_n914), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT104), .B1(new_n914), .B2(new_n932), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n913), .B(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n887), .B1(new_n942), .B2(G868), .ZN(G295));
  AOI21_X1  g518(.A(new_n887), .B1(new_n942), .B2(G868), .ZN(G331));
  NAND2_X1  g519(.A1(G168), .A2(G171), .ZN(new_n945));
  OAI21_X1  g520(.A(G286), .B1(new_n553), .B2(new_n549), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n841), .B2(new_n845), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n837), .A2(new_n566), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n844), .A2(new_n835), .A3(new_n558), .A4(new_n836), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n946), .A4(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(new_n930), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n932), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n932), .B2(new_n952), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n960), .B(new_n954), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n912), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n932), .A2(new_n952), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n932), .A2(new_n952), .A3(new_n955), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n912), .A2(new_n966), .A3(new_n954), .ZN(new_n967));
  INV_X1    g542(.A(G37), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n962), .C2(new_n969), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n931), .A2(new_n926), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n952), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n948), .A2(new_n951), .A3(new_n935), .A4(new_n936), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n978), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n905), .B(new_n911), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n967), .A2(new_n975), .A3(new_n968), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n953), .B1(new_n964), .B2(new_n965), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n986), .B2(new_n912), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(KEYINPUT112), .A3(new_n975), .A4(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n962), .A2(new_n969), .A3(KEYINPUT43), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n975), .B1(new_n987), .B2(new_n982), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(G397));
  NAND4_X1  g569(.A1(new_n474), .A2(G40), .A3(new_n466), .A4(new_n470), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n501), .A2(KEYINPUT116), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT116), .B1(new_n501), .B2(new_n997), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n588), .A2(G1976), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(G8), .A3(new_n1003), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1002), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n601), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n600), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n592), .A2(G651), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n594), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n592), .A2(KEYINPUT77), .A3(G651), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1012), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT118), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n601), .A2(new_n1012), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1010), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1022), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1009), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n889), .A2(G8), .A3(new_n890), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n501), .A2(new_n997), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n501), .A2(KEYINPUT116), .A3(new_n997), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT50), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n996), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1033), .B1(new_n1041), .B2(G2090), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1034), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT115), .A3(new_n996), .ZN(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(new_n995), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1039), .B1(new_n998), .B2(new_n999), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1040), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n995), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(KEYINPUT117), .A3(new_n696), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1042), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1032), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1027), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(G8), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1043), .B1(new_n998), .B2(new_n999), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1045), .A2(KEYINPUT119), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1045), .A2(KEYINPUT119), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1063), .A2(new_n996), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n722), .ZN(new_n1067));
  INV_X1    g642(.A(G2084), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1055), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G8), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G286), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1059), .A2(KEYINPUT63), .A3(new_n1062), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1036), .A2(KEYINPUT50), .A3(new_n1037), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n996), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1052), .B1(G2090), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1061), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1027), .A2(new_n1080), .A3(new_n1058), .A4(new_n1072), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT120), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1081), .A2(KEYINPUT120), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1073), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(new_n1004), .A3(new_n588), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1010), .B1(new_n1088), .B2(new_n1020), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1058), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1027), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1041), .A2(new_n782), .ZN(new_n1092));
  INV_X1    g667(.A(G2078), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(KEYINPUT53), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n1066), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n1097), .B2(new_n1093), .ZN(new_n1098));
  OAI21_X1  g673(.A(G171), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(G286), .A2(G8), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT51), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1071), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1102), .C1(new_n1070), .C2(G286), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1070), .A2(G8), .A3(G286), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1104), .A2(KEYINPUT62), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1099), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  INV_X1    g687(.A(G1348), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1041), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n996), .A2(new_n1000), .A3(new_n765), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1112), .B(new_n1115), .C1(new_n1055), .C2(G1348), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1050), .A2(new_n995), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT56), .B(G2072), .Z(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1077), .A2(new_n755), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1124), .B(new_n577), .C1(new_n580), .C2(new_n550), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT121), .B1(new_n915), .B2(new_n917), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n575), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n1128), .B2(G299), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1123), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1119), .A2(new_n623), .A3(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1136), .A2(KEYINPUT122), .B1(KEYINPUT57), .B2(new_n920), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n995), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1046), .A2(new_n996), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1138), .A2(G1956), .B1(new_n1139), .B2(new_n1121), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1132), .A3(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1116), .A2(new_n1118), .A3(KEYINPUT60), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT60), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n623), .ZN(new_n1145));
  OAI211_X1 g720(.A(KEYINPUT60), .B(new_n617), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1134), .A2(new_n1141), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1134), .A2(new_n1141), .A3(KEYINPUT61), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1139), .A2(G1996), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT58), .B(G1341), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n996), .B2(new_n1000), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n567), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT59), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1150), .A2(new_n1151), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1142), .B1(new_n1147), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1095), .B(new_n1050), .C1(KEYINPUT125), .C2(new_n996), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(KEYINPUT125), .B2(new_n996), .ZN(new_n1160));
  XOR2_X1   g735(.A(G171), .B(KEYINPUT54), .Z(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1092), .A3(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(new_n1098), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1161), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1107), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1111), .B1(new_n1158), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1059), .A2(new_n1080), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1086), .B(new_n1091), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n858), .B(G2067), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n995), .A2(new_n1044), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1172), .A2(KEYINPUT113), .ZN(new_n1173));
  INV_X1    g748(.A(G1996), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n708), .B(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1171), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1172), .B2(KEYINPUT113), .ZN(new_n1177));
  OR3_X1    g752(.A1(new_n1173), .A2(new_n1177), .A3(KEYINPUT114), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT114), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n811), .B(new_n814), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1171), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(G1986), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(new_n1171), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1169), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1171), .B1(new_n1170), .B2(new_n862), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT46), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1188));
  NOR4_X1   g763(.A1(new_n995), .A2(new_n1044), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT47), .ZN(new_n1191));
  NOR2_X1   g766(.A1(G290), .A2(G1986), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1171), .A2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT48), .Z(new_n1194));
  OAI21_X1  g769(.A(new_n1191), .B1(new_n1182), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n812), .A2(new_n814), .ZN(new_n1197));
  OAI22_X1  g772(.A1(new_n1196), .A2(new_n1197), .B1(G2067), .B2(new_n858), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n1198), .B2(new_n1171), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1185), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(G319), .ZN(new_n1202));
  OR2_X1    g776(.A1(G227), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OR2_X1    g779(.A1(G229), .A2(G401), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1207));
  NOR3_X1   g781(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n885), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n989), .A2(new_n974), .ZN(new_n1210));
  INV_X1    g784(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1209), .B1(new_n972), .B2(new_n1211), .ZN(G308));
  INV_X1    g786(.A(new_n972), .ZN(new_n1213));
  OAI211_X1 g787(.A(new_n885), .B(new_n1208), .C1(new_n1213), .C2(new_n1210), .ZN(G225));
endmodule


