//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G143), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n189), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n190), .A2(new_n192), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n194), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n197), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n193), .A2(G128), .A3(new_n210), .A4(new_n196), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT69), .B(G128), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n193), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n211), .B1(new_n214), .B2(new_n202), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n207), .B1(G125), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G224), .ZN(new_n218));
  XOR2_X1   g032(.A(new_n218), .B(KEYINPUT80), .Z(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT81), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n216), .B(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(G107), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n226), .A2(new_n224), .A3(G107), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n228), .A2(G104), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  OAI22_X1  g045(.A1(new_n228), .A2(G104), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n226), .B1(new_n224), .B2(G107), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n228), .A2(KEYINPUT77), .A3(KEYINPUT3), .A4(G104), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n237), .A3(KEYINPUT4), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n230), .A2(new_n239), .A3(G101), .ZN(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT70), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT2), .B(G113), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n245), .A2(new_n249), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n238), .A2(new_n240), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n228), .A2(G104), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n224), .A2(G107), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n236), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n235), .B2(new_n236), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n246), .B2(new_n248), .ZN(new_n259));
  OAI21_X1  g073(.A(G113), .B1(new_n242), .B2(KEYINPUT5), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n257), .B(new_n251), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n253), .A2(KEYINPUT79), .A3(new_n261), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G122), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n253), .A2(new_n261), .A3(new_n266), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n262), .B2(new_n263), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT6), .B1(new_n271), .B2(new_n265), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n221), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT7), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n219), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n216), .B(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n266), .B(KEYINPUT8), .Z(new_n277));
  NOR2_X1   g091(.A1(new_n245), .A2(new_n258), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n251), .B1(new_n278), .B2(new_n260), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n257), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n251), .B1(new_n259), .B2(new_n260), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n257), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n269), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n273), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT82), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n273), .A2(new_n284), .A3(new_n286), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n188), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT9), .B(G234), .ZN(new_n291));
  INV_X1    g105(.A(G217), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n291), .A2(new_n292), .A3(G953), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G122), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G116), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n243), .A2(G122), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(G107), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n212), .A2(G143), .ZN(new_n300));
  INV_X1    g114(.A(G134), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n201), .A2(G128), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n201), .A2(KEYINPUT13), .A3(G128), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT13), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n212), .A2(G143), .B1(new_n308), .B2(new_n302), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n301), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n296), .A2(KEYINPUT14), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n298), .A2(new_n312), .A3(G107), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n296), .B(new_n297), .C1(KEYINPUT14), .C2(new_n228), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n300), .A2(new_n302), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G134), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n317), .B2(new_n303), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n294), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n314), .B(new_n313), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n322), .B(new_n293), .C1(new_n310), .C2(new_n304), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT89), .ZN(new_n326));
  INV_X1    g140(.A(G902), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT87), .B(new_n294), .C1(new_n311), .C2(new_n318), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G478), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n329), .B(KEYINPUT88), .C1(KEYINPUT15), .C2(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n329), .A2(KEYINPUT88), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(KEYINPUT15), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(KEYINPUT88), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n331), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n217), .A2(G952), .ZN(new_n337));
  NAND2_X1  g151(.A1(G234), .A2(G237), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT21), .B(G898), .Z(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(G902), .A3(G953), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n343));
  NOR2_X1   g157(.A1(G237), .A2(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G143), .A3(G214), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(G143), .B1(new_n344), .B2(G214), .ZN(new_n347));
  OAI21_X1  g161(.A(G131), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(G214), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n201), .ZN(new_n350));
  INV_X1    g164(.A(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n345), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT17), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G125), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G140), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT16), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n356), .A2(KEYINPUT16), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n189), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G125), .B(G140), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n362), .B2(KEYINPUT16), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G146), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT17), .B(G131), .C1(new_n346), .C2(new_n347), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n354), .A2(new_n361), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n356), .A2(new_n358), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n362), .A2(KEYINPUT74), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT64), .B(G146), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n362), .B2(new_n189), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n367), .A2(KEYINPUT83), .A3(G146), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT18), .A2(G131), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n346), .B2(new_n347), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n350), .A2(KEYINPUT18), .A3(G131), .A4(new_n345), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n366), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n224), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n343), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g200(.A(KEYINPUT85), .B(new_n384), .C1(new_n366), .C2(new_n381), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n382), .A2(new_n385), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n327), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G475), .A2(G902), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n348), .A2(new_n352), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT19), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n369), .A2(new_n370), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n396), .B(new_n371), .C1(new_n395), .C2(new_n362), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT84), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n394), .A2(new_n397), .A3(new_n364), .A4(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n384), .B1(new_n399), .B2(new_n381), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n391), .B1(new_n400), .B2(new_n389), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT20), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n403), .B(new_n391), .C1(new_n400), .C2(new_n389), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n390), .A2(G475), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n336), .A2(new_n342), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n386), .ZN(new_n409));
  INV_X1    g223(.A(new_n387), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n389), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G475), .B1(new_n411), .B2(G902), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n404), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n412), .A2(new_n413), .A3(new_n342), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT90), .B1(new_n414), .B2(new_n336), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n290), .B1(new_n408), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G469), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n195), .B1(new_n371), .B2(G143), .ZN(new_n418));
  INV_X1    g232(.A(G128), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n211), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n257), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n215), .B2(new_n257), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT66), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT11), .A2(G134), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(G137), .ZN(new_n426));
  INV_X1    g240(.A(G137), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n427), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n427), .B2(G134), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n301), .A2(KEYINPUT67), .A3(G137), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(G134), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT11), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n427), .C2(G134), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n429), .B(new_n433), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G131), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n436), .B1(new_n301), .B2(G137), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT65), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n435), .A2(new_n434), .A3(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(new_n351), .A3(new_n429), .A4(new_n433), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n423), .A2(KEYINPUT12), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT12), .B1(new_n423), .B2(new_n446), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT10), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n422), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n198), .B1(new_n371), .B2(G143), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n452), .A2(new_n204), .B1(new_n418), .B2(new_n194), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n238), .A2(new_n240), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n445), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n442), .A2(new_n443), .B1(new_n431), .B2(new_n432), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n351), .B1(new_n456), .B2(new_n429), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n215), .A2(KEYINPUT10), .A3(new_n257), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n451), .A2(new_n454), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G140), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n217), .A2(G227), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n461), .B(new_n462), .Z(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n449), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n451), .A2(new_n454), .A3(new_n459), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n446), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n468), .B2(new_n460), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n417), .B(new_n327), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n460), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n463), .B1(new_n449), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n460), .A2(new_n464), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(G469), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n417), .A2(new_n327), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(KEYINPUT78), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT91), .B1(new_n416), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n292), .B1(G234), .B2(new_n327), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n362), .B(new_n368), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n487), .A2(new_n371), .B1(G146), .B2(new_n363), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n419), .A2(KEYINPUT69), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G128), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n491), .A3(G119), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(G119), .B2(new_n419), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT73), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT24), .B(G110), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n212), .A2(KEYINPUT23), .A3(G119), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT23), .B1(new_n419), .B2(G119), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n241), .B2(G128), .ZN(new_n499));
  INV_X1    g313(.A(G110), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n488), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n364), .A2(new_n361), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n497), .A2(new_n499), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G110), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n493), .A2(new_n495), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT76), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n504), .A2(new_n512), .A3(new_n509), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT75), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(KEYINPUT76), .A3(new_n517), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT25), .B1(new_n521), .B2(new_n327), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n523), .B(G902), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n486), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n486), .A2(G902), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n529));
  INV_X1    g343(.A(new_n435), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n427), .A2(G134), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n215), .A2(new_n445), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n206), .B1(new_n440), .B2(new_n445), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT30), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n453), .B1(new_n455), .B2(new_n457), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n215), .A2(new_n445), .A3(new_n532), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n252), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n252), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n344), .A2(G210), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT27), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(G101), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT31), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n540), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n546), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT28), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n252), .B1(new_n533), .B2(new_n534), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(new_n542), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n533), .A2(new_n534), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT28), .B1(new_n555), .B2(new_n541), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT30), .B1(new_n533), .B2(new_n534), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n537), .A2(new_n536), .A3(new_n538), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n541), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT31), .B1(new_n560), .B2(new_n547), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n550), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT71), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n529), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI211_X1 g381(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n562), .C2(new_n564), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(KEYINPUT32), .A3(new_n564), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G472), .ZN(new_n572));
  OR3_X1    g386(.A1(new_n554), .A2(new_n556), .A3(new_n551), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT29), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n533), .A2(new_n534), .A3(new_n252), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n551), .B1(new_n560), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n554), .A2(new_n556), .A3(new_n551), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n578), .B2(KEYINPUT29), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n572), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n528), .B1(new_n569), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n478), .A2(KEYINPUT78), .A3(new_n479), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT78), .B1(new_n478), .B2(new_n479), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n406), .A2(new_n407), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n414), .A2(KEYINPUT90), .A3(new_n336), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(new_n586), .A3(new_n589), .A4(new_n290), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n485), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  INV_X1    g406(.A(new_n289), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n286), .B1(new_n273), .B2(new_n284), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n187), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n342), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n325), .A2(new_n598), .A3(new_n328), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n319), .A2(new_n323), .A3(KEYINPUT33), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(G478), .A3(new_n327), .A4(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT92), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n334), .A2(new_n602), .A3(new_n330), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n334), .B2(new_n330), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(new_n405), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n597), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n562), .A2(new_n327), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n565), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n528), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n585), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n404), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT94), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n404), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n402), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n402), .A3(new_n622), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n412), .A3(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n597), .A2(new_n336), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n614), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n518), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n510), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n526), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n513), .A2(new_n518), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n512), .B1(new_n504), .B2(new_n509), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n520), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n327), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n523), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n521), .A2(KEYINPUT25), .A3(new_n327), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n635), .B1(new_n643), .B2(new_n486), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n612), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n485), .A2(new_n590), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT95), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  NAND2_X1  g463(.A1(new_n569), .A2(new_n581), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n339), .B1(G900), .B2(new_n341), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n625), .A2(new_n412), .A3(new_n626), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n336), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n595), .A2(new_n644), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n650), .A2(new_n585), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  XNOR2_X1  g470(.A(new_n651), .B(KEYINPUT39), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n585), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n288), .A2(new_n289), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT38), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n525), .A2(new_n634), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n663), .A2(new_n336), .A3(new_n405), .A4(new_n188), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n659), .A2(new_n660), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n546), .B1(new_n553), .B2(new_n542), .ZN(new_n666));
  OAI22_X1  g480(.A1(KEYINPUT96), .A2(new_n666), .B1(new_n560), .B2(new_n547), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(KEYINPUT96), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n327), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G472), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n570), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n565), .A2(new_n566), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT72), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n565), .A2(new_n529), .A3(new_n566), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT97), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n569), .A2(KEYINPUT97), .A3(new_n671), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n665), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT98), .B(G143), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G45));
  NAND2_X1  g497(.A1(new_n412), .A2(new_n413), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n605), .A2(new_n684), .A3(new_n651), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n650), .A2(new_n585), .A3(new_n654), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  OAI21_X1  g501(.A(new_n473), .B1(new_n447), .B2(new_n448), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n468), .A2(new_n460), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n463), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n417), .ZN(new_n692));
  INV_X1    g506(.A(new_n470), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n479), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n528), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n694), .A2(KEYINPUT99), .A3(new_n479), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n650), .A2(new_n697), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n609), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n628), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND2_X1  g519(.A1(new_n697), .A2(new_n699), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n595), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n644), .B1(new_n587), .B2(new_n588), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n650), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n336), .B2(new_n405), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n329), .A2(KEYINPUT88), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n713), .B(new_n333), .C1(KEYINPUT88), .C2(new_n334), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n684), .A2(new_n714), .A3(KEYINPUT100), .A4(new_n331), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n342), .A2(new_n613), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AOI22_X1  g532(.A1(new_n610), .A2(G472), .B1(new_n562), .B2(new_n564), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n685), .A2(new_n663), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n697), .A3(new_n596), .A4(new_n699), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n581), .A2(new_n672), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n698), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n288), .A2(new_n187), .A3(new_n289), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n480), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n685), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT42), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n685), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n582), .A2(new_n731), .A3(new_n727), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n723), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n723), .A3(new_n732), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n351), .ZN(G33));
  NAND3_X1  g551(.A1(new_n582), .A2(new_n653), .A3(new_n727), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  NAND2_X1  g553(.A1(new_n472), .A2(new_n474), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n417), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT102), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n741), .B2(new_n740), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n742), .A2(KEYINPUT102), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n477), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n693), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n747), .B2(new_n746), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n479), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(KEYINPUT103), .A3(new_n657), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n479), .A3(new_n657), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n605), .B(new_n405), .C1(new_n755), .C2(KEYINPUT43), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n606), .A2(new_n684), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n612), .A3(new_n663), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(new_n726), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n751), .A2(new_n754), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(KEYINPUT105), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(KEYINPUT105), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n750), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n650), .A2(new_n730), .A3(new_n698), .A4(new_n726), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n771), .B(new_n772), .C1(new_n750), .C2(new_n770), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  OAI21_X1  g588(.A(new_n771), .B1(new_n750), .B2(new_n770), .ZN(new_n775));
  INV_X1    g589(.A(new_n479), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n694), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT116), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT116), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n759), .A2(new_n338), .A3(new_n337), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT113), .Z(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n613), .ZN(new_n783));
  INV_X1    g597(.A(new_n726), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n779), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n706), .A2(new_n187), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT114), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n662), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n783), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT50), .Z(new_n791));
  NOR2_X1   g605(.A1(new_n706), .A2(new_n726), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT115), .Z(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n645), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n528), .A2(new_n339), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n680), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n797), .A2(new_n684), .A3(new_n605), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n786), .A2(KEYINPUT51), .A3(new_n791), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n783), .A2(new_n707), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n801), .B(new_n337), .C1(new_n608), .C2(new_n797), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n794), .A2(new_n698), .A3(new_n724), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT48), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT48), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n778), .A2(new_n785), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n799), .A2(new_n791), .A3(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n800), .B(new_n806), .C1(new_n808), .C2(KEYINPUT51), .ZN(new_n809));
  INV_X1    g623(.A(new_n735), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n733), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n701), .A2(new_n709), .A3(new_n704), .A4(new_n717), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n784), .A2(new_n336), .A3(new_n663), .ZN(new_n813));
  INV_X1    g627(.A(new_n652), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n650), .A3(new_n585), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n720), .A2(new_n727), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n738), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n811), .A2(new_n812), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n290), .A2(new_n342), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n614), .A2(new_n607), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n591), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT106), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n591), .A2(KEYINPUT106), .A3(new_n822), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n336), .A2(new_n684), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT107), .Z(new_n828));
  NAND3_X1  g642(.A1(new_n614), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n646), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n825), .A2(new_n826), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT108), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT106), .B1(new_n591), .B2(new_n822), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n830), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT108), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n826), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n819), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n655), .A2(new_n686), .A3(new_n721), .ZN(new_n839));
  INV_X1    g653(.A(new_n286), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n285), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n289), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n712), .A3(new_n715), .A4(new_n187), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n476), .B1(new_n691), .B2(new_n417), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n776), .B1(new_n844), .B2(new_n475), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n644), .A3(new_n651), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT97), .B1(new_n569), .B2(new_n671), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT97), .A2(new_n671), .A3(new_n673), .A4(new_n674), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n848), .B1(new_n679), .B2(new_n847), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n839), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n847), .B1(new_n850), .B2(new_n849), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT109), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n851), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(KEYINPUT110), .A3(new_n839), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n838), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n860), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n861), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n865), .B2(new_n866), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n709), .A2(new_n704), .A3(new_n701), .A4(new_n717), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n736), .A2(new_n874), .A3(new_n817), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n836), .B1(new_n835), .B2(new_n826), .ZN(new_n876));
  INV_X1    g690(.A(new_n826), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n877), .A2(new_n834), .A3(KEYINPUT108), .A4(new_n830), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n854), .A2(new_n855), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT110), .B1(new_n859), .B2(new_n839), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n860), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n873), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n729), .A2(KEYINPUT53), .A3(new_n732), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n874), .A2(new_n817), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n864), .B(new_n888), .C1(new_n878), .C2(new_n876), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n872), .A2(new_n891), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n809), .A2(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n694), .B(KEYINPUT49), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n776), .A2(new_n188), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n698), .A3(new_n757), .A4(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(new_n662), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n679), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n217), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT53), .B1(new_n869), .B2(new_n838), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n888), .B1(new_n876), .B2(new_n878), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n883), .A2(new_n862), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n327), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n906), .A2(new_n287), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n270), .A2(new_n272), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n221), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n900), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(G210), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n914), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(G51));
  INV_X1    g730(.A(new_n890), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n901), .B2(new_n904), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(KEYINPUT117), .A3(new_n891), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n917), .C1(new_n901), .C2(new_n904), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n476), .B(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT118), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n919), .A2(new_n925), .A3(new_n921), .A4(new_n922), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n466), .A2(new_n469), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT119), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n744), .A2(new_n745), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n906), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n899), .B1(new_n929), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n400), .A2(new_n389), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n933), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n899), .ZN(G60));
  NAND2_X1  g752(.A1(new_n599), .A2(new_n600), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT59), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n892), .B2(new_n942), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n940), .A2(new_n919), .A3(new_n921), .A4(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n944), .A3(new_n899), .ZN(G63));
  XNOR2_X1  g759(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n905), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n633), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n521), .B(KEYINPUT121), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n905), .B2(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n900), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G66));
  AOI21_X1  g769(.A(new_n217), .B1(new_n340), .B2(G224), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n874), .B1(new_n833), .B2(new_n837), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n958), .B2(new_n217), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n908), .B1(G898), .B2(new_n217), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT122), .Z(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  NOR2_X1   g776(.A1(new_n535), .A2(new_n539), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n396), .B1(new_n395), .B2(new_n362), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n839), .B(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n665), .A2(new_n680), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n773), .B(new_n765), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n828), .A2(new_n607), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n972), .A2(new_n658), .A3(new_n726), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n582), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n967), .B1(new_n680), .B2(new_n665), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(KEYINPUT62), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n965), .B1(new_n977), .B2(G953), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n965), .B1(G900), .B2(G953), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n967), .A2(new_n811), .A3(new_n738), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n725), .A2(new_n843), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n751), .A2(new_n754), .A3(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n980), .A2(new_n773), .A3(new_n765), .A4(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n979), .B1(new_n983), .B2(G953), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n978), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G72));
  AOI21_X1  g802(.A(new_n551), .B1(new_n540), .B2(new_n542), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n977), .A2(new_n957), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  AOI21_X1  g806(.A(KEYINPUT125), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n994));
  INV_X1    g808(.A(new_n992), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n994), .B(new_n995), .C1(new_n977), .C2(new_n957), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n989), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n576), .A2(new_n998), .B1(new_n540), .B2(new_n548), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n998), .B2(new_n576), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n992), .B(new_n1000), .C1(new_n867), .C2(new_n871), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n992), .B1(new_n983), .B2(new_n958), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n560), .A2(new_n575), .A3(new_n546), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n899), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n997), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(KEYINPUT127), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n997), .A2(new_n1007), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(G57));
endmodule


