

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742;

  AND2_X1 U365 ( .A1(n368), .A2(KEYINPUT80), .ZN(n661) );
  XNOR2_X1 U366 ( .A(n563), .B(n562), .ZN(n737) );
  BUF_X1 U367 ( .A(n495), .Z(n554) );
  XNOR2_X1 U368 ( .A(n484), .B(KEYINPUT4), .ZN(n723) );
  INV_X2 U369 ( .A(G953), .ZN(n717) );
  AND2_X2 U370 ( .A1(n363), .A2(n352), .ZN(n351) );
  NOR2_X1 U371 ( .A1(n575), .A2(KEYINPUT76), .ZN(n576) );
  NOR2_X2 U372 ( .A1(n589), .A2(n739), .ZN(n378) );
  NOR2_X2 U373 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X2 U374 ( .A1(n353), .A2(n658), .ZN(n728) );
  XNOR2_X2 U375 ( .A(n355), .B(n354), .ZN(n353) );
  XNOR2_X2 U376 ( .A(n491), .B(n490), .ZN(n538) );
  XNOR2_X2 U377 ( .A(n554), .B(KEYINPUT38), .ZN(n667) );
  NOR2_X1 U378 ( .A1(n688), .A2(n535), .ZN(n514) );
  INV_X1 U379 ( .A(KEYINPUT84), .ZN(n354) );
  NAND2_X1 U380 ( .A1(n357), .A2(n356), .ZN(n355) );
  AND2_X1 U381 ( .A1(n386), .A2(n385), .ZN(n384) );
  NOR2_X1 U382 ( .A1(n529), .A2(n528), .ZN(n386) );
  NOR2_X2 U383 ( .A1(n595), .A2(n741), .ZN(n596) );
  NOR2_X1 U384 ( .A1(n675), .A2(n535), .ZN(n537) );
  AND2_X1 U385 ( .A1(n561), .A2(n590), .ZN(n563) );
  XNOR2_X1 U386 ( .A(n534), .B(n533), .ZN(n675) );
  XNOR2_X1 U387 ( .A(n542), .B(n541), .ZN(n555) );
  XNOR2_X1 U388 ( .A(n516), .B(KEYINPUT1), .ZN(n375) );
  XNOR2_X1 U389 ( .A(n450), .B(n449), .ZN(n716) );
  XNOR2_X1 U390 ( .A(n429), .B(n428), .ZN(n450) );
  INV_X1 U391 ( .A(KEYINPUT109), .ZN(n562) );
  OR2_X1 U392 ( .A1(n540), .A2(n538), .ZN(n653) );
  XNOR2_X2 U393 ( .A(n421), .B(n420), .ZN(n484) );
  OR2_X1 U394 ( .A1(n637), .A2(G902), .ZN(n447) );
  XOR2_X1 U395 ( .A(KEYINPUT81), .B(n669), .Z(n572) );
  NAND2_X1 U396 ( .A1(n548), .A2(KEYINPUT66), .ZN(n371) );
  INV_X1 U397 ( .A(KEYINPUT73), .ZN(n369) );
  NOR2_X2 U398 ( .A1(G953), .A2(G237), .ZN(n465) );
  OR2_X1 U399 ( .A1(n685), .A2(n558), .ZN(n559) );
  INV_X1 U400 ( .A(KEYINPUT2), .ZN(n367) );
  NAND2_X1 U401 ( .A1(n494), .A2(n667), .ZN(n360) );
  NAND2_X1 U402 ( .A1(n590), .A2(n667), .ZN(n592) );
  AND2_X1 U403 ( .A1(n448), .A2(n516), .ZN(n565) );
  NAND2_X1 U404 ( .A1(n701), .A2(G472), .ZN(n625) );
  NAND2_X1 U405 ( .A1(n530), .A2(KEYINPUT66), .ZN(n546) );
  XNOR2_X1 U406 ( .A(G119), .B(G116), .ZN(n426) );
  XNOR2_X1 U407 ( .A(G146), .B(G125), .ZN(n452) );
  NAND2_X1 U408 ( .A1(n389), .A2(n630), .ZN(n388) );
  NAND2_X1 U409 ( .A1(n519), .A2(n653), .ZN(n669) );
  INV_X1 U410 ( .A(G237), .ZN(n460) );
  NAND2_X1 U411 ( .A1(G953), .A2(G902), .ZN(n497) );
  XOR2_X1 U412 ( .A(G137), .B(KEYINPUT5), .Z(n424) );
  XNOR2_X1 U413 ( .A(n452), .B(n382), .ZN(n403) );
  INV_X1 U414 ( .A(KEYINPUT10), .ZN(n382) );
  XNOR2_X1 U415 ( .A(G134), .B(G131), .ZN(n724) );
  XNOR2_X1 U416 ( .A(n376), .B(n597), .ZN(n357) );
  AND2_X1 U417 ( .A1(n372), .A2(n374), .ZN(n682) );
  NAND2_X1 U418 ( .A1(n509), .A2(n678), .ZN(n679) );
  NAND2_X1 U419 ( .A1(n375), .A2(n681), .ZN(n531) );
  XNOR2_X1 U420 ( .A(G128), .B(G119), .ZN(n407) );
  XNOR2_X1 U421 ( .A(n403), .B(n442), .ZN(n727) );
  XNOR2_X1 U422 ( .A(G122), .B(KEYINPUT7), .ZN(n479) );
  XOR2_X1 U423 ( .A(KEYINPUT9), .B(KEYINPUT98), .Z(n480) );
  XNOR2_X1 U424 ( .A(G116), .B(G134), .ZN(n482) );
  INV_X1 U425 ( .A(G128), .ZN(n420) );
  XOR2_X1 U426 ( .A(KEYINPUT12), .B(G140), .Z(n472) );
  XOR2_X1 U427 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n467) );
  XNOR2_X1 U428 ( .A(G143), .B(G131), .ZN(n469) );
  XOR2_X1 U429 ( .A(G137), .B(G140), .Z(n442) );
  OR2_X1 U430 ( .A1(n372), .A2(n373), .ZN(n524) );
  XNOR2_X1 U431 ( .A(n507), .B(n391), .ZN(n361) );
  INV_X1 U432 ( .A(KEYINPUT22), .ZN(n391) );
  XNOR2_X1 U433 ( .A(n559), .B(n380), .ZN(n379) );
  INV_X1 U434 ( .A(KEYINPUT30), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n478), .B(n477), .ZN(n540) );
  NAND2_X1 U436 ( .A1(n366), .A2(n362), .ZN(n349) );
  NOR2_X1 U437 ( .A1(n728), .A2(n367), .ZN(n362) );
  AND2_X1 U438 ( .A1(n612), .A2(G953), .ZN(n705) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n394) );
  XNOR2_X1 U440 ( .A(n359), .B(n358), .ZN(n595) );
  INV_X1 U441 ( .A(KEYINPUT42), .ZN(n358) );
  XNOR2_X1 U442 ( .A(n594), .B(n593), .ZN(n741) );
  AND2_X1 U443 ( .A1(n540), .A2(n538), .ZN(n646) );
  AND2_X1 U444 ( .A1(n546), .A2(n550), .ZN(n344) );
  XOR2_X1 U445 ( .A(n409), .B(n408), .Z(n345) );
  INV_X1 U446 ( .A(n681), .ZN(n374) );
  INV_X1 U447 ( .A(n509), .ZN(n373) );
  NOR2_X1 U448 ( .A1(n582), .A2(n509), .ZN(n346) );
  XOR2_X1 U449 ( .A(n504), .B(KEYINPUT0), .Z(n347) );
  XOR2_X1 U450 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n348) );
  AND2_X4 U451 ( .A1(n350), .A2(n349), .ZN(n701) );
  AND2_X2 U452 ( .A1(n364), .A2(n351), .ZN(n350) );
  INV_X1 U453 ( .A(n607), .ZN(n352) );
  INV_X1 U454 ( .A(n375), .ZN(n372) );
  AND2_X1 U455 ( .A1(n553), .A2(n629), .ZN(n389) );
  XNOR2_X2 U456 ( .A(n545), .B(n544), .ZN(n629) );
  INV_X1 U457 ( .A(n742), .ZN(n356) );
  NAND2_X1 U458 ( .A1(n690), .A2(n565), .ZN(n359) );
  XNOR2_X2 U459 ( .A(n360), .B(KEYINPUT41), .ZN(n690) );
  NAND2_X1 U460 ( .A1(n361), .A2(n526), .ZN(n527) );
  AND2_X1 U461 ( .A1(n361), .A2(n372), .ZN(n511) );
  INV_X1 U462 ( .A(n706), .ZN(n366) );
  NAND2_X1 U463 ( .A1(n728), .A2(n367), .ZN(n363) );
  NAND2_X1 U464 ( .A1(n706), .A2(n367), .ZN(n364) );
  NAND2_X1 U465 ( .A1(n366), .A2(n365), .ZN(n368) );
  INV_X1 U466 ( .A(n728), .ZN(n365) );
  OR2_X2 U467 ( .A1(n531), .A2(n685), .ZN(n513) );
  NAND2_X1 U468 ( .A1(n344), .A2(n371), .ZN(n370) );
  NAND2_X1 U469 ( .A1(n547), .A2(KEYINPUT44), .ZN(n385) );
  OR2_X2 U470 ( .A1(n579), .A2(n578), .ZN(n589) );
  NOR2_X2 U471 ( .A1(n512), .A2(n509), .ZN(n681) );
  NOR2_X1 U472 ( .A1(n557), .A2(n560), .ZN(n381) );
  AND2_X1 U473 ( .A1(n381), .A2(n379), .ZN(n590) );
  NAND2_X1 U474 ( .A1(n370), .A2(n369), .ZN(n390) );
  NOR2_X1 U475 ( .A1(n375), .A2(n598), .ZN(n599) );
  NAND2_X1 U476 ( .A1(n587), .A2(n375), .ZN(n588) );
  NAND2_X1 U477 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U478 ( .A(n596), .B(KEYINPUT46), .ZN(n377) );
  INV_X1 U479 ( .A(n403), .ZN(n473) );
  XNOR2_X2 U480 ( .A(n383), .B(n348), .ZN(n706) );
  NAND2_X1 U481 ( .A1(n387), .A2(n384), .ZN(n383) );
  NAND2_X1 U482 ( .A1(n390), .A2(n388), .ZN(n387) );
  XNOR2_X1 U483 ( .A(n583), .B(n496), .ZN(n566) );
  OR2_X2 U484 ( .A1(n495), .A2(n558), .ZN(n583) );
  XNOR2_X2 U485 ( .A(n592), .B(n591), .ZN(n606) );
  XNOR2_X1 U486 ( .A(n464), .B(n463), .ZN(n495) );
  NAND2_X1 U487 ( .A1(n459), .A2(n607), .ZN(n464) );
  NAND2_X1 U488 ( .A1(n570), .A2(KEYINPUT47), .ZN(n392) );
  XNOR2_X1 U489 ( .A(n737), .B(KEYINPUT82), .ZN(n564) );
  NAND2_X1 U490 ( .A1(n630), .A2(n549), .ZN(n530) );
  BUF_X1 U491 ( .A(n566), .Z(n567) );
  INV_X1 U492 ( .A(KEYINPUT40), .ZN(n593) );
  INV_X1 U493 ( .A(KEYINPUT14), .ZN(n393) );
  XNOR2_X1 U494 ( .A(n394), .B(n393), .ZN(n697) );
  NOR2_X1 U495 ( .A1(n697), .A2(n497), .ZN(n395) );
  XNOR2_X1 U496 ( .A(n395), .B(KEYINPUT105), .ZN(n396) );
  NOR2_X1 U497 ( .A1(G900), .A2(n396), .ZN(n397) );
  XNOR2_X1 U498 ( .A(n397), .B(KEYINPUT106), .ZN(n399) );
  NAND2_X1 U499 ( .A1(n717), .A2(G952), .ZN(n498) );
  NOR2_X1 U500 ( .A1(n498), .A2(n697), .ZN(n398) );
  NOR2_X1 U501 ( .A1(n399), .A2(n398), .ZN(n560) );
  XNOR2_X1 U502 ( .A(KEYINPUT15), .B(G902), .ZN(n607) );
  NAND2_X1 U503 ( .A1(G234), .A2(n607), .ZN(n400) );
  XNOR2_X1 U504 ( .A(KEYINPUT20), .B(n400), .ZN(n414) );
  NAND2_X1 U505 ( .A1(G221), .A2(n414), .ZN(n401) );
  XNOR2_X1 U506 ( .A(n401), .B(KEYINPUT21), .ZN(n678) );
  NOR2_X1 U507 ( .A1(n560), .A2(n678), .ZN(n402) );
  XNOR2_X1 U508 ( .A(KEYINPUT68), .B(n402), .ZN(n419) );
  XOR2_X1 U509 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n405) );
  XNOR2_X1 U510 ( .A(G110), .B(KEYINPUT70), .ZN(n404) );
  XNOR2_X1 U511 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U512 ( .A(n727), .B(n406), .ZN(n413) );
  XNOR2_X1 U513 ( .A(n407), .B(KEYINPUT24), .ZN(n409) );
  XOR2_X1 U514 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n408) );
  NAND2_X1 U515 ( .A1(G234), .A2(n717), .ZN(n410) );
  XOR2_X1 U516 ( .A(KEYINPUT8), .B(n410), .Z(n485) );
  NAND2_X1 U517 ( .A1(n485), .A2(G221), .ZN(n411) );
  XOR2_X1 U518 ( .A(n345), .B(n411), .Z(n412) );
  XNOR2_X1 U519 ( .A(n413), .B(n412), .ZN(n632) );
  INV_X1 U520 ( .A(G902), .ZN(n489) );
  NAND2_X1 U521 ( .A1(n632), .A2(n489), .ZN(n418) );
  NAND2_X1 U522 ( .A1(G217), .A2(n414), .ZN(n416) );
  XOR2_X1 U523 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n415) );
  XNOR2_X1 U524 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X2 U525 ( .A(n418), .B(n417), .ZN(n509) );
  NAND2_X1 U526 ( .A1(n419), .A2(n509), .ZN(n580) );
  XNOR2_X2 U527 ( .A(G143), .B(KEYINPUT65), .ZN(n421) );
  XNOR2_X1 U528 ( .A(KEYINPUT67), .B(G101), .ZN(n422) );
  XNOR2_X2 U529 ( .A(n723), .B(n422), .ZN(n440) );
  XNOR2_X1 U530 ( .A(n724), .B(G146), .ZN(n444) );
  NAND2_X1 U531 ( .A1(n465), .A2(G210), .ZN(n423) );
  XNOR2_X1 U532 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U533 ( .A(n444), .B(n425), .ZN(n430) );
  XNOR2_X1 U534 ( .A(n426), .B(KEYINPUT3), .ZN(n429) );
  INV_X1 U535 ( .A(KEYINPUT88), .ZN(n427) );
  XNOR2_X1 U536 ( .A(n427), .B(G113), .ZN(n428) );
  XNOR2_X1 U537 ( .A(n430), .B(n450), .ZN(n431) );
  XNOR2_X1 U538 ( .A(n440), .B(n431), .ZN(n623) );
  NAND2_X1 U539 ( .A1(n623), .A2(n489), .ZN(n435) );
  XNOR2_X1 U540 ( .A(KEYINPUT75), .B(KEYINPUT95), .ZN(n433) );
  INV_X1 U541 ( .A(G472), .ZN(n432) );
  XNOR2_X1 U542 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X2 U543 ( .A(n435), .B(n434), .ZN(n685) );
  NOR2_X1 U544 ( .A1(n580), .A2(n685), .ZN(n436) );
  XNOR2_X1 U545 ( .A(n436), .B(KEYINPUT28), .ZN(n448) );
  XNOR2_X1 U546 ( .A(G104), .B(G110), .ZN(n437) );
  XNOR2_X1 U547 ( .A(n437), .B(G107), .ZN(n714) );
  XNOR2_X1 U548 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n438) );
  XNOR2_X1 U549 ( .A(n714), .B(n438), .ZN(n439) );
  XNOR2_X2 U550 ( .A(n440), .B(n439), .ZN(n458) );
  NAND2_X1 U551 ( .A1(G227), .A2(n717), .ZN(n441) );
  XNOR2_X1 U552 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U554 ( .A(n458), .B(n445), .ZN(n637) );
  XOR2_X1 U555 ( .A(KEYINPUT69), .B(G469), .Z(n446) );
  XNOR2_X2 U556 ( .A(n447), .B(n446), .ZN(n516) );
  XNOR2_X1 U557 ( .A(KEYINPUT16), .B(G122), .ZN(n449) );
  XNOR2_X1 U558 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n452), .B(n451), .ZN(n455) );
  NAND2_X1 U560 ( .A1(n717), .A2(G224), .ZN(n453) );
  XNOR2_X1 U561 ( .A(n453), .B(KEYINPUT89), .ZN(n454) );
  XNOR2_X1 U562 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U563 ( .A(n716), .B(n456), .ZN(n457) );
  XNOR2_X1 U564 ( .A(n458), .B(n457), .ZN(n608) );
  INV_X1 U565 ( .A(n608), .ZN(n459) );
  NAND2_X1 U566 ( .A1(n489), .A2(n460), .ZN(n493) );
  NAND2_X1 U567 ( .A1(n493), .A2(G210), .ZN(n462) );
  INV_X1 U568 ( .A(KEYINPUT79), .ZN(n461) );
  XNOR2_X1 U569 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U570 ( .A1(G214), .A2(n465), .ZN(n466) );
  XNOR2_X1 U571 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U572 ( .A(n468), .B(G104), .Z(n470) );
  XNOR2_X1 U573 ( .A(n470), .B(n469), .ZN(n476) );
  XNOR2_X1 U574 ( .A(G113), .B(G122), .ZN(n471) );
  XNOR2_X1 U575 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U576 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U577 ( .A(n476), .B(n475), .ZN(n617) );
  NAND2_X1 U578 ( .A1(n617), .A2(n489), .ZN(n478) );
  XNOR2_X1 U579 ( .A(KEYINPUT13), .B(G475), .ZN(n477) );
  INV_X1 U580 ( .A(n540), .ZN(n492) );
  XNOR2_X1 U581 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U582 ( .A(n481), .B(G107), .Z(n483) );
  XNOR2_X1 U583 ( .A(n483), .B(n482), .ZN(n488) );
  AND2_X1 U584 ( .A1(G217), .A2(n485), .ZN(n486) );
  XNOR2_X1 U585 ( .A(n484), .B(n486), .ZN(n487) );
  XNOR2_X1 U586 ( .A(n488), .B(n487), .ZN(n703) );
  NAND2_X1 U587 ( .A1(n703), .A2(n489), .ZN(n491) );
  XOR2_X1 U588 ( .A(KEYINPUT99), .B(G478), .Z(n490) );
  OR2_X1 U589 ( .A1(n492), .A2(n538), .ZN(n664) );
  NAND2_X1 U590 ( .A1(n493), .A2(G214), .ZN(n668) );
  INV_X1 U591 ( .A(n668), .ZN(n558) );
  NOR2_X1 U592 ( .A1(n664), .A2(n558), .ZN(n494) );
  XOR2_X1 U593 ( .A(n595), .B(G137), .Z(G39) );
  INV_X1 U594 ( .A(KEYINPUT19), .ZN(n496) );
  INV_X1 U595 ( .A(n697), .ZN(n502) );
  NOR2_X1 U596 ( .A1(G898), .A2(n497), .ZN(n500) );
  INV_X1 U597 ( .A(n498), .ZN(n499) );
  OR2_X1 U598 ( .A1(n500), .A2(n499), .ZN(n501) );
  NAND2_X1 U599 ( .A1(n502), .A2(n501), .ZN(n503) );
  OR2_X2 U600 ( .A1(n566), .A2(n503), .ZN(n505) );
  INV_X1 U601 ( .A(KEYINPUT87), .ZN(n504) );
  XNOR2_X2 U602 ( .A(n505), .B(n347), .ZN(n515) );
  XNOR2_X1 U603 ( .A(n678), .B(KEYINPUT94), .ZN(n512) );
  NOR2_X1 U604 ( .A1(n664), .A2(n512), .ZN(n506) );
  NAND2_X1 U605 ( .A1(n515), .A2(n506), .ZN(n507) );
  XOR2_X1 U606 ( .A(KEYINPUT6), .B(KEYINPUT101), .Z(n508) );
  XNOR2_X1 U607 ( .A(n685), .B(n508), .ZN(n582) );
  NAND2_X1 U608 ( .A1(n511), .A2(n346), .ZN(n521) );
  XNOR2_X1 U609 ( .A(n521), .B(G101), .ZN(G3) );
  INV_X1 U610 ( .A(n685), .ZN(n517) );
  NOR2_X1 U611 ( .A1(n517), .A2(n373), .ZN(n510) );
  NAND2_X1 U612 ( .A1(n511), .A2(n510), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(G110), .ZN(G12) );
  XNOR2_X1 U614 ( .A(n513), .B(KEYINPUT96), .ZN(n688) );
  INV_X1 U615 ( .A(n515), .ZN(n535) );
  XNOR2_X1 U616 ( .A(n514), .B(KEYINPUT31), .ZN(n655) );
  NAND2_X1 U617 ( .A1(n516), .A2(n681), .ZN(n557) );
  NOR2_X1 U618 ( .A1(n557), .A2(n517), .ZN(n518) );
  NAND2_X1 U619 ( .A1(n515), .A2(n518), .ZN(n642) );
  NAND2_X1 U620 ( .A1(n655), .A2(n642), .ZN(n520) );
  XNOR2_X1 U621 ( .A(n646), .B(KEYINPUT100), .ZN(n605) );
  INV_X1 U622 ( .A(n605), .ZN(n519) );
  NAND2_X1 U623 ( .A1(n520), .A2(n572), .ZN(n522) );
  NAND2_X1 U624 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U625 ( .A(n523), .B(KEYINPUT102), .ZN(n529) );
  XNOR2_X1 U626 ( .A(n582), .B(KEYINPUT78), .ZN(n525) );
  NOR2_X1 U627 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X2 U628 ( .A(n527), .B(KEYINPUT32), .ZN(n630) );
  NOR2_X1 U629 ( .A1(n530), .A2(KEYINPUT66), .ZN(n528) );
  INV_X1 U630 ( .A(n531), .ZN(n532) );
  NAND2_X1 U631 ( .A1(n532), .A2(n582), .ZN(n534) );
  XNOR2_X1 U632 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n533) );
  XOR2_X1 U633 ( .A(KEYINPUT77), .B(KEYINPUT34), .Z(n536) );
  XNOR2_X1 U634 ( .A(n537), .B(n536), .ZN(n543) );
  INV_X1 U635 ( .A(n538), .ZN(n539) );
  OR2_X1 U636 ( .A1(n540), .A2(n539), .ZN(n542) );
  INV_X1 U637 ( .A(KEYINPUT104), .ZN(n541) );
  NAND2_X1 U638 ( .A1(n543), .A2(n555), .ZN(n545) );
  XNOR2_X1 U639 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n544) );
  NAND2_X1 U640 ( .A1(n546), .A2(n629), .ZN(n547) );
  INV_X1 U641 ( .A(n629), .ZN(n548) );
  INV_X1 U642 ( .A(KEYINPUT44), .ZN(n550) );
  INV_X1 U643 ( .A(n549), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n550), .A2(KEYINPUT73), .ZN(n551) );
  NOR2_X1 U645 ( .A1(n552), .A2(n551), .ZN(n553) );
  INV_X1 U646 ( .A(n555), .ZN(n556) );
  NOR2_X1 U647 ( .A1(n554), .A2(n556), .ZN(n561) );
  INV_X1 U648 ( .A(n564), .ZN(n571) );
  INV_X1 U649 ( .A(n565), .ZN(n568) );
  NOR2_X4 U650 ( .A1(n568), .A2(n567), .ZN(n651) );
  AND2_X1 U651 ( .A1(n669), .A2(KEYINPUT76), .ZN(n569) );
  NAND2_X1 U652 ( .A1(n651), .A2(n569), .ZN(n570) );
  NAND2_X1 U653 ( .A1(n571), .A2(n392), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n651), .A2(n572), .ZN(n575) );
  NOR2_X1 U655 ( .A1(n575), .A2(KEYINPUT47), .ZN(n574) );
  INV_X1 U656 ( .A(KEYINPUT76), .ZN(n573) );
  NOR2_X1 U657 ( .A1(n574), .A2(n573), .ZN(n577) );
  NOR2_X1 U658 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U659 ( .A1(n580), .A2(n653), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n598) );
  XNOR2_X1 U661 ( .A(KEYINPUT110), .B(n598), .ZN(n584) );
  NOR2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U663 ( .A(KEYINPUT86), .B(KEYINPUT36), .ZN(n585) );
  XNOR2_X1 U664 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U665 ( .A(n588), .B(KEYINPUT111), .ZN(n739) );
  XNOR2_X1 U666 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n591) );
  INV_X1 U667 ( .A(n653), .ZN(n650) );
  NAND2_X1 U668 ( .A1(n606), .A2(n650), .ZN(n594) );
  INV_X1 U669 ( .A(KEYINPUT48), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n668), .A2(n599), .ZN(n600) );
  XOR2_X1 U671 ( .A(KEYINPUT107), .B(n600), .Z(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT43), .B(n601), .Z(n603) );
  INV_X1 U673 ( .A(n554), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT108), .ZN(n742) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n658) );
  NAND2_X1 U677 ( .A1(n701), .A2(G210), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n609) );
  XNOR2_X1 U679 ( .A(n608), .B(n609), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U681 ( .A(G952), .ZN(n612) );
  NOR2_X2 U682 ( .A1(n613), .A2(n705), .ZN(n615) );
  XOR2_X1 U683 ( .A(KEYINPUT85), .B(KEYINPUT56), .Z(n614) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(G51) );
  NAND2_X1 U685 ( .A1(n701), .A2(G475), .ZN(n619) );
  XOR2_X1 U686 ( .A(KEYINPUT119), .B(KEYINPUT59), .Z(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X2 U689 ( .A1(n620), .A2(n705), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n621), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U691 ( .A(KEYINPUT112), .B(KEYINPUT62), .Z(n622) );
  XNOR2_X1 U692 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U694 ( .A1(n626), .A2(n705), .ZN(n628) );
  XNOR2_X1 U695 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(G57) );
  XNOR2_X1 U697 ( .A(n629), .B(G122), .ZN(G24) );
  XNOR2_X1 U698 ( .A(G119), .B(KEYINPUT127), .ZN(n631) );
  XOR2_X1 U699 ( .A(n631), .B(n630), .Z(G21) );
  NAND2_X1 U700 ( .A1(n701), .A2(G217), .ZN(n634) );
  XOR2_X1 U701 ( .A(n632), .B(KEYINPUT120), .Z(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X1 U703 ( .A1(n635), .A2(n705), .ZN(G66) );
  NAND2_X1 U704 ( .A1(n701), .A2(G469), .ZN(n639) );
  XOR2_X1 U705 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n636) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U708 ( .A1(n640), .A2(n705), .ZN(G54) );
  NOR2_X1 U709 ( .A1(n653), .A2(n642), .ZN(n641) );
  XOR2_X1 U710 ( .A(G104), .B(n641), .Z(G6) );
  INV_X1 U711 ( .A(n646), .ZN(n656) );
  NOR2_X1 U712 ( .A1(n656), .A2(n642), .ZN(n644) );
  XNOR2_X1 U713 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U715 ( .A(G107), .B(n645), .ZN(G9) );
  XOR2_X1 U716 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U717 ( .A1(n651), .A2(n646), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(G128), .B(n649), .ZN(G30) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n652), .B(G146), .ZN(G48) );
  NOR2_X1 U722 ( .A1(n653), .A2(n655), .ZN(n654) );
  XOR2_X1 U723 ( .A(G113), .B(n654), .Z(G15) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U725 ( .A(G116), .B(n657), .Z(G18) );
  XNOR2_X1 U726 ( .A(G134), .B(n658), .ZN(G36) );
  INV_X1 U727 ( .A(n690), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n675), .A2(n659), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n660), .A2(G953), .ZN(n663) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n661), .Z(n662) );
  NAND2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n699) );
  NOR2_X1 U732 ( .A1(n667), .A2(n668), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U734 ( .A(KEYINPUT117), .B(n666), .Z(n673) );
  INV_X1 U735 ( .A(n667), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U739 ( .A(KEYINPUT118), .B(n674), .Z(n677) );
  INV_X1 U740 ( .A(n675), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n693) );
  XNOR2_X1 U742 ( .A(n679), .B(KEYINPUT116), .ZN(n680) );
  XNOR2_X1 U743 ( .A(KEYINPUT49), .B(n680), .ZN(n684) );
  XNOR2_X1 U744 ( .A(KEYINPUT50), .B(n682), .ZN(n683) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U748 ( .A(KEYINPUT51), .B(n689), .Z(n691) );
  NAND2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U751 ( .A(KEYINPUT52), .B(n694), .ZN(n695) );
  NAND2_X1 U752 ( .A1(n695), .A2(G952), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U754 ( .A(KEYINPUT53), .B(n700), .ZN(G75) );
  NAND2_X1 U755 ( .A1(n701), .A2(G478), .ZN(n702) );
  XOR2_X1 U756 ( .A(n703), .B(n702), .Z(n704) );
  NOR2_X1 U757 ( .A1(n705), .A2(n704), .ZN(G63) );
  NOR2_X1 U758 ( .A1(n706), .A2(G953), .ZN(n712) );
  XOR2_X1 U759 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n708) );
  NAND2_X1 U760 ( .A1(G224), .A2(G953), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U762 ( .A1(G898), .A2(n709), .ZN(n710) );
  XOR2_X1 U763 ( .A(KEYINPUT122), .B(n710), .Z(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n713), .B(KEYINPUT123), .ZN(n721) );
  XOR2_X1 U766 ( .A(G101), .B(n714), .Z(n715) );
  XNOR2_X1 U767 ( .A(n716), .B(n715), .ZN(n719) );
  NOR2_X1 U768 ( .A1(G898), .A2(n717), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(KEYINPUT124), .B(n722), .ZN(G69) );
  INV_X1 U772 ( .A(n724), .ZN(n725) );
  XNOR2_X1 U773 ( .A(n723), .B(n725), .ZN(n726) );
  XNOR2_X1 U774 ( .A(n727), .B(n726), .ZN(n730) );
  XNOR2_X1 U775 ( .A(n728), .B(n730), .ZN(n729) );
  NOR2_X1 U776 ( .A1(n729), .A2(G953), .ZN(n735) );
  XNOR2_X1 U777 ( .A(n730), .B(KEYINPUT125), .ZN(n731) );
  XNOR2_X1 U778 ( .A(G227), .B(n731), .ZN(n733) );
  NAND2_X1 U779 ( .A1(G900), .A2(G953), .ZN(n732) );
  NOR2_X1 U780 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U781 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U782 ( .A(KEYINPUT126), .B(n736), .ZN(G72) );
  XNOR2_X1 U783 ( .A(G143), .B(n737), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n738), .B(KEYINPUT115), .ZN(G45) );
  XNOR2_X1 U785 ( .A(G125), .B(n739), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n740), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U787 ( .A(G131), .B(n741), .Z(G33) );
  XOR2_X1 U788 ( .A(G140), .B(n742), .Z(G42) );
endmodule

