//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT78), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT78), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  AOI21_X1  g006(.A(G107), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(G101), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n189), .A2(KEYINPUT3), .A3(G107), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n193), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n190), .A2(new_n192), .A3(G107), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n196), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT81), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT81), .B(new_n196), .C1(new_n200), .C2(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(G113), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT5), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(G119), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT5), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n212), .A2(KEYINPUT84), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT84), .B1(new_n212), .B2(new_n216), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G113), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n207), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT85), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n190), .A2(new_n192), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n194), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n197), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  INV_X1    g043(.A(new_n203), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n201), .B(new_n198), .C1(new_n193), .C2(new_n199), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(G101), .B1(new_n232), .B2(new_n233), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n219), .B(new_n220), .Z(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n233), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT78), .B(G104), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(new_n240), .B2(G107), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n241), .A2(KEYINPUT79), .A3(new_n201), .A4(new_n198), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n239), .A2(new_n226), .A3(G101), .A4(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n236), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n206), .A2(KEYINPUT85), .A3(new_n222), .A4(new_n207), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n225), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G110), .B(G122), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT86), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n225), .A2(new_n244), .A3(new_n250), .A4(new_n245), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n246), .A2(new_n253), .A3(new_n248), .ZN(new_n254));
  XNOR2_X1  g068(.A(G143), .B(G146), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G128), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(G143), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT64), .B1(new_n268), .B2(new_n255), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n258), .A2(G143), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G146), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n266), .A4(new_n267), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT65), .B1(new_n273), .B2(new_n267), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n255), .A2(new_n278), .A3(KEYINPUT0), .A4(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n265), .B1(new_n281), .B2(new_n264), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G224), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT87), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n282), .B(new_n285), .Z(new_n286));
  NAND3_X1  g100(.A1(new_n252), .A2(new_n254), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT88), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n252), .A2(KEYINPUT88), .A3(new_n254), .A4(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(KEYINPUT7), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n248), .B(KEYINPUT8), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n222), .A2(new_n204), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n221), .B1(new_n216), .B2(new_n212), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(new_n295), .C1(new_n204), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n282), .A2(new_n292), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n299), .B2(new_n251), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT89), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT90), .ZN(new_n304));
  INV_X1    g118(.A(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n289), .B2(new_n290), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT89), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n304), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n188), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT11), .ZN(new_n314));
  INV_X1    g128(.A(G134), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G137), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT11), .A3(G134), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(G131), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n316), .A2(new_n318), .A3(new_n322), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n276), .A2(new_n324), .A3(new_n280), .ZN(new_n325));
  INV_X1    g139(.A(new_n319), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n315), .A2(G137), .ZN(new_n327));
  OAI21_X1  g141(.A(G131), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n262), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n238), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n237), .A3(new_n329), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n313), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n313), .B2(new_n332), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n335));
  INV_X1    g149(.A(G210), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n336), .A2(G237), .A3(G953), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n335), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(G101), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT69), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n332), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n332), .B2(new_n340), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n330), .A2(new_n346), .A3(KEYINPUT30), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT66), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(KEYINPUT30), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n325), .A2(new_n329), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT67), .B1(new_n352), .B2(new_n238), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n354), .B(new_n237), .C1(new_n347), .C2(new_n351), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n345), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT31), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI211_X1 g172(.A(KEYINPUT66), .B(new_n348), .C1(new_n325), .C2(new_n329), .ZN(new_n359));
  AND4_X1   g173(.A1(new_n325), .A2(new_n329), .A3(new_n349), .A4(new_n350), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n238), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n354), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n352), .A2(KEYINPUT67), .A3(new_n238), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(KEYINPUT31), .A3(new_n345), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n341), .B1(new_n358), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT70), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n341), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT31), .B1(new_n364), .B2(new_n345), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n343), .A2(new_n344), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n357), .B(new_n372), .C1(new_n362), .C2(new_n363), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n367), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT32), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n369), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G472), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n331), .A2(new_n332), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT28), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT71), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n332), .A2(new_n313), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n333), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n334), .B2(new_n340), .ZN(new_n389));
  INV_X1    g203(.A(new_n332), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n362), .B2(new_n363), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n391), .B2(new_n340), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n379), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n366), .A2(new_n368), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(KEYINPUT32), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n378), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  INV_X1    g211(.A(G902), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(G234), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G125), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n264), .A2(G140), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT75), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n401), .A2(KEYINPUT75), .A3(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n404), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G146), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n258), .B(new_n404), .C1(new_n409), .C2(new_n403), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n213), .A2(G128), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n213), .A2(G128), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n414), .B(new_n415), .C1(new_n416), .C2(KEYINPUT23), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G110), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT24), .B(G110), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n416), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n426), .A2(new_n415), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n424), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n413), .B(new_n422), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n402), .A2(new_n405), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n258), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n417), .A2(G110), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n427), .B1(new_n425), .B2(new_n428), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n411), .B(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT22), .B(G137), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n438), .B(new_n439), .Z(new_n440));
  NAND3_X1  g254(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n432), .B2(new_n437), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT25), .A3(new_n398), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n398), .A3(new_n441), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n400), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n444), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n399), .A2(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT76), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n396), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n206), .A2(new_n262), .A3(new_n207), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT10), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n461));
  OAI21_X1  g275(.A(G128), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n259), .A2(KEYINPUT80), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n273), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n464), .A2(new_n257), .ZN(new_n465));
  OR3_X1    g279(.A1(new_n465), .A2(KEYINPUT10), .A3(new_n204), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n324), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n236), .A2(new_n281), .A3(new_n243), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT12), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n464), .A2(new_n257), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n229), .A2(new_n230), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n196), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n204), .A2(new_n263), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n472), .B1(new_n477), .B2(new_n324), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n479));
  AOI211_X1 g293(.A(new_n468), .B(new_n479), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n470), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G110), .B(G140), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n283), .A2(G227), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n457), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n465), .A2(new_n204), .A3(KEYINPUT10), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n458), .B2(KEYINPUT10), .ZN(new_n488));
  INV_X1    g302(.A(new_n469), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n324), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n470), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n485), .ZN(new_n492));
  INV_X1    g306(.A(new_n485), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n470), .A2(new_n481), .A3(KEYINPUT83), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n486), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G469), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n398), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n482), .A2(new_n485), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n470), .A3(new_n493), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(G469), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G469), .A2(G902), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G221), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT9), .B(G234), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n504), .B1(new_n506), .B2(new_n398), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT77), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT20), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT91), .B(G143), .ZN(new_n512));
  INV_X1    g326(.A(G214), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n513), .A2(G237), .A3(G953), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G237), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n283), .A3(G214), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G143), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n514), .B1(new_n518), .B2(G143), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(new_n322), .C1(new_n512), .C2(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT19), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n407), .B2(new_n408), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n433), .A2(KEYINPUT19), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n258), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n411), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n530));
  OAI221_X1 g344(.A(new_n522), .B1(new_n530), .B2(new_n322), .C1(new_n514), .C2(new_n512), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n434), .B1(new_n409), .B2(new_n258), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n531), .B(new_n532), .C1(new_n530), .C2(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G113), .B(G122), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n189), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n521), .A2(new_n523), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT17), .B(G131), .C1(new_n515), .C2(new_n520), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n540), .A2(new_n411), .A3(new_n412), .A4(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n536), .B(KEYINPUT92), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n533), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G475), .A2(G902), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n511), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n511), .A3(new_n546), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(KEYINPUT93), .B2(new_n548), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n548), .A2(KEYINPUT93), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n544), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n536), .B1(new_n542), .B2(new_n533), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n398), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G475), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT95), .B(G952), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  NAND2_X1  g371(.A1(G234), .A2(G237), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT21), .B(G898), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(G902), .A3(G953), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n505), .A2(new_n397), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G116), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n209), .A2(G122), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n194), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n271), .A2(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n260), .A2(G143), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n315), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n315), .B1(new_n569), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT94), .B1(new_n567), .B2(KEYINPUT14), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT14), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n209), .A4(G122), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n567), .A2(KEYINPUT14), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n575), .A2(new_n566), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n574), .B1(G107), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n566), .A2(new_n567), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G107), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n568), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n260), .B2(G143), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n570), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n569), .A2(new_n585), .ZN(new_n588));
  OAI21_X1  g402(.A(G134), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n589), .A3(new_n571), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n564), .B1(new_n581), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n564), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n580), .A2(G107), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n590), .B(new_n593), .C1(new_n594), .C2(new_n574), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n398), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G478), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(KEYINPUT15), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n598), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n592), .A2(new_n398), .A3(new_n595), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n551), .A2(new_n555), .A3(new_n563), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n510), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n312), .A2(new_n456), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  AOI21_X1  g421(.A(new_n310), .B1(new_n291), .B2(new_n300), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n304), .B(new_n305), .C1(new_n289), .C2(new_n290), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n187), .B(new_n563), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n596), .A2(new_n597), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n592), .A2(new_n612), .A3(new_n595), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n613), .A2(KEYINPUT96), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT97), .B1(new_n581), .B2(new_n591), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n615), .A2(new_n564), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n564), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(KEYINPUT33), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(KEYINPUT96), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n597), .A2(G902), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n614), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n551), .A2(new_n555), .B1(new_n611), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n610), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n366), .B2(G902), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n369), .A2(new_n625), .A3(new_n376), .A4(new_n455), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n510), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n545), .A2(new_n546), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT20), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n548), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n555), .A3(new_n602), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n610), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n627), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NAND3_X1  g452(.A1(new_n369), .A2(new_n625), .A3(new_n376), .ZN(new_n639));
  INV_X1    g453(.A(new_n453), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n432), .A2(new_n437), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  INV_X1    g456(.A(new_n440), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n642), .A2(KEYINPUT36), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(KEYINPUT36), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n640), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n445), .A2(new_n449), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n399), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n639), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n312), .A2(new_n605), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(new_n634), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n562), .A2(G900), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n559), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(KEYINPUT99), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  INV_X1    g475(.A(new_n659), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n634), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n652), .B(new_n664), .C1(new_n378), .C2(new_n395), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n508), .B1(new_n497), .B2(new_n502), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n666), .B(new_n187), .C1(new_n609), .C2(new_n608), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  NAND2_X1  g484(.A1(new_n309), .A2(new_n311), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n309), .A2(new_n673), .A3(new_n311), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n659), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  INV_X1    g493(.A(new_n340), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n380), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n356), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n379), .B1(new_n682), .B2(new_n398), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n394), .B2(KEYINPUT32), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n378), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n603), .B1(new_n551), .B2(new_n555), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n652), .A2(new_n686), .A3(new_n187), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n675), .A2(new_n678), .A3(new_n679), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NAND3_X1  g504(.A1(new_n651), .A2(new_n622), .A3(new_n659), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n396), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT100), .B1(new_n693), .B2(new_n667), .ZN(new_n694));
  INV_X1    g508(.A(new_n608), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n188), .B1(new_n695), .B2(new_n311), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n691), .B1(new_n378), .B2(new_n395), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n666), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NAND2_X1  g515(.A1(new_n495), .A2(new_n398), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G469), .ZN(new_n703));
  INV_X1    g517(.A(new_n507), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n497), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n396), .A2(new_n705), .A3(new_n455), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n624), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n635), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  AOI211_X1 g525(.A(new_n652), .B(new_n604), .C1(new_n378), .C2(new_n395), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n187), .B1(new_n608), .B2(new_n609), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n703), .A2(new_n704), .A3(new_n497), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NAND3_X1  g531(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n358), .A2(new_n365), .B1(new_n680), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT101), .B1(new_n719), .B2(new_n368), .ZN(new_n720));
  OAI22_X1  g534(.A1(new_n371), .A2(new_n373), .B1(new_n340), .B2(new_n386), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n722), .A3(new_n367), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n454), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n650), .A2(new_n725), .A3(KEYINPUT102), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n450), .B2(new_n454), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n724), .A2(new_n729), .A3(new_n625), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n703), .A2(new_n704), .A3(new_n686), .A4(new_n497), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n610), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NAND2_X1  g549(.A1(new_n551), .A2(new_n555), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n621), .A2(new_n611), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n736), .A2(new_n737), .A3(new_n659), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n724), .A2(new_n738), .A3(new_n625), .A4(new_n651), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n715), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  NAND2_X1  g556(.A1(new_n396), .A2(new_n455), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n188), .B1(new_n306), .B2(new_n310), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n507), .B1(new_n497), .B2(new_n502), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n746));
  AOI211_X1 g560(.A(KEYINPUT89), .B(new_n305), .C1(new_n289), .C2(new_n290), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n738), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n395), .B1(KEYINPUT32), .B2(new_n394), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n738), .A3(new_n729), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT42), .B1(new_n753), .B2(new_n748), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n322), .ZN(G33));
  NOR3_X1   g570(.A1(new_n743), .A2(new_n748), .A3(new_n664), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT103), .B(G134), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G36));
  NAND2_X1  g573(.A1(new_n309), .A2(new_n744), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n551), .A2(new_n555), .A3(new_n737), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n761), .A2(KEYINPUT106), .A3(new_n762), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n761), .A2(KEYINPUT105), .A3(new_n762), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT105), .B1(new_n761), .B2(new_n762), .ZN(new_n768));
  OAI22_X1  g582(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT107), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  OAI221_X1 g585(.A(new_n771), .B1(new_n767), .B2(new_n768), .C1(new_n765), .C2(new_n766), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n639), .A2(new_n651), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n760), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  INV_X1    g591(.A(new_n497), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n498), .A2(new_n499), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n499), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(G469), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n501), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n778), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n704), .ZN(new_n788));
  INV_X1    g602(.A(new_n676), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n777), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n787), .A2(KEYINPUT104), .A3(new_n704), .A4(new_n676), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n770), .A2(new_n772), .A3(KEYINPUT44), .A4(new_n773), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n776), .A2(new_n790), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n787), .A2(KEYINPUT47), .A3(new_n704), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n738), .B1(new_n454), .B2(new_n450), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n760), .A2(new_n396), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT108), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n798), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  NAND2_X1  g620(.A1(new_n703), .A2(new_n497), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT109), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n796), .B(new_n797), .C1(new_n509), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n311), .A2(new_n187), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n310), .B1(new_n301), .B2(KEYINPUT89), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(new_n308), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n730), .A2(new_n559), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n769), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n810), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  MUX2_X1   g631(.A(KEYINPUT116), .B(new_n817), .S(KEYINPUT51), .Z(new_n818));
  NOR3_X1   g632(.A1(new_n760), .A2(new_n559), .A3(new_n714), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n455), .A3(new_n685), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n736), .A3(new_n737), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n724), .A2(new_n625), .A3(new_n651), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n819), .A2(new_n769), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n714), .A2(new_n187), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n672), .A2(new_n674), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n672), .A2(KEYINPUT115), .A3(new_n674), .A4(new_n826), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n815), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(KEYINPUT50), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(KEYINPUT50), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n818), .B(new_n825), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n665), .A2(new_n668), .B1(new_n715), .B2(new_n740), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n659), .B(KEYINPUT112), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n648), .A2(new_n650), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n648), .A2(new_n650), .A3(new_n839), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n685), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n696), .A3(new_n686), .A4(new_n745), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n700), .A2(new_n835), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n700), .A2(new_n835), .A3(new_n843), .A4(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n664), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n599), .A2(new_n601), .A3(new_n659), .ZN(new_n850));
  INV_X1    g664(.A(new_n546), .ZN(new_n851));
  AOI211_X1 g665(.A(KEYINPUT20), .B(new_n851), .C1(new_n538), .C2(new_n544), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n555), .B(new_n850), .C1(new_n852), .C2(new_n547), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n633), .A2(KEYINPUT110), .A3(new_n555), .A4(new_n850), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n508), .B(new_n857), .C1(new_n497), .C2(new_n502), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n396), .A2(new_n858), .A3(new_n651), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n749), .A2(new_n849), .B1(new_n859), .B2(new_n813), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n813), .A2(new_n740), .A3(new_n861), .A4(new_n745), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT111), .B1(new_n748), .B2(new_n739), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n860), .A2(new_n864), .A3(new_n754), .A4(new_n751), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n736), .A2(new_n603), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n563), .B1(new_n866), .B2(new_n622), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n626), .A2(new_n867), .A3(new_n510), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n635), .A2(new_n706), .B1(new_n312), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n715), .A2(new_n712), .B1(new_n732), .B2(new_n733), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n312), .B(new_n605), .C1(new_n456), .C2(new_n653), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n707), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n848), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n848), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n848), .A2(new_n873), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n848), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n880));
  XNOR2_X1  g694(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n816), .A2(new_n715), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n557), .B(new_n883), .C1(new_n820), .C2(new_n623), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n824), .A2(new_n729), .A3(new_n752), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT48), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(KEYINPUT48), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n834), .A2(new_n876), .A3(new_n882), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n825), .B1(new_n833), .B2(new_n832), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT51), .B1(new_n892), .B2(new_n817), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n889), .A2(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  INV_X1    g708(.A(new_n675), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n729), .A2(new_n187), .A3(new_n509), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n761), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n685), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n809), .B2(KEYINPUT49), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n895), .B(new_n899), .C1(KEYINPUT49), .C2(new_n809), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n894), .A2(new_n900), .ZN(G75));
  OAI211_X1 g715(.A(G902), .B(new_n304), .C1(new_n874), .C2(new_n875), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n252), .A2(new_n254), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n286), .ZN(new_n904));
  XNOR2_X1  g718(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n904), .B(new_n905), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT119), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n908), .A2(KEYINPUT119), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n902), .A2(new_n907), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n283), .A2(G952), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n398), .B1(new_n879), .B2(new_n880), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n915), .B2(new_n304), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT118), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n902), .A2(new_n908), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n906), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n917), .B2(new_n920), .ZN(G51));
  XOR2_X1   g735(.A(new_n501), .B(KEYINPUT57), .Z(new_n922));
  AND3_X1   g736(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n495), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n783), .B(KEYINPUT121), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n912), .B1(new_n926), .B2(new_n928), .ZN(G54));
  NAND2_X1  g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n915), .A2(new_n545), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n545), .B1(new_n915), .B2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n912), .ZN(G60));
  NAND3_X1  g748(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT59), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n936), .B(new_n938), .C1(new_n923), .C2(new_n924), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n913), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n876), .A2(new_n882), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n936), .B1(new_n941), .B2(new_n938), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n879), .B2(new_n880), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT122), .B(new_n913), .C1(new_n946), .C2(new_n444), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n644), .A2(new_n647), .ZN(new_n948));
  INV_X1    g762(.A(new_n945), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n948), .B(new_n949), .C1(new_n874), .C2(new_n875), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n950), .B(new_n913), .C1(new_n946), .C2(new_n444), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n947), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n913), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n949), .B1(new_n874), .B2(new_n875), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n451), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n956), .B(new_n950), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(G224), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n560), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n872), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n903), .B1(G898), .B2(new_n283), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  NAND2_X1  g778(.A1(G900), .A2(G953), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n526), .A2(new_n527), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n352), .B(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n755), .A2(new_n757), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n696), .A2(new_n686), .A3(new_n729), .A4(new_n752), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n790), .A2(new_n791), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n700), .A2(new_n835), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n805), .A2(new_n793), .A3(new_n970), .A4(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n965), .B(new_n969), .C1(new_n975), .C2(G953), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n866), .A2(new_n622), .ZN(new_n977));
  OR4_X1    g791(.A1(new_n743), .A2(new_n760), .A3(new_n677), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n793), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n793), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n973), .A2(new_n689), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n973), .A2(KEYINPUT62), .A3(new_n689), .ZN(new_n987));
  AOI22_X1  g801(.A1(new_n986), .A2(new_n987), .B1(new_n804), .B2(new_n802), .ZN(new_n988));
  AOI21_X1  g802(.A(G953), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n969), .B(KEYINPUT125), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n976), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n975), .B2(new_n872), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n391), .A2(new_n680), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT127), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n912), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n356), .B1(new_n391), .B2(new_n340), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n995), .B(new_n1000), .C1(new_n874), .C2(new_n875), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n983), .A2(new_n988), .A3(new_n961), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n680), .B(new_n391), .C1(new_n1003), .C2(new_n995), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n1004), .ZN(G57));
endmodule


