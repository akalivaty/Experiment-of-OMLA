

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778;

  AND2_X1 U374 ( .A1(n514), .A2(n592), .ZN(n404) );
  XNOR2_X1 U375 ( .A(n501), .B(n379), .ZN(n763) );
  INV_X1 U376 ( .A(G953), .ZN(n765) );
  BUF_X1 U377 ( .A(n671), .Z(n351) );
  XNOR2_X2 U378 ( .A(G143), .B(G128), .ZN(n439) );
  XNOR2_X2 U379 ( .A(n425), .B(G125), .ZN(n444) );
  AND2_X1 U380 ( .A1(n418), .A2(n358), .ZN(n416) );
  NOR2_X1 U381 ( .A1(n628), .A2(n625), .ZN(n568) );
  XNOR2_X1 U382 ( .A(n548), .B(KEYINPUT99), .ZN(n776) );
  NAND2_X1 U383 ( .A1(n416), .A2(n413), .ZN(n548) );
  OR2_X1 U384 ( .A1(n585), .A2(n670), .ZN(n586) );
  XNOR2_X1 U385 ( .A(n374), .B(n528), .ZN(n532) );
  AND2_X1 U386 ( .A1(n369), .A2(n368), .ZN(n367) );
  XNOR2_X1 U387 ( .A(n440), .B(G131), .ZN(n486) );
  XNOR2_X1 U388 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n465) );
  XNOR2_X1 U389 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n464) );
  XNOR2_X2 U390 ( .A(n433), .B(n432), .ZN(n517) );
  INV_X1 U391 ( .A(G237), .ZN(n431) );
  XNOR2_X1 U392 ( .A(n444), .B(n390), .ZN(n761) );
  XNOR2_X1 U393 ( .A(G140), .B(KEYINPUT10), .ZN(n390) );
  NOR2_X1 U394 ( .A1(n776), .A2(n563), .ZN(n564) );
  NAND2_X1 U395 ( .A1(n570), .A2(KEYINPUT0), .ZN(n393) );
  NAND2_X1 U396 ( .A1(n402), .A2(n400), .ZN(n399) );
  NAND2_X1 U397 ( .A1(n401), .A2(n427), .ZN(n400) );
  NAND2_X1 U398 ( .A1(n395), .A2(n756), .ZN(n394) );
  NAND2_X1 U399 ( .A1(n397), .A2(n396), .ZN(n395) );
  NAND2_X1 U400 ( .A1(n426), .A2(n401), .ZN(n397) );
  NOR2_X1 U401 ( .A1(n582), .A2(n580), .ZN(n598) );
  NAND2_X2 U402 ( .A1(n367), .A2(n365), .ZN(n513) );
  OR2_X1 U403 ( .A1(n636), .A2(n366), .ZN(n365) );
  NAND2_X1 U404 ( .A1(G472), .A2(n443), .ZN(n366) );
  OR2_X2 U405 ( .A1(n570), .A2(n352), .ZN(n359) );
  XNOR2_X1 U406 ( .A(n363), .B(G107), .ZN(n754) );
  XNOR2_X1 U407 ( .A(G110), .B(G104), .ZN(n363) );
  XNOR2_X1 U408 ( .A(n364), .B(n754), .ZN(n438) );
  XNOR2_X1 U409 ( .A(n466), .B(KEYINPUT70), .ZN(n364) );
  XNOR2_X1 U410 ( .A(n454), .B(n453), .ZN(n703) );
  XOR2_X1 U411 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n482) );
  XNOR2_X1 U412 ( .A(n377), .B(n566), .ZN(n628) );
  NAND2_X1 U413 ( .A1(n524), .A2(KEYINPUT0), .ZN(n412) );
  INV_X1 U414 ( .A(G146), .ZN(n425) );
  XNOR2_X1 U415 ( .A(n486), .B(n441), .ZN(n379) );
  XNOR2_X1 U416 ( .A(KEYINPUT68), .B(G137), .ZN(n441) );
  INV_X1 U417 ( .A(G475), .ZN(n387) );
  XNOR2_X1 U418 ( .A(G113), .B(G116), .ZN(n421) );
  XNOR2_X1 U419 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X1 U420 ( .A(KEYINPUT24), .B(KEYINPUT73), .ZN(n409) );
  XNOR2_X1 U421 ( .A(G119), .B(G110), .ZN(n408) );
  XNOR2_X1 U422 ( .A(n446), .B(KEYINPUT23), .ZN(n410) );
  XNOR2_X1 U423 ( .A(G128), .B(G137), .ZN(n446) );
  XNOR2_X1 U424 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U425 ( .A(n485), .B(n388), .ZN(n491) );
  XNOR2_X1 U426 ( .A(n438), .B(n360), .ZN(n430) );
  XNOR2_X1 U427 ( .A(n361), .B(n439), .ZN(n360) );
  AND2_X1 U428 ( .A1(n592), .A2(n591), .ZN(n612) );
  NAND2_X1 U429 ( .A1(n525), .A2(KEYINPUT34), .ZN(n385) );
  NAND2_X1 U430 ( .A1(n370), .A2(n391), .ZN(n374) );
  AND2_X1 U431 ( .A1(n359), .A2(n598), .ZN(n370) );
  OR2_X1 U432 ( .A1(n703), .A2(n354), .ZN(n554) );
  OR2_X1 U433 ( .A1(n699), .A2(KEYINPUT83), .ZN(n417) );
  INV_X1 U434 ( .A(KEYINPUT83), .ZN(n414) );
  NAND2_X1 U435 ( .A1(n426), .A2(n444), .ZN(n402) );
  NOR2_X1 U436 ( .A1(n676), .A2(n673), .ZN(n693) );
  NAND2_X1 U437 ( .A1(n636), .A2(n473), .ZN(n369) );
  NAND2_X1 U438 ( .A1(n473), .A2(G902), .ZN(n368) );
  AND2_X1 U439 ( .A1(n621), .A2(n620), .ZN(n629) );
  INV_X1 U440 ( .A(KEYINPUT67), .ZN(n440) );
  XNOR2_X1 U441 ( .A(n761), .B(n389), .ZN(n388) );
  INV_X1 U442 ( .A(G113), .ZN(n389) );
  XOR2_X1 U443 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n483) );
  XNOR2_X1 U444 ( .A(G104), .B(G122), .ZN(n481) );
  XNOR2_X1 U445 ( .A(G902), .B(KEYINPUT15), .ZN(n625) );
  XNOR2_X1 U446 ( .A(n429), .B(n362), .ZN(n361) );
  XNOR2_X1 U447 ( .A(KEYINPUT74), .B(KEYINPUT17), .ZN(n362) );
  BUF_X1 U448 ( .A(n628), .Z(n749) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n457) );
  AND2_X1 U450 ( .A1(n393), .A2(n356), .ZN(n391) );
  INV_X1 U451 ( .A(n702), .ZN(n392) );
  NOR2_X1 U452 ( .A1(G237), .A2(G953), .ZN(n468) );
  XNOR2_X1 U453 ( .A(G122), .B(KEYINPUT97), .ZN(n494) );
  XOR2_X1 U454 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n495) );
  XNOR2_X1 U455 ( .A(n439), .B(G134), .ZN(n501) );
  XNOR2_X1 U456 ( .A(n504), .B(n375), .ZN(n580) );
  XNOR2_X1 U457 ( .A(n376), .B(KEYINPUT98), .ZN(n375) );
  INV_X1 U458 ( .A(G478), .ZN(n376) );
  INV_X1 U459 ( .A(KEYINPUT19), .ZN(n518) );
  NAND2_X1 U460 ( .A1(n517), .A2(n688), .ZN(n519) );
  XNOR2_X1 U461 ( .A(n492), .B(n386), .ZN(n582) );
  XNOR2_X1 U462 ( .A(n493), .B(n387), .ZN(n386) );
  XNOR2_X1 U463 ( .A(KEYINPUT16), .B(G122), .ZN(n424) );
  XNOR2_X1 U464 ( .A(n410), .B(n407), .ZN(n447) );
  XNOR2_X1 U465 ( .A(n436), .B(n435), .ZN(n437) );
  INV_X1 U466 ( .A(G140), .ZN(n435) );
  XNOR2_X1 U467 ( .A(n511), .B(n510), .ZN(n605) );
  OR2_X1 U468 ( .A1(n594), .A2(n699), .ZN(n679) );
  XNOR2_X1 U469 ( .A(n553), .B(KEYINPUT31), .ZN(n677) );
  NOR2_X1 U470 ( .A1(n582), .A2(n506), .ZN(n676) );
  NAND2_X1 U471 ( .A1(n415), .A2(n414), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n739), .B(n738), .ZN(n372) );
  OR2_X1 U473 ( .A1(n524), .A2(KEYINPUT0), .ZN(n352) );
  INV_X1 U474 ( .A(n406), .ZN(n699) );
  XNOR2_X1 U475 ( .A(n571), .B(KEYINPUT1), .ZN(n406) );
  AND2_X1 U476 ( .A1(n582), .A2(n580), .ZN(n353) );
  NAND2_X1 U477 ( .A1(n391), .A2(n359), .ZN(n354) );
  AND2_X1 U478 ( .A1(n393), .A2(n412), .ZN(n355) );
  AND2_X1 U479 ( .A1(n392), .A2(n412), .ZN(n356) );
  AND2_X1 U480 ( .A1(n385), .A2(n353), .ZN(n357) );
  AND2_X1 U481 ( .A1(n417), .A2(n547), .ZN(n358) );
  NAND2_X1 U482 ( .A1(n355), .A2(n359), .ZN(n525) );
  XNOR2_X2 U483 ( .A(n428), .B(G101), .ZN(n466) );
  XNOR2_X2 U484 ( .A(n513), .B(KEYINPUT6), .ZN(n592) );
  XNOR2_X2 U485 ( .A(n373), .B(n472), .ZN(n636) );
  NAND2_X1 U486 ( .A1(n371), .A2(n477), .ZN(n583) );
  XNOR2_X1 U487 ( .A(n476), .B(n475), .ZN(n371) );
  NOR2_X1 U488 ( .A1(n372), .A2(n745), .ZN(G63) );
  INV_X2 U489 ( .A(KEYINPUT4), .ZN(n428) );
  XNOR2_X2 U490 ( .A(n463), .B(n424), .ZN(n756) );
  XNOR2_X2 U491 ( .A(n423), .B(n422), .ZN(n463) );
  NAND2_X1 U492 ( .A1(n403), .A2(n399), .ZN(n398) );
  XNOR2_X1 U493 ( .A(n471), .B(n463), .ZN(n373) );
  NAND2_X1 U494 ( .A1(n406), .A2(n404), .ZN(n405) );
  NAND2_X1 U495 ( .A1(n398), .A2(n394), .ZN(n411) );
  NAND2_X1 U496 ( .A1(n564), .A2(n565), .ZN(n377) );
  XNOR2_X2 U497 ( .A(n519), .B(n518), .ZN(n570) );
  XNOR2_X1 U498 ( .A(n411), .B(n430), .ZN(n644) );
  XNOR2_X2 U499 ( .A(n378), .B(G469), .ZN(n571) );
  NAND2_X1 U500 ( .A1(n734), .A2(n443), .ZN(n378) );
  XNOR2_X2 U501 ( .A(n763), .B(G146), .ZN(n472) );
  NAND2_X1 U502 ( .A1(n723), .A2(KEYINPUT34), .ZN(n381) );
  XNOR2_X2 U503 ( .A(n405), .B(n516), .ZN(n723) );
  NOR2_X2 U504 ( .A1(n382), .A2(n380), .ZN(n527) );
  NAND2_X1 U505 ( .A1(n381), .A2(n357), .ZN(n380) );
  NOR2_X1 U506 ( .A1(n723), .A2(n383), .ZN(n382) );
  NAND2_X1 U507 ( .A1(n384), .A2(n526), .ZN(n383) );
  INV_X1 U508 ( .A(n525), .ZN(n384) );
  XNOR2_X2 U509 ( .A(n629), .B(KEYINPUT80), .ZN(n764) );
  NAND2_X1 U510 ( .A1(n444), .A2(n427), .ZN(n396) );
  INV_X1 U511 ( .A(n444), .ZN(n401) );
  INV_X1 U512 ( .A(n756), .ZN(n403) );
  INV_X1 U513 ( .A(n420), .ZN(n415) );
  NAND2_X1 U514 ( .A1(n420), .A2(n419), .ZN(n418) );
  AND2_X1 U515 ( .A1(n699), .A2(KEYINPUT83), .ZN(n419) );
  XNOR2_X1 U516 ( .A(n546), .B(KEYINPUT82), .ZN(n420) );
  XNOR2_X1 U517 ( .A(n568), .B(n567), .ZN(n622) );
  INV_X1 U518 ( .A(KEYINPUT79), .ZN(n567) );
  XNOR2_X1 U519 ( .A(n466), .B(n467), .ZN(n470) );
  NAND2_X1 U520 ( .A1(n609), .A2(n608), .ZN(n611) );
  XNOR2_X1 U521 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U522 ( .A(n438), .B(n437), .ZN(n442) );
  INV_X1 U523 ( .A(KEYINPUT34), .ZN(n526) );
  INV_X1 U524 ( .A(n421), .ZN(n423) );
  XNOR2_X1 U525 ( .A(KEYINPUT3), .B(G119), .ZN(n422) );
  XOR2_X1 U526 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n427) );
  INV_X1 U527 ( .A(n427), .ZN(n426) );
  NAND2_X1 U528 ( .A1(G224), .A2(n765), .ZN(n429) );
  NAND2_X1 U529 ( .A1(n644), .A2(n625), .ZN(n433) );
  INV_X1 U530 ( .A(G902), .ZN(n443) );
  NAND2_X1 U531 ( .A1(n443), .A2(n431), .ZN(n474) );
  AND2_X1 U532 ( .A1(n474), .A2(G210), .ZN(n432) );
  BUF_X1 U533 ( .A(n517), .Z(n615) );
  INV_X1 U534 ( .A(KEYINPUT38), .ZN(n434) );
  XNOR2_X1 U535 ( .A(n615), .B(n434), .ZN(n689) );
  NAND2_X1 U536 ( .A1(G227), .A2(n765), .ZN(n436) );
  XNOR2_X1 U537 ( .A(n442), .B(n472), .ZN(n734) );
  NAND2_X1 U538 ( .A1(G234), .A2(n765), .ZN(n445) );
  XOR2_X1 U539 ( .A(KEYINPUT8), .B(n445), .Z(n499) );
  NAND2_X1 U540 ( .A1(n499), .A2(G221), .ZN(n448) );
  XNOR2_X1 U541 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U542 ( .A(n761), .B(n449), .ZN(n741) );
  NOR2_X1 U543 ( .A1(n741), .A2(G902), .ZN(n454) );
  XOR2_X1 U544 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n452) );
  NAND2_X1 U545 ( .A1(n625), .A2(G234), .ZN(n450) );
  XNOR2_X1 U546 ( .A(n450), .B(KEYINPUT20), .ZN(n455) );
  NAND2_X1 U547 ( .A1(G217), .A2(n455), .ZN(n451) );
  XNOR2_X1 U548 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U549 ( .A1(G221), .A2(n455), .ZN(n456) );
  XNOR2_X1 U550 ( .A(n456), .B(KEYINPUT21), .ZN(n702) );
  OR2_X1 U551 ( .A1(n703), .A2(n702), .ZN(n709) );
  XNOR2_X1 U552 ( .A(n457), .B(KEYINPUT14), .ZN(n460) );
  NAND2_X1 U553 ( .A1(G902), .A2(n460), .ZN(n520) );
  NOR2_X1 U554 ( .A1(G900), .A2(n520), .ZN(n458) );
  NAND2_X1 U555 ( .A1(G953), .A2(n458), .ZN(n459) );
  XNOR2_X1 U556 ( .A(n459), .B(KEYINPUT101), .ZN(n461) );
  NAND2_X1 U557 ( .A1(G952), .A2(n460), .ZN(n720) );
  NOR2_X1 U558 ( .A1(n720), .A2(G953), .ZN(n522) );
  NOR2_X1 U559 ( .A1(n461), .A2(n522), .ZN(n572) );
  NOR2_X1 U560 ( .A1(n709), .A2(n572), .ZN(n462) );
  AND2_X1 U561 ( .A1(n571), .A2(n462), .ZN(n477) );
  XNOR2_X1 U562 ( .A(n465), .B(n464), .ZN(n467) );
  XNOR2_X1 U563 ( .A(KEYINPUT72), .B(n468), .ZN(n487) );
  NAND2_X1 U564 ( .A1(n487), .A2(G210), .ZN(n469) );
  INV_X1 U565 ( .A(G472), .ZN(n473) );
  BUF_X2 U566 ( .A(n513), .Z(n708) );
  INV_X1 U567 ( .A(n513), .ZN(n555) );
  NAND2_X1 U568 ( .A1(n474), .A2(G214), .ZN(n688) );
  NAND2_X1 U569 ( .A1(n555), .A2(n688), .ZN(n476) );
  XNOR2_X1 U570 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n475) );
  INV_X1 U571 ( .A(n583), .ZN(n478) );
  NAND2_X1 U572 ( .A1(n689), .A2(n478), .ZN(n480) );
  INV_X1 U573 ( .A(KEYINPUT39), .ZN(n479) );
  XNOR2_X1 U574 ( .A(n480), .B(n479), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U576 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U577 ( .A(G143), .B(n486), .ZN(n489) );
  NAND2_X1 U578 ( .A1(n487), .A2(G214), .ZN(n488) );
  XNOR2_X1 U579 ( .A(n491), .B(n490), .ZN(n654) );
  NOR2_X1 U580 ( .A1(G902), .A2(n654), .ZN(n492) );
  INV_X1 U581 ( .A(KEYINPUT13), .ZN(n493) );
  XNOR2_X1 U582 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U583 ( .A(n496), .B(KEYINPUT96), .Z(n498) );
  XNOR2_X1 U584 ( .A(G116), .B(G107), .ZN(n497) );
  XNOR2_X1 U585 ( .A(n498), .B(n497), .ZN(n503) );
  NAND2_X1 U586 ( .A1(G217), .A2(n499), .ZN(n500) );
  XOR2_X1 U587 ( .A(n501), .B(n500), .Z(n502) );
  XNOR2_X1 U588 ( .A(n503), .B(n502), .ZN(n738) );
  NOR2_X1 U589 ( .A1(G902), .A2(n738), .ZN(n504) );
  INV_X1 U590 ( .A(n580), .ZN(n506) );
  INV_X1 U591 ( .A(n676), .ZN(n505) );
  OR2_X1 U592 ( .A1(n508), .A2(n505), .ZN(n619) );
  XNOR2_X1 U593 ( .A(n619), .B(G134), .ZN(G36) );
  AND2_X1 U594 ( .A1(n582), .A2(n506), .ZN(n673) );
  INV_X1 U595 ( .A(n673), .ZN(n507) );
  OR2_X1 U596 ( .A1(n508), .A2(n507), .ZN(n511) );
  INV_X1 U597 ( .A(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U598 ( .A(n509), .B(KEYINPUT40), .ZN(n510) );
  XOR2_X1 U599 ( .A(G131), .B(KEYINPUT127), .Z(n512) );
  XNOR2_X1 U600 ( .A(n605), .B(n512), .ZN(G33) );
  INV_X1 U601 ( .A(n709), .ZN(n514) );
  XNOR2_X1 U602 ( .A(KEYINPUT100), .B(KEYINPUT33), .ZN(n515) );
  XNOR2_X1 U603 ( .A(n515), .B(KEYINPUT85), .ZN(n516) );
  XOR2_X1 U604 ( .A(G898), .B(KEYINPUT88), .Z(n748) );
  NAND2_X1 U605 ( .A1(G953), .A2(n748), .ZN(n758) );
  NOR2_X1 U606 ( .A1(n758), .A2(n520), .ZN(n521) );
  NOR2_X1 U607 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U608 ( .A(KEYINPUT89), .B(n523), .Z(n524) );
  XNOR2_X2 U609 ( .A(n527), .B(KEYINPUT35), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n541), .B(G122), .ZN(G24) );
  XNOR2_X1 U611 ( .A(n541), .B(KEYINPUT66), .ZN(n536) );
  XOR2_X1 U612 ( .A(KEYINPUT22), .B(KEYINPUT71), .Z(n528) );
  NOR2_X2 U613 ( .A1(n532), .A2(n592), .ZN(n546) );
  INV_X1 U614 ( .A(n703), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n699), .A2(n547), .ZN(n529) );
  NAND2_X1 U616 ( .A1(n546), .A2(n529), .ZN(n531) );
  INV_X1 U617 ( .A(KEYINPUT32), .ZN(n530) );
  XNOR2_X1 U618 ( .A(n531), .B(n530), .ZN(n777) );
  AND2_X1 U619 ( .A1(n708), .A2(n703), .ZN(n533) );
  NAND2_X1 U620 ( .A1(n699), .A2(n533), .ZN(n534) );
  NOR2_X1 U621 ( .A1(n532), .A2(n534), .ZN(n666) );
  NOR2_X1 U622 ( .A1(n777), .A2(n666), .ZN(n535) );
  NAND2_X1 U623 ( .A1(n536), .A2(n535), .ZN(n538) );
  INV_X1 U624 ( .A(KEYINPUT44), .ZN(n537) );
  NAND2_X1 U625 ( .A1(n538), .A2(n537), .ZN(n545) );
  NAND2_X1 U626 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n539) );
  OR2_X1 U627 ( .A1(n666), .A2(n539), .ZN(n540) );
  NOR2_X1 U628 ( .A1(n777), .A2(n540), .ZN(n543) );
  INV_X1 U629 ( .A(n541), .ZN(n549) );
  NAND2_X1 U630 ( .A1(n549), .A2(KEYINPUT84), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U632 ( .A1(n545), .A2(n544), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n549), .A2(KEYINPUT44), .ZN(n551) );
  INV_X1 U634 ( .A(KEYINPUT84), .ZN(n550) );
  NAND2_X1 U635 ( .A1(n551), .A2(n550), .ZN(n562) );
  NOR2_X1 U636 ( .A1(n554), .A2(n708), .ZN(n552) );
  NAND2_X1 U637 ( .A1(n406), .A2(n552), .ZN(n553) );
  INV_X1 U638 ( .A(n677), .ZN(n558) );
  NOR2_X1 U639 ( .A1(n555), .A2(n554), .ZN(n556) );
  AND2_X1 U640 ( .A1(n571), .A2(n556), .ZN(n662) );
  INV_X1 U641 ( .A(n662), .ZN(n557) );
  NAND2_X1 U642 ( .A1(n558), .A2(n557), .ZN(n560) );
  INV_X1 U643 ( .A(n693), .ZN(n559) );
  NAND2_X1 U644 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U645 ( .A1(n562), .A2(n561), .ZN(n563) );
  INV_X1 U646 ( .A(KEYINPUT45), .ZN(n566) );
  NAND2_X1 U647 ( .A1(n693), .A2(KEYINPUT47), .ZN(n569) );
  XOR2_X1 U648 ( .A(n569), .B(KEYINPUT77), .Z(n579) );
  XNOR2_X1 U649 ( .A(n571), .B(KEYINPUT104), .ZN(n576) );
  NOR2_X1 U650 ( .A1(n702), .A2(n572), .ZN(n573) );
  NAND2_X1 U651 ( .A1(n703), .A2(n573), .ZN(n588) );
  NOR2_X1 U652 ( .A1(n588), .A2(n708), .ZN(n574) );
  XNOR2_X1 U653 ( .A(n574), .B(KEYINPUT28), .ZN(n575) );
  NAND2_X1 U654 ( .A1(n576), .A2(n575), .ZN(n601) );
  NOR2_X1 U655 ( .A1(n570), .A2(n601), .ZN(n671) );
  INV_X1 U656 ( .A(n351), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n577), .A2(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n585) );
  AND2_X1 U659 ( .A1(n615), .A2(n580), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n584) );
  NOR2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n670) );
  XNOR2_X1 U662 ( .A(n586), .B(KEYINPUT76), .ZN(n597) );
  NOR2_X1 U663 ( .A1(KEYINPUT47), .A2(n693), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n587), .A2(n351), .ZN(n595) );
  INV_X1 U665 ( .A(n588), .ZN(n589) );
  AND2_X1 U666 ( .A1(n673), .A2(n589), .ZN(n590) );
  AND2_X1 U667 ( .A1(n688), .A2(n590), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n615), .A2(n612), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT36), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n679), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n609) );
  INV_X1 U672 ( .A(n598), .ZN(n691) );
  NAND2_X1 U673 ( .A1(n689), .A2(n688), .ZN(n692) );
  NOR2_X1 U674 ( .A1(n691), .A2(n692), .ZN(n600) );
  XNOR2_X1 U675 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n600), .B(n599), .ZN(n724) );
  OR2_X1 U677 ( .A1(n724), .A2(n601), .ZN(n604) );
  INV_X1 U678 ( .A(KEYINPUT107), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT42), .ZN(n603) );
  XNOR2_X1 U680 ( .A(n604), .B(n603), .ZN(n774) );
  NAND2_X1 U681 ( .A1(n774), .A2(n605), .ZN(n607) );
  INV_X1 U682 ( .A(KEYINPUT46), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(n621) );
  NAND2_X1 U686 ( .A1(n699), .A2(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(KEYINPUT43), .B(KEYINPUT102), .ZN(n613) );
  XNOR2_X1 U688 ( .A(n614), .B(n613), .ZN(n617) );
  INV_X1 U689 ( .A(n615), .ZN(n616) );
  AND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n682) );
  INV_X1 U691 ( .A(n682), .ZN(n618) );
  AND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n622), .A2(n764), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT78), .ZN(n627) );
  INV_X1 U695 ( .A(KEYINPUT2), .ZN(n624) );
  OR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n633) );
  INV_X1 U698 ( .A(n749), .ZN(n632) );
  NAND2_X1 U699 ( .A1(n629), .A2(KEYINPUT2), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT81), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n685) );
  AND2_X2 U702 ( .A1(n633), .A2(n685), .ZN(n731) );
  NAND2_X1 U703 ( .A1(n731), .A2(G472), .ZN(n638) );
  XOR2_X1 U704 ( .A(KEYINPUT86), .B(KEYINPUT108), .Z(n634) );
  XNOR2_X1 U705 ( .A(n634), .B(KEYINPUT62), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n638), .B(n637), .ZN(n642) );
  INV_X1 U708 ( .A(G952), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n639), .A2(G953), .ZN(n641) );
  INV_X1 U710 ( .A(KEYINPUT87), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n730) );
  NAND2_X1 U712 ( .A1(n642), .A2(n730), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U714 ( .A1(n731), .A2(G210), .ZN(n649) );
  BUF_X1 U715 ( .A(n644), .Z(n645) );
  XNOR2_X1 U716 ( .A(KEYINPUT117), .B(KEYINPUT54), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT55), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n645), .B(n647), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n650), .A2(n730), .ZN(n652) );
  INV_X1 U721 ( .A(KEYINPUT56), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(G51) );
  NAND2_X1 U723 ( .A1(n731), .A2(G475), .ZN(n656) );
  XNOR2_X1 U724 ( .A(KEYINPUT64), .B(KEYINPUT59), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n657), .A2(n730), .ZN(n660) );
  XOR2_X1 U728 ( .A(KEYINPUT119), .B(KEYINPUT60), .Z(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(KEYINPUT65), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G60) );
  NAND2_X1 U731 ( .A1(n662), .A2(n673), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n661), .B(G104), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n664) );
  NAND2_X1 U734 ( .A1(n662), .A2(n676), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(G107), .B(n665), .ZN(G9) );
  XOR2_X1 U737 ( .A(G110), .B(n666), .Z(G12) );
  XOR2_X1 U738 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n668) );
  NAND2_X1 U739 ( .A1(n351), .A2(n676), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U741 ( .A(G128), .B(n669), .Z(G30) );
  XOR2_X1 U742 ( .A(G143), .B(n670), .Z(G45) );
  NAND2_X1 U743 ( .A1(n351), .A2(n673), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n672), .B(G146), .ZN(G48) );
  NAND2_X1 U745 ( .A1(n677), .A2(n673), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT110), .ZN(n675) );
  XNOR2_X1 U747 ( .A(G113), .B(n675), .ZN(G15) );
  NAND2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n678), .B(G116), .ZN(G18) );
  XNOR2_X1 U750 ( .A(KEYINPUT37), .B(KEYINPUT111), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U752 ( .A(G125), .B(n681), .ZN(G27) );
  XOR2_X1 U753 ( .A(G140), .B(n682), .Z(G42) );
  INV_X1 U754 ( .A(n764), .ZN(n683) );
  NOR2_X1 U755 ( .A1(n749), .A2(n683), .ZN(n684) );
  NOR2_X1 U756 ( .A1(n684), .A2(KEYINPUT2), .ZN(n687) );
  INV_X1 U757 ( .A(n685), .ZN(n686) );
  NOR2_X1 U758 ( .A1(n687), .A2(n686), .ZN(n722) );
  NOR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U763 ( .A(n696), .B(KEYINPUT114), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n697), .A2(n723), .ZN(n698) );
  XOR2_X1 U765 ( .A(KEYINPUT115), .B(n698), .Z(n717) );
  XOR2_X1 U766 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n701) );
  NAND2_X1 U767 ( .A1(n699), .A2(n709), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n701), .B(n700), .ZN(n706) );
  AND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U770 ( .A(KEYINPUT49), .B(n704), .Z(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n707), .A2(n708), .ZN(n712) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n406), .A2(n710), .ZN(n711) );
  NAND2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U776 ( .A(KEYINPUT51), .B(n713), .ZN(n714) );
  NOR2_X1 U777 ( .A1(n724), .A2(n714), .ZN(n715) );
  XOR2_X1 U778 ( .A(KEYINPUT113), .B(n715), .Z(n716) );
  NOR2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U780 ( .A(n718), .B(KEYINPUT52), .ZN(n719) );
  NOR2_X1 U781 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n727) );
  NOR2_X1 U783 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U784 ( .A(KEYINPUT116), .B(n725), .Z(n726) );
  NAND2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U786 ( .A1(n728), .A2(G953), .ZN(n729) );
  XNOR2_X1 U787 ( .A(n729), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U788 ( .A(n730), .ZN(n745) );
  BUF_X2 U789 ( .A(n731), .Z(n740) );
  NAND2_X1 U790 ( .A1(n740), .A2(G469), .ZN(n736) );
  XOR2_X1 U791 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n732) );
  XOR2_X1 U792 ( .A(n732), .B(KEYINPUT118), .Z(n733) );
  XNOR2_X1 U793 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U794 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U795 ( .A1(n745), .A2(n737), .ZN(G54) );
  NAND2_X1 U796 ( .A1(n740), .A2(G478), .ZN(n739) );
  NAND2_X1 U797 ( .A1(n740), .A2(G217), .ZN(n743) );
  XNOR2_X1 U798 ( .A(n741), .B(KEYINPUT120), .ZN(n742) );
  XNOR2_X1 U799 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U800 ( .A1(n745), .A2(n744), .ZN(G66) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n746) );
  XOR2_X1 U802 ( .A(KEYINPUT61), .B(n746), .Z(n747) );
  NOR2_X1 U803 ( .A1(n748), .A2(n747), .ZN(n752) );
  NOR2_X1 U804 ( .A1(n749), .A2(G953), .ZN(n750) );
  XOR2_X1 U805 ( .A(KEYINPUT121), .B(n750), .Z(n751) );
  NOR2_X1 U806 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U807 ( .A(KEYINPUT122), .B(n753), .Z(n760) );
  XNOR2_X1 U808 ( .A(G101), .B(n754), .ZN(n755) );
  XNOR2_X1 U809 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U811 ( .A(n760), .B(n759), .Z(G69) );
  XNOR2_X1 U812 ( .A(n761), .B(KEYINPUT4), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(n767) );
  XNOR2_X1 U814 ( .A(n764), .B(n767), .ZN(n766) );
  NAND2_X1 U815 ( .A1(n766), .A2(n765), .ZN(n772) );
  XNOR2_X1 U816 ( .A(G227), .B(n767), .ZN(n768) );
  NAND2_X1 U817 ( .A1(n768), .A2(G900), .ZN(n769) );
  XNOR2_X1 U818 ( .A(KEYINPUT123), .B(n769), .ZN(n770) );
  NAND2_X1 U819 ( .A1(G953), .A2(n770), .ZN(n771) );
  NAND2_X1 U820 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U821 ( .A(KEYINPUT124), .B(n773), .Z(G72) );
  XNOR2_X1 U822 ( .A(G137), .B(n774), .ZN(n775) );
  XNOR2_X1 U823 ( .A(n775), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U824 ( .A(n776), .B(G101), .Z(G3) );
  XNOR2_X1 U825 ( .A(G119), .B(KEYINPUT125), .ZN(n778) );
  XNOR2_X1 U826 ( .A(n778), .B(n777), .ZN(G21) );
endmodule

