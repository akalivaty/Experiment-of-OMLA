//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT64), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  AND2_X1   g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G45), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n249), .A2(new_n208), .A3(G274), .A4(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n249), .A2(G226), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n217), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(G222), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(G223), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n262), .B(new_n263), .C1(new_n264), .C2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n256), .B1(new_n258), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G179), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n217), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G150), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n209), .A2(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G58), .A2(G68), .ZN(new_n281));
  INV_X1    g0081(.A(G50), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n209), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n275), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n274), .A2(new_n217), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n208), .A2(G20), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n285), .A2(G50), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n208), .A2(new_n282), .A3(G13), .A4(G20), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT65), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n286), .A2(new_n217), .A3(new_n274), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(G50), .ZN(new_n292));
  OAI211_X1 g0092(.A(KEYINPUT65), .B(new_n289), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n284), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n273), .B(new_n295), .C1(G169), .C2(new_n271), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n285), .A2(G77), .A3(new_n286), .A4(new_n287), .ZN(new_n297));
  INV_X1    g0097(.A(new_n286), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n264), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G20), .A2(G77), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n209), .A2(new_n266), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT15), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G87), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n301), .B1(new_n278), .B2(new_n302), .C1(new_n306), .C2(new_n279), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n300), .B1(new_n307), .B2(new_n275), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G244), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n254), .B1(new_n217), .B2(new_n257), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n253), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n269), .A2(G232), .A3(new_n259), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n269), .A2(G238), .A3(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G107), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n269), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n316), .B2(new_n258), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n309), .B1(new_n317), .B2(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n272), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n317), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G200), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n309), .B1(G190), .B2(new_n317), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT67), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT9), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n284), .B(new_n328), .C1(new_n290), .C2(new_n294), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n270), .A2(new_n258), .ZN(new_n332));
  INV_X1    g0132(.A(new_n256), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(G190), .B2(new_n271), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT66), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n330), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n335), .A3(KEYINPUT67), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n326), .A2(new_n337), .B1(new_n338), .B2(KEYINPUT10), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n337), .A2(new_n326), .A3(KEYINPUT10), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n296), .B(new_n325), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT68), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n326), .A3(KEYINPUT10), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n332), .A2(G190), .A3(new_n333), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n331), .B2(new_n271), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n327), .B2(new_n329), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT67), .B1(new_n347), .B2(new_n336), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n347), .B2(KEYINPUT67), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n344), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n351), .A2(KEYINPUT68), .A3(new_n296), .A4(new_n325), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n267), .A2(new_n209), .A3(new_n268), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n268), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n202), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(G20), .B1(new_n360), .B2(new_n281), .ZN(new_n361));
  INV_X1    g0161(.A(G159), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(new_n302), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n354), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n355), .A2(new_n365), .A3(new_n356), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G68), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n260), .A2(new_n261), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT7), .B1(new_n368), .B2(new_n209), .ZN(new_n369));
  INV_X1    g0169(.A(new_n358), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n367), .B1(new_n371), .B2(KEYINPUT72), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n209), .B1(new_n203), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n302), .A2(new_n362), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n361), .B(KEYINPUT73), .C1(new_n362), .C2(new_n302), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT16), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n275), .B(new_n364), .C1(new_n372), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n287), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n278), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n291), .B1(new_n382), .B2(KEYINPUT75), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n278), .B2(new_n381), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n383), .A2(new_n385), .B1(new_n298), .B2(new_n278), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(G223), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n388));
  OAI211_X1 g0188(.A(G226), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n388), .B(new_n389), .C1(new_n266), .C2(new_n222), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n258), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n249), .A2(G232), .A3(new_n254), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n253), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n253), .A2(KEYINPUT76), .A3(new_n392), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G169), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n253), .A2(new_n392), .A3(KEYINPUT76), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT76), .B1(new_n253), .B2(new_n392), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(G179), .A3(new_n391), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n387), .A2(KEYINPUT18), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT77), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT77), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n387), .A2(new_n406), .A3(new_n403), .A4(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n387), .A2(new_n403), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n401), .A2(G190), .A3(new_n391), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n397), .A2(G200), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n380), .A2(new_n386), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n331), .B1(new_n401), .B2(new_n391), .ZN(new_n417));
  AND4_X1   g0217(.A1(G190), .A2(new_n391), .A3(new_n395), .A4(new_n396), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n386), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT16), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n357), .A2(KEYINPUT72), .A3(new_n358), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(G68), .A3(new_n366), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n285), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n420), .B1(new_n424), .B2(new_n364), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(new_n425), .A3(KEYINPUT17), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n411), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT78), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n264), .B2(new_n279), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT71), .A3(new_n275), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT71), .B1(new_n431), .B2(new_n275), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT11), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n275), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT71), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT11), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n432), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n291), .A2(new_n202), .A3(new_n381), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT12), .B1(new_n286), .B2(G68), .ZN(new_n442));
  OR3_X1    g0242(.A1(new_n286), .A2(KEYINPUT12), .A3(G68), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n435), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT13), .ZN(new_n447));
  INV_X1    g0247(.A(new_n253), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n208), .A2(new_n252), .B1(new_n247), .B2(new_n248), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n221), .B1(new_n449), .B2(KEYINPUT69), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT69), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n311), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G232), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n454));
  OAI211_X1 g0254(.A(G226), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G97), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n258), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n447), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n249), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n452), .A2(G238), .A3(new_n460), .ZN(new_n461));
  AND4_X1   g0261(.A1(new_n447), .A2(new_n458), .A3(new_n253), .A4(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n446), .B(G169), .C1(new_n459), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n461), .A3(new_n253), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT13), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n453), .A2(new_n447), .A3(new_n458), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(G179), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n466), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n446), .B1(new_n469), .B2(G169), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n445), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n459), .A2(new_n462), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n445), .B1(new_n472), .B2(G190), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT70), .B1(new_n469), .B2(G200), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT70), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n331), .C1(new_n465), .C2(new_n466), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n416), .A2(new_n426), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT18), .B1(new_n387), .B2(new_n403), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(KEYINPUT77), .B2(new_n404), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(new_n407), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT78), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n353), .A2(new_n429), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n208), .A2(G33), .ZN(new_n487));
  AND4_X1   g0287(.A1(new_n217), .A2(new_n286), .A3(new_n274), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G97), .ZN(new_n489));
  INV_X1    g0289(.A(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n298), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  AND2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n205), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n315), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n371), .B2(new_n315), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n499), .B2(new_n275), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT79), .B1(new_n502), .B2(G41), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT79), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n250), .A3(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(G41), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n251), .A2(G1), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G257), .A3(new_n249), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n508), .A2(KEYINPUT80), .A3(G257), .A4(new_n249), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n249), .A2(G274), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(G244), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G250), .A2(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(KEYINPUT4), .A2(G244), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(G1698), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n269), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n515), .B1(new_n525), .B2(new_n258), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G169), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n513), .A2(new_n526), .A3(new_n272), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n501), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n532));
  OAI211_X1 g0332(.A(G238), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n533));
  INV_X1    g0333(.A(G116), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n266), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n258), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n208), .A2(G45), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT82), .A2(G250), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n258), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G274), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n507), .B(new_n540), .C1(KEYINPUT82), .C2(new_n223), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n303), .A2(new_n305), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n286), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n209), .B1(new_n456), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G87), .B2(new_n206), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n209), .B(G68), .C1(new_n260), .C2(new_n261), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n279), .B2(new_n490), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI221_X4 g0352(.A(new_n546), .B1(new_n488), .B2(G87), .C1(new_n552), .C2(new_n275), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n535), .A2(new_n258), .B1(new_n539), .B2(new_n541), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G190), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n544), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n275), .ZN(new_n557));
  INV_X1    g0357(.A(new_n546), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n488), .A2(new_n545), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n536), .A2(new_n272), .A3(new_n542), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(G169), .C2(new_n554), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G190), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n331), .B1(new_n513), .B2(new_n526), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  OAI221_X1 g0366(.A(new_n500), .B1(new_n527), .B2(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n531), .B(new_n563), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n571));
  OAI211_X1 g0371(.A(G257), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n267), .A2(G303), .A3(new_n268), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n574), .A2(new_n258), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n508), .A2(G270), .A3(new_n249), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n537), .B1(new_n502), .B2(G41), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n540), .B1(new_n247), .B2(new_n248), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n505), .A4(new_n503), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(KEYINPUT21), .B(G169), .C1(new_n575), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n574), .A2(new_n258), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(G179), .A3(new_n579), .A4(new_n576), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n298), .A2(new_n534), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n285), .A2(G116), .A3(new_n286), .A4(new_n487), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n274), .A2(new_n217), .B1(G20), .B2(new_n534), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n519), .B(new_n209), .C1(G33), .C2(new_n490), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n587), .A2(KEYINPUT20), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT20), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n585), .B(new_n586), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n582), .A2(new_n579), .A3(new_n576), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(new_n593), .B2(G200), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n564), .B2(new_n593), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n591), .B(G169), .C1(new_n575), .C2(new_n580), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT83), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n597), .B1(new_n596), .B2(new_n598), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n592), .B(new_n595), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n209), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n269), .A2(new_n604), .A3(new_n209), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT23), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n209), .B2(G107), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n315), .A2(KEYINPUT23), .A3(G20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(KEYINPUT84), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n612), .B1(new_n603), .B2(new_n605), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT24), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g0419(.A(KEYINPUT84), .B(new_n612), .C1(new_n603), .C2(new_n605), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n616), .B(new_n275), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n622));
  OAI211_X1 g0422(.A(G250), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n623));
  XOR2_X1   g0423(.A(KEYINPUT85), .B(G294), .Z(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n266), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n258), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n508), .A2(G264), .A3(new_n249), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n579), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n331), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n626), .A2(new_n564), .A3(new_n579), .A4(new_n627), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT25), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n286), .B2(G107), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n286), .A2(new_n632), .A3(G107), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n633), .A2(new_n635), .B1(new_n488), .B2(G107), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n621), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n636), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n617), .A2(new_n618), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(KEYINPUT24), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n617), .A2(new_n618), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n285), .B1(new_n642), .B2(new_n615), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n638), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n628), .A2(new_n528), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(G179), .B2(new_n628), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n637), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n570), .A2(new_n601), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n486), .A2(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n562), .ZN(new_n650));
  INV_X1    g0450(.A(new_n530), .ZN(new_n651));
  AOI21_X1  g0451(.A(G169), .B1(new_n513), .B2(new_n526), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n651), .A2(new_n652), .A3(new_n500), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n563), .A2(new_n653), .A3(KEYINPUT26), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n556), .A2(new_n562), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n531), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n650), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n592), .B1(new_n599), .B2(new_n600), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n644), .A2(new_n646), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n513), .A2(new_n526), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT81), .B1(new_n662), .B2(new_n331), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(G190), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n500), .A3(new_n568), .A4(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(new_n531), .A3(new_n563), .A4(new_n637), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n658), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n486), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT86), .Z(new_n669));
  NAND2_X1  g0469(.A1(new_n477), .A2(new_n321), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n479), .B1(new_n670), .B2(new_n471), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n528), .B1(new_n401), .B2(new_n391), .ZN(new_n672));
  AND4_X1   g0472(.A1(G179), .A2(new_n391), .A3(new_n395), .A4(new_n396), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n674), .A2(new_n425), .A3(new_n409), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n480), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT87), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT87), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n410), .A2(new_n404), .ZN(new_n679));
  INV_X1    g0479(.A(new_n470), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n467), .A3(new_n463), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n681), .A2(new_n445), .B1(new_n477), .B2(new_n321), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n678), .B(new_n679), .C1(new_n682), .C2(new_n479), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n677), .A2(new_n683), .A3(new_n351), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT88), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n296), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n684), .B2(new_n296), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n669), .B1(new_n687), .B2(new_n688), .ZN(G369));
  INV_X1    g0489(.A(new_n647), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n690), .B1(new_n644), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n621), .A2(new_n636), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n628), .A2(G179), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n528), .B2(new_n628), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n698), .B1(new_n702), .B2(new_n697), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n591), .A2(new_n696), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n659), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n601), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g0507(.A(KEYINPUT89), .B(G330), .Z(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT90), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT90), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n596), .A2(new_n598), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT83), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n696), .B1(new_n718), .B2(new_n592), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n690), .A2(new_n719), .B1(new_n660), .B2(new_n697), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n714), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n212), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n215), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n565), .A2(new_n566), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n527), .A2(new_n564), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n729), .A2(new_n501), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n653), .B1(new_n731), .B2(new_n568), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n702), .A2(new_n718), .A3(new_n592), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(new_n563), .A4(new_n637), .ZN(new_n734));
  AOI211_X1 g0534(.A(KEYINPUT29), .B(new_n696), .C1(new_n734), .C2(new_n658), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n667), .B2(new_n697), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n648), .A2(new_n697), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n543), .A2(new_n593), .A3(new_n272), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n527), .A2(new_n628), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT91), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n527), .A2(KEYINPUT91), .A3(new_n628), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n508), .A2(new_n249), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n747), .A2(G264), .B1(new_n625), .B2(new_n258), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(new_n513), .A3(new_n526), .A4(new_n554), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n746), .B1(new_n749), .B2(new_n583), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n554), .A2(new_n627), .A3(new_n626), .ZN(new_n751));
  INV_X1    g0551(.A(new_n583), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n662), .A2(new_n751), .A3(new_n752), .A4(KEYINPUT30), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n696), .B1(new_n745), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(KEYINPUT31), .B(new_n696), .C1(new_n745), .C2(new_n754), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n739), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n709), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n738), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n728), .B1(new_n761), .B2(G1), .ZN(G364));
  AND2_X1   g0562(.A1(new_n209), .A2(G13), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n208), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n723), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n217), .B1(G20), .B2(new_n528), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(G20), .A2(G179), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n564), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(KEYINPUT95), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(KEYINPUT95), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n771), .A2(G190), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n778), .A2(KEYINPUT94), .A3(new_n331), .ZN(new_n779));
  AOI21_X1  g0579(.A(KEYINPUT94), .B1(new_n778), .B2(new_n331), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n264), .B1(new_n201), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT96), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT98), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G179), .A2(G200), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G20), .A3(new_n564), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(G159), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n786), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n490), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n331), .A2(G179), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(G20), .A3(G190), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n222), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n793), .A2(new_n368), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n785), .A2(G159), .A3(new_n788), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n794), .A2(G20), .A3(new_n564), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT99), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n789), .B(new_n799), .C1(G107), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n778), .A2(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n772), .A2(new_n331), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n807), .A2(G50), .B1(G68), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n783), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n781), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G322), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n792), .A2(new_n624), .ZN(new_n813));
  INV_X1    g0613(.A(G329), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n368), .B1(new_n787), .B2(new_n814), .C1(new_n795), .C2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n813), .B(new_n816), .C1(new_n805), .C2(G283), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT33), .B(G317), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n808), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n807), .A2(G326), .B1(G311), .B2(new_n773), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n812), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n769), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n212), .A2(new_n269), .ZN(new_n823));
  INV_X1    g0623(.A(G355), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n824), .B1(G116), .B2(new_n212), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n722), .A2(new_n269), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n251), .B2(new_n216), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n242), .A2(new_n251), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n832));
  NOR2_X1   g0632(.A1(G13), .A2(G33), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n768), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n767), .B(new_n822), .C1(new_n831), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n835), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n707), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n710), .A2(new_n766), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n709), .B2(new_n707), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  AOI22_X1  g0645(.A1(new_n807), .A2(G137), .B1(G150), .B2(new_n808), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n781), .C1(new_n777), .C2(new_n362), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT34), .Z(new_n849));
  NAND2_X1  g0649(.A1(new_n805), .A2(G68), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n795), .A2(new_n282), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n368), .B(new_n851), .C1(G132), .C2(new_n788), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n852), .C1(new_n201), .C2(new_n792), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n807), .A2(G303), .B1(G283), .B2(new_n808), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n777), .B2(new_n534), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT100), .Z(new_n857));
  NAND2_X1  g0657(.A1(new_n805), .A2(G87), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n368), .B1(new_n795), .B2(new_n315), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n859), .B(new_n793), .C1(G311), .C2(new_n788), .ZN(new_n860));
  INV_X1    g0660(.A(G294), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n860), .C1(new_n781), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n768), .B1(new_n854), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n769), .A2(new_n834), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(G77), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n317), .A2(G190), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n323), .A2(new_n867), .A3(new_n308), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n309), .A2(new_n696), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n308), .B1(new_n322), .B2(new_n528), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n868), .A2(new_n869), .B1(new_n870), .B2(new_n319), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n318), .A2(new_n320), .A3(new_n696), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT101), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n321), .A2(new_n697), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT101), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n324), .A2(new_n323), .B1(new_n309), .B2(new_n696), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n321), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n834), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n766), .B1(new_n866), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n667), .A2(new_n697), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n760), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n767), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n882), .A2(new_n760), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(G384));
  OR2_X1    g0691(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n218), .A4(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT36), .Z(new_n895));
  NAND3_X1  g0695(.A1(new_n216), .A2(G77), .A3(new_n374), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n282), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n208), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n486), .A2(new_n759), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT104), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n445), .A2(new_n696), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n471), .A2(new_n477), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n471), .A2(new_n477), .A3(KEYINPUT103), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n468), .A2(new_n470), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n903), .B1(new_n477), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n759), .A3(new_n878), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n377), .A2(new_n378), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n423), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n354), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n420), .B1(new_n916), .B2(new_n424), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n414), .B1(new_n917), .B2(new_n694), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n674), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT37), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n694), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n387), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT37), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n408), .A2(new_n922), .A3(new_n923), .A4(new_n414), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n275), .B1(new_n372), .B2(new_n379), .ZN(new_n926));
  INV_X1    g0726(.A(new_n354), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n423), .B2(new_n914), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n386), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n921), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n925), .B1(new_n482), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n930), .B1(new_n411), .B2(new_n427), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n920), .B2(new_n924), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n931), .A2(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n902), .B1(new_n913), .B2(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n921), .A2(new_n929), .B1(new_n419), .B2(new_n425), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n403), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n923), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND4_X1   g0740(.A1(new_n923), .A2(new_n408), .A3(new_n922), .A4(new_n414), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT38), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n933), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n425), .A2(new_n694), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n676), .B2(new_n479), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n414), .B1(new_n425), .B2(new_n674), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT37), .B1(new_n946), .B2(new_n944), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n924), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT40), .B1(new_n943), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n937), .B1(new_n913), .B2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n901), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n901), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n709), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n666), .A2(new_n661), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT26), .B1(new_n563), .B2(new_n653), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n531), .A2(new_n656), .A3(new_n655), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n562), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n697), .B(new_n878), .C1(new_n955), .C2(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n959), .A2(new_n874), .B1(new_n908), .B2(new_n911), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n940), .A2(new_n941), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n932), .B1(new_n933), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n935), .B1(new_n482), .B2(new_n930), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n960), .A2(new_n964), .B1(new_n676), .B2(new_n694), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n943), .B2(new_n949), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n962), .A2(KEYINPUT39), .A3(new_n963), .ZN(new_n968));
  INV_X1    g0768(.A(new_n471), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n697), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n965), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n738), .A2(new_n485), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n684), .A2(new_n296), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT88), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n977), .B2(new_n686), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n974), .B(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n954), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT105), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n208), .B2(new_n763), .C1(new_n979), .C2(new_n954), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n980), .A2(KEYINPUT105), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n899), .B1(new_n982), .B2(new_n983), .ZN(G367));
  NOR2_X1   g0784(.A1(new_n792), .A2(new_n202), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n368), .B1(new_n788), .B2(G137), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n201), .B2(new_n795), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(new_n805), .C2(G77), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n807), .A2(G143), .B1(G159), .B2(new_n808), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(G150), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n282), .B2(new_n777), .C1(new_n991), .C2(new_n781), .ZN(new_n992));
  INV_X1    g0792(.A(new_n795), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT46), .B1(new_n993), .B2(G116), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n269), .B(new_n994), .C1(G317), .C2(new_n788), .ZN(new_n995));
  INV_X1    g0795(.A(new_n808), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(new_n315), .B2(new_n792), .C1(new_n996), .C2(new_n624), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n805), .A2(G97), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n993), .A2(KEYINPUT46), .A3(G116), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT110), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n999), .A2(new_n1000), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n997), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(G283), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n1005), .B2(new_n777), .ZN(new_n1006));
  INV_X1    g0806(.A(G311), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n807), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n781), .A2(new_n815), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT109), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n992), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n769), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n553), .A2(new_n697), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n656), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n650), .A2(new_n1015), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n835), .A3(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n238), .A2(new_n827), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n837), .B1(new_n722), .B2(new_n545), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n767), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n1014), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n531), .A2(new_n697), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT107), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n732), .B1(new_n500), .B2(new_n697), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n720), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT45), .Z(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n720), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT44), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(new_n714), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n690), .A2(new_n719), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n703), .B2(new_n719), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(new_n710), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n761), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT108), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1033), .A2(KEYINPUT108), .A3(new_n1038), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n761), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n723), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n765), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1027), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n714), .A2(KEYINPUT106), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT106), .B1(new_n714), .B2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n1051), .A2(KEYINPUT43), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(KEYINPUT43), .B2(new_n1052), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1048), .A2(new_n1034), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT42), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n531), .B1(new_n1048), .B2(new_n702), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n697), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1057), .A2(new_n1059), .B1(KEYINPUT43), .B2(new_n1052), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1055), .B(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1023), .B1(new_n1047), .B2(new_n1062), .ZN(G387));
  NAND2_X1  g0863(.A1(new_n1036), .A2(new_n765), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n792), .A2(new_n1005), .B1(new_n795), .B2(new_n624), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n807), .A2(G322), .B1(G311), .B2(new_n808), .ZN(new_n1066));
  INV_X1    g0866(.A(G317), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1066), .B1(new_n1067), .B2(new_n781), .C1(new_n777), .C2(new_n815), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT49), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n269), .B1(new_n788), .B2(G326), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n534), .C2(new_n804), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n791), .A2(new_n545), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n795), .A2(new_n264), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n368), .B(new_n1076), .C1(G150), .C2(new_n788), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n998), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n807), .A2(G159), .B1(G68), .B2(new_n773), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n278), .B2(new_n996), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(G50), .C2(new_n811), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT113), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n769), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n823), .A2(new_n725), .B1(G107), .B2(new_n212), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT111), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n234), .A2(new_n251), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n725), .ZN(new_n1087));
  AOI211_X1 g0887(.A(G45), .B(new_n1087), .C1(G68), .C2(G77), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n278), .A2(G50), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT50), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n827), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1085), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n766), .B1(new_n1092), .B2(new_n837), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT112), .Z(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n703), .B2(new_n840), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n723), .B(KEYINPUT114), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1037), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n761), .A2(new_n1036), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1064), .B1(new_n1083), .B2(new_n1095), .C1(new_n1097), .C2(new_n1098), .ZN(G393));
  NAND2_X1  g0899(.A1(new_n1033), .A2(new_n765), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n836), .B1(new_n490), .B2(new_n212), .C1(new_n827), .C2(new_n245), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n766), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n781), .A2(new_n1007), .B1(new_n1067), .B2(new_n1008), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT52), .Z(new_n1104));
  AOI22_X1  g0904(.A1(new_n808), .A2(G303), .B1(G116), .B2(new_n791), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1106), .A2(KEYINPUT115), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(KEYINPUT115), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n368), .B1(new_n795), .B2(new_n1005), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G322), .B2(new_n788), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n804), .B2(new_n315), .C1(new_n774), .C2(new_n861), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n781), .A2(new_n362), .B1(new_n991), .B2(new_n1008), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT51), .Z(new_n1114));
  NAND2_X1  g0914(.A1(new_n791), .A2(G77), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n269), .B1(new_n787), .B2(new_n847), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G68), .B2(new_n993), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n858), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G50), .B2(new_n808), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n278), .B2(new_n777), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1104), .A2(new_n1112), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1102), .B1(new_n1121), .B2(new_n768), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n840), .B2(new_n1027), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1100), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1096), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1124), .B1(new_n1043), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G390));
  INV_X1    g0929(.A(new_n968), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n947), .A2(new_n924), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n922), .B1(new_n427), .B2(new_n679), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n932), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT39), .B1(new_n1133), .B2(new_n963), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1130), .A2(new_n1134), .B1(new_n971), .B2(new_n960), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n959), .A2(new_n874), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n912), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n970), .C1(new_n943), .C2(new_n949), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n757), .A2(new_n758), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n570), .A2(new_n647), .A3(new_n601), .A4(new_n696), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n878), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n910), .B1(new_n906), .B2(new_n907), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n709), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1135), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(G330), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n913), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n759), .A2(new_n709), .A3(new_n878), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1142), .A2(new_n959), .A3(new_n874), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1137), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1142), .A2(new_n959), .A3(new_n874), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n960), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n759), .A2(G330), .A3(new_n878), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n484), .A2(new_n429), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1159), .A2(G330), .A3(new_n353), .A4(new_n759), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n978), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1126), .B1(new_n1151), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1145), .B1(new_n1164), .B2(new_n1149), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1161), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1151), .A2(new_n765), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n834), .B1(new_n967), .B2(new_n968), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n807), .A2(G283), .B1(G107), .B2(new_n808), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n269), .B(new_n796), .C1(G294), .C2(new_n788), .ZN(new_n1171));
  AND4_X1   g0971(.A1(new_n850), .A2(new_n1170), .A3(new_n1115), .A4(new_n1171), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n490), .B2(new_n777), .C1(new_n534), .C2(new_n781), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n795), .A2(new_n991), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT53), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n368), .B1(new_n788), .B2(G125), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n362), .C2(new_n792), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G50), .B2(new_n805), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n811), .A2(G132), .ZN(new_n1179));
  XOR2_X1   g0979(.A(KEYINPUT54), .B(G143), .Z(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n775), .B2(new_n776), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n807), .A2(G128), .B1(G137), .B2(new_n808), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n769), .B1(new_n1173), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n278), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n766), .B1(new_n1185), .B2(new_n865), .ZN(new_n1186));
  OR3_X1    g0986(.A1(new_n1169), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1167), .A2(new_n1168), .A3(new_n1187), .ZN(G378));
  OAI21_X1  g0988(.A(new_n766), .B1(G50), .B2(new_n865), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n269), .A2(G41), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G50), .B(new_n1190), .C1(new_n266), .C2(new_n250), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1008), .A2(new_n534), .B1(new_n306), .B2(new_n774), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G97), .B2(new_n808), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n804), .A2(new_n201), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1190), .B1(new_n1005), .B2(new_n787), .C1(new_n264), .C2(new_n795), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1194), .A2(new_n985), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(new_n315), .C2(new_n781), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1191), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n792), .A2(new_n991), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n993), .A2(new_n1180), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT116), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G137), .C2(new_n773), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n807), .A2(G125), .B1(G132), .B2(new_n808), .ZN(new_n1204));
  INV_X1    g1004(.A(G128), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1204), .C1(new_n1205), .C2(new_n781), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n362), .C2(new_n804), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(new_n1198), .B2(new_n1197), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1189), .B1(new_n1211), .B2(new_n768), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n351), .A2(new_n296), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n295), .A2(new_n921), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n351), .A2(new_n296), .A3(new_n1214), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1212), .B1(new_n1222), .B2(new_n834), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(G330), .B1(new_n913), .B2(new_n950), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT40), .B1(new_n1143), .B2(new_n964), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1222), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n902), .B1(new_n1133), .B2(new_n963), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1147), .B1(new_n1143), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n937), .A2(new_n1229), .A3(new_n1221), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n973), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT117), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1227), .A2(new_n1230), .A3(KEYINPUT117), .A4(new_n973), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT118), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(new_n974), .ZN(new_n1237));
  AOI211_X1 g1037(.A(KEYINPUT118), .B(new_n973), .C1(new_n1227), .C2(new_n1230), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1233), .B(new_n1234), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1224), .B1(new_n1239), .B2(new_n765), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1157), .B1(new_n1137), .B2(new_n1153), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1156), .B2(new_n1152), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n978), .B(new_n1160), .C1(new_n1165), .C2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1236), .A2(new_n974), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1231), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT57), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1159), .B(new_n353), .C1(new_n737), .C2(new_n735), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1160), .B(new_n1248), .C1(new_n687), .C2(new_n688), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1151), .B2(new_n1162), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1096), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1240), .B1(new_n1244), .B2(new_n1251), .ZN(G375));
  XNOR2_X1  g1052(.A(new_n1249), .B(new_n1158), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1046), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n807), .A2(G294), .B1(G116), .B2(new_n808), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n777), .B2(new_n315), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT119), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1075), .B1(new_n490), .B2(new_n795), .C1(new_n815), .C2(new_n787), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n368), .B1(new_n804), .B2(new_n264), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT120), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G283), .C2(new_n811), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n807), .A2(G132), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT121), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n269), .B1(new_n787), .B2(new_n1205), .C1(new_n795), .C2(new_n362), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1264), .B(new_n1194), .C1(G50), .C2(new_n791), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G150), .A2(new_n773), .B1(new_n808), .B2(new_n1180), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G137), .B2(new_n811), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1257), .A2(new_n1261), .B1(new_n1263), .B2(new_n1268), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n766), .B1(G68), .B2(new_n865), .C1(new_n1269), .C2(new_n769), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n833), .B2(new_n1142), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1158), .B2(new_n765), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1254), .A2(new_n1272), .ZN(G381));
  NOR3_X1   g1073(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1128), .A2(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(G387), .A2(G381), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1168), .A2(new_n1187), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1278));
  INV_X1    g1078(.A(G375), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .ZN(G407));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(G343), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1278), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(G213), .A3(new_n1283), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT122), .Z(G409));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1240), .C1(new_n1244), .C2(new_n1251), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1046), .B(new_n1243), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1224), .B1(new_n1246), .B2(new_n765), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1278), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1282), .B1(new_n1287), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1158), .B1(new_n978), .B2(new_n1160), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1096), .B1(new_n1295), .B2(KEYINPUT60), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1242), .A2(new_n1249), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1298), .B2(new_n1161), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1272), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n888), .A2(KEYINPUT123), .A3(new_n889), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT123), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n889), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n887), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1126), .B1(new_n1298), .B2(new_n1297), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1253), .B2(new_n1297), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1307), .A2(new_n890), .A3(new_n1302), .A4(new_n1272), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1282), .A2(G2897), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1305), .A2(new_n1308), .A3(G2897), .A4(new_n1282), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1286), .B1(new_n1294), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(KEYINPUT125), .B(new_n1286), .C1(new_n1294), .C2(new_n1313), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1287), .A2(new_n1293), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1282), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1309), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1319), .B1(new_n1322), .B2(KEYINPUT126), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1294), .A2(new_n1309), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(KEYINPUT62), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT127), .B1(new_n1318), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT127), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1323), .A4(new_n1326), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1055), .B(new_n1060), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n761), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1333), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n764), .B1(new_n1334), .B2(new_n1045), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1022), .B1(new_n1332), .B2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT124), .B1(new_n1336), .B2(G390), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(G393), .B(new_n844), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1336), .A2(G390), .ZN(new_n1340));
  AOI211_X1 g1140(.A(new_n1022), .B(new_n1128), .C1(new_n1332), .C2(new_n1335), .ZN(new_n1341));
  OAI22_X1  g1141(.A1(new_n1337), .A2(new_n1339), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G387), .A2(new_n1128), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1336), .A2(G390), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1343), .A2(KEYINPUT124), .A3(new_n1344), .A4(new_n1338), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1328), .A2(new_n1331), .A3(new_n1346), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1322), .B(KEYINPUT63), .ZN(new_n1348));
  OR3_X1    g1148(.A1(new_n1348), .A2(new_n1346), .A3(new_n1314), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(G405));
  INV_X1    g1150(.A(new_n1309), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1346), .A2(new_n1351), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(G375), .B(G378), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1342), .A2(new_n1309), .A3(new_n1345), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1353), .B1(new_n1352), .B2(new_n1354), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1356), .ZN(G402));
endmodule


