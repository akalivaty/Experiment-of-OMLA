

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U322 ( .A(n358), .B(n292), .ZN(n359) );
  XNOR2_X1 U323 ( .A(n411), .B(n290), .ZN(n569) );
  XNOR2_X1 U324 ( .A(n328), .B(n291), .ZN(n329) );
  XNOR2_X1 U325 ( .A(n364), .B(n363), .ZN(n553) );
  XNOR2_X1 U326 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U327 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U328 ( .A(KEYINPUT117), .B(KEYINPUT54), .ZN(n290) );
  XOR2_X1 U329 ( .A(n327), .B(n326), .Z(n291) );
  AND2_X1 U330 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U331 ( .A(n320), .B(KEYINPUT72), .Z(n293) );
  XNOR2_X1 U332 ( .A(n389), .B(KEYINPUT46), .ZN(n390) );
  NOR2_X1 U333 ( .A1(n391), .A2(n553), .ZN(n392) );
  XNOR2_X1 U334 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n313) );
  XOR2_X1 U335 ( .A(G92GAT), .B(G85GAT), .Z(n353) );
  XNOR2_X1 U336 ( .A(n313), .B(KEYINPUT69), .ZN(n376) );
  XOR2_X1 U337 ( .A(KEYINPUT36), .B(n553), .Z(n583) );
  XNOR2_X1 U338 ( .A(n330), .B(n329), .ZN(n576) );
  NOR2_X1 U339 ( .A1(n530), .A2(n450), .ZN(n565) );
  XOR2_X1 U340 ( .A(n445), .B(n444), .Z(n525) );
  XNOR2_X1 U341 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U342 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n294), .B(KEYINPUT88), .ZN(n295) );
  XOR2_X1 U345 ( .A(n295), .B(KEYINPUT18), .Z(n297) );
  XNOR2_X1 U346 ( .A(G183GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n405) );
  XOR2_X1 U348 ( .A(G113GAT), .B(G15GAT), .Z(n334) );
  XOR2_X1 U349 ( .A(G176GAT), .B(KEYINPUT86), .Z(n299) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n334), .B(n300), .Z(n302) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U355 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n304) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(KEYINPUT87), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(n306), .B(n305), .Z(n311) );
  XNOR2_X1 U359 ( .A(G99GAT), .B(G71GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n307), .B(G120GAT), .ZN(n321) );
  XOR2_X1 U361 ( .A(G127GAT), .B(KEYINPUT0), .Z(n309) );
  XNOR2_X1 U362 ( .A(G134GAT), .B(KEYINPUT83), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n437) );
  XNOR2_X1 U364 ( .A(n321), .B(n437), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n405), .B(n312), .ZN(n530) );
  XOR2_X1 U367 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n448) );
  INV_X1 U368 ( .A(n353), .ZN(n314) );
  NAND2_X1 U369 ( .A1(n376), .A2(n314), .ZN(n317) );
  INV_X1 U370 ( .A(n376), .ZN(n315) );
  NAND2_X1 U371 ( .A1(n315), .A2(n353), .ZN(n316) );
  NAND2_X1 U372 ( .A1(n317), .A2(n316), .ZN(n319) );
  NAND2_X1 U373 ( .A1(G230GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(KEYINPUT32), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n293), .B(n322), .ZN(n330) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G78GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n323), .B(G148GAT), .ZN(n418) );
  XOR2_X1 U379 ( .A(G64GAT), .B(KEYINPUT73), .Z(n325) );
  XNOR2_X1 U380 ( .A(G176GAT), .B(G204GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n400) );
  XNOR2_X1 U382 ( .A(n418), .B(n400), .ZN(n328) );
  XOR2_X1 U383 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n327) );
  XNOR2_X1 U384 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n326) );
  XOR2_X1 U385 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n332) );
  XNOR2_X1 U386 ( .A(KEYINPUT65), .B(KEYINPUT30), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n341) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n333), .B(G8GAT), .ZN(n401) );
  XOR2_X1 U390 ( .A(n334), .B(n401), .Z(n336) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n337), .B(G1GAT), .Z(n339) );
  XOR2_X1 U394 ( .A(G141GAT), .B(G22GAT), .Z(n415) );
  XNOR2_X1 U395 ( .A(n415), .B(G197GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n346) );
  XOR2_X1 U398 ( .A(G29GAT), .B(KEYINPUT66), .Z(n343) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G43GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n345) );
  XOR2_X1 U401 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n364) );
  XOR2_X1 U403 ( .A(n346), .B(n364), .Z(n502) );
  INV_X1 U404 ( .A(n502), .ZN(n572) );
  XNOR2_X1 U405 ( .A(KEYINPUT68), .B(n572), .ZN(n556) );
  XOR2_X1 U406 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n348) );
  XNOR2_X1 U407 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n350) );
  XNOR2_X1 U410 ( .A(G99GAT), .B(KEYINPUT64), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n362) );
  XOR2_X1 U413 ( .A(n353), .B(G218GAT), .Z(n355) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(G134GAT), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n357) );
  XNOR2_X1 U417 ( .A(G190GAT), .B(G162GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U420 ( .A(G78GAT), .B(G211GAT), .Z(n366) );
  XNOR2_X1 U421 ( .A(G22GAT), .B(G155GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U423 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n368) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(G64GAT), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U426 ( .A(n370), .B(n369), .Z(n375) );
  XOR2_X1 U427 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n372) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U430 ( .A(KEYINPUT79), .B(n373), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U432 ( .A(n376), .B(G127GAT), .Z(n378) );
  XNOR2_X1 U433 ( .A(G183GAT), .B(G71GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U435 ( .A(n380), .B(n379), .Z(n385) );
  XOR2_X1 U436 ( .A(KEYINPUT12), .B(KEYINPUT82), .Z(n382) );
  XNOR2_X1 U437 ( .A(G1GAT), .B(KEYINPUT81), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U439 ( .A(G15GAT), .B(n383), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n535) );
  NOR2_X1 U441 ( .A1(n583), .A2(n535), .ZN(n386) );
  XOR2_X1 U442 ( .A(KEYINPUT45), .B(n386), .Z(n387) );
  NOR2_X1 U443 ( .A1(n556), .A2(n387), .ZN(n388) );
  NAND2_X1 U444 ( .A1(n576), .A2(n388), .ZN(n395) );
  XNOR2_X1 U445 ( .A(KEYINPUT110), .B(KEYINPUT47), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n576), .B(KEYINPUT41), .ZN(n549) );
  NAND2_X1 U447 ( .A1(n549), .A2(n572), .ZN(n389) );
  NAND2_X1 U448 ( .A1(n390), .A2(n535), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n394) );
  NAND2_X1 U450 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n396), .B(KEYINPUT48), .ZN(n524) );
  XOR2_X1 U452 ( .A(KEYINPUT78), .B(KEYINPUT94), .Z(n398) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(n399), .B(G92GAT), .Z(n403) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n410) );
  XOR2_X1 U459 ( .A(KEYINPUT90), .B(G218GAT), .Z(n407) );
  XNOR2_X1 U460 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U462 ( .A(G197GAT), .B(n408), .Z(n426) );
  INV_X1 U463 ( .A(n426), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n516) );
  NAND2_X1 U465 ( .A1(n524), .A2(n516), .ZN(n411) );
  XOR2_X1 U466 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n413) );
  XNOR2_X1 U467 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U469 ( .A(n414), .B(KEYINPUT24), .Z(n417) );
  XNOR2_X1 U470 ( .A(G50GAT), .B(n415), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U472 ( .A(n418), .B(G204GAT), .Z(n420) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U475 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U476 ( .A(KEYINPUT2), .B(G162GAT), .Z(n424) );
  XNOR2_X1 U477 ( .A(KEYINPUT91), .B(G155GAT), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(KEYINPUT3), .B(n425), .Z(n441) );
  XNOR2_X1 U480 ( .A(n441), .B(n426), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n463) );
  XOR2_X1 U482 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n430) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n445) );
  XOR2_X1 U485 ( .A(KEYINPUT75), .B(G85GAT), .Z(n432) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(G120GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U488 ( .A(G57GAT), .B(G148GAT), .Z(n434) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(G113GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U491 ( .A(n436), .B(n435), .Z(n443) );
  XOR2_X1 U492 ( .A(n437), .B(KEYINPUT5), .Z(n439) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  INV_X1 U497 ( .A(n525), .ZN(n568) );
  AND2_X1 U498 ( .A1(n463), .A2(n568), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n569), .A2(n446), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT55), .B(n449), .Z(n450) );
  NAND2_X1 U502 ( .A1(n565), .A2(n553), .ZN(n454) );
  XOR2_X1 U503 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n452) );
  XNOR2_X1 U504 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n451) );
  NAND2_X1 U505 ( .A1(n556), .A2(n576), .ZN(n488) );
  NOR2_X1 U506 ( .A1(n553), .A2(n535), .ZN(n455) );
  XNOR2_X1 U507 ( .A(KEYINPUT16), .B(n455), .ZN(n473) );
  XNOR2_X1 U508 ( .A(n463), .B(KEYINPUT28), .ZN(n528) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(n516), .ZN(n527) );
  XNOR2_X1 U511 ( .A(KEYINPUT89), .B(n530), .ZN(n457) );
  NOR2_X1 U512 ( .A1(n527), .A2(n457), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n528), .A2(n458), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n459), .A2(n525), .ZN(n471) );
  INV_X1 U515 ( .A(n530), .ZN(n518) );
  NAND2_X1 U516 ( .A1(n516), .A2(n518), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n460), .A2(n463), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(KEYINPUT97), .ZN(n462) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(n462), .ZN(n469) );
  NOR2_X1 U520 ( .A1(n518), .A2(n463), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n465), .B(n464), .ZN(n570) );
  INV_X1 U523 ( .A(n570), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n466), .A2(n527), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n525), .A2(n467), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n485) );
  INV_X1 U528 ( .A(n485), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n504) );
  NOR2_X1 U530 ( .A1(n488), .A2(n504), .ZN(n483) );
  NAND2_X1 U531 ( .A1(n483), .A2(n525), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n516), .A2(n483), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT98), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n479) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n483), .A2(n518), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT99), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  INV_X1 U543 ( .A(n528), .ZN(n520) );
  NAND2_X1 U544 ( .A1(n483), .A2(n520), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n492) );
  NOR2_X1 U547 ( .A1(n583), .A2(n485), .ZN(n486) );
  NAND2_X1 U548 ( .A1(n486), .A2(n535), .ZN(n487) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n487), .Z(n513) );
  NOR2_X1 U550 ( .A1(n513), .A2(n488), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n499) );
  NAND2_X1 U553 ( .A1(n499), .A2(n525), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U555 ( .A(G29GAT), .B(n493), .Z(G1328GAT) );
  NAND2_X1 U556 ( .A1(n516), .A2(n499), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U560 ( .A1(n499), .A2(n518), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n501) );
  NAND2_X1 U564 ( .A1(n520), .A2(n499), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  XOR2_X1 U567 ( .A(KEYINPUT107), .B(n549), .Z(n560) );
  NAND2_X1 U568 ( .A1(n560), .A2(n502), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(KEYINPUT108), .ZN(n514) );
  NOR2_X1 U570 ( .A1(n514), .A2(n504), .ZN(n510) );
  NAND2_X1 U571 ( .A1(n525), .A2(n510), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n516), .A2(n510), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT109), .Z(n509) );
  NAND2_X1 U576 ( .A1(n510), .A2(n518), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U579 ( .A1(n510), .A2(n520), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n525), .A2(n521), .ZN(n515) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n516), .A2(n521), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n525), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n542), .A2(n528), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n538), .A2(n556), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT111), .Z(n533) );
  NAND2_X1 U598 ( .A1(n538), .A2(n560), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  INV_X1 U601 ( .A(n535), .ZN(n580) );
  NAND2_X1 U602 ( .A1(n580), .A2(n538), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT112), .Z(n540) );
  NAND2_X1 U606 ( .A1(n538), .A2(n553), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n541), .ZN(G1343GAT) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT114), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n570), .A2(n542), .ZN(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT113), .B(n543), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n554), .A2(n572), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U617 ( .A(KEYINPUT115), .B(n548), .Z(n551) );
  NAND2_X1 U618 ( .A1(n554), .A2(n549), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n580), .A2(n554), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n565), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n557) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XNOR2_X1 U627 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n564) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .Z(n562) );
  NAND2_X1 U629 ( .A1(n565), .A2(n560), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .Z(n567) );
  NAND2_X1 U633 ( .A1(n565), .A2(n580), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  AND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n582) );
  INV_X1 U638 ( .A(n582), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  OR2_X1 U643 ( .A1(n582), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

