//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(new_n202), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n209), .A2(new_n213), .A3(new_n221), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n227), .B(new_n230), .Z(G358));
  XOR2_X1   g0031(.A(G87), .B(G97), .Z(new_n232));
  XNOR2_X1  g0032(.A(G107), .B(G116), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(G50), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(G68), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n234), .B(new_n241), .ZN(G351));
  OR2_X1    g0042(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g0043(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n243), .A2(G33), .A3(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT73), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT73), .A2(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(KEYINPUT3), .A3(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n245), .A2(new_n250), .A3(new_n211), .A4(G68), .ZN(new_n251));
  NAND3_X1  g0051(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n211), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT84), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G97), .A2(G107), .ZN(new_n255));
  INV_X1    g0055(.A(G87), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT84), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n252), .A2(new_n258), .A3(new_n211), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT19), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n211), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G97), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n251), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n212), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT15), .B(G87), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT68), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n211), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n269), .B(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n273), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n267), .B(KEYINPUT67), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n247), .A2(G1), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n276), .A2(new_n277), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n268), .A2(new_n274), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT85), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n265), .A2(new_n267), .B1(new_n273), .B2(new_n270), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(KEYINPUT85), .A3(new_n281), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n271), .A2(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G250), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(G274), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT83), .B1(new_n293), .B2(new_n290), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  AND2_X1   g0095(.A1(G1), .A2(G13), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n287), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT83), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n292), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G238), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G244), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G1698), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n245), .A2(new_n250), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n248), .A2(new_n249), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G116), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(G179), .B(new_n302), .C1(new_n311), .C2(new_n288), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n298), .B1(new_n297), .B2(new_n300), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n289), .B2(new_n291), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n288), .B1(new_n308), .B2(new_n310), .ZN(new_n316));
  OAI21_X1  g0116(.A(G169), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n284), .A2(new_n286), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n315), .A2(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G190), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n266), .A2(new_n212), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n266), .A2(KEYINPUT67), .A3(new_n212), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n323), .A2(new_n273), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n280), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G87), .ZN(new_n328));
  OAI21_X1  g0128(.A(G200), .B1(new_n315), .B2(new_n316), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n321), .A2(new_n328), .A3(new_n285), .A4(new_n329), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n319), .A2(KEYINPUT86), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT86), .B1(new_n319), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G41), .ZN(new_n334));
  AOI21_X1  g0134(.A(G1), .B1(new_n334), .B2(new_n299), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n288), .A3(G274), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n288), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(G226), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G33), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(G222), .A3(new_n304), .ZN(new_n346));
  INV_X1    g0146(.A(G77), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(G1698), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT66), .B(G223), .Z(new_n349));
  OAI221_X1 g0149(.A(new_n346), .B1(new_n347), .B2(new_n345), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AOI211_X1 g0150(.A(new_n337), .B(new_n341), .C1(new_n350), .C2(new_n289), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G190), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n211), .A2(G1), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n325), .A2(G50), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n278), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n211), .B1(new_n201), .B2(new_n235), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT8), .B(G58), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G20), .A2(G33), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n358), .A2(new_n262), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n356), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n355), .B(new_n363), .C1(G50), .C2(new_n277), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT9), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n352), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n351), .A2(new_n368), .B1(new_n364), .B2(new_n365), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g0170(.A(new_n370), .B(KEYINPUT10), .Z(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n351), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n364), .C1(G169), .C2(new_n351), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n348), .A2(new_n303), .B1(new_n376), .B2(new_n345), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n342), .A2(new_n344), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n378), .A2(new_n224), .A3(G1698), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n289), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n337), .B1(G244), .B2(new_n340), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n276), .A2(new_n211), .A3(G33), .ZN(new_n385));
  INV_X1    g0185(.A(new_n358), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(new_n360), .B1(G20), .B2(G77), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n322), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n273), .A2(new_n267), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(G77), .A3(new_n354), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G77), .B2(new_n277), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n384), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n382), .A2(G179), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n382), .A2(G200), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n388), .A2(new_n391), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(new_n382), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT69), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n342), .A2(new_n344), .A3(G232), .A4(G1698), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n342), .A2(new_n344), .A3(G226), .A4(new_n304), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n289), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT70), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT70), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n409), .A3(new_n289), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n288), .A2(G238), .A3(new_n338), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n336), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT71), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT71), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n336), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n402), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n406), .A2(new_n409), .A3(new_n289), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n409), .B1(new_n406), .B2(new_n289), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n417), .B(new_n402), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(G169), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT14), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT72), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT72), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n428), .A3(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n427), .A2(G179), .A3(new_n429), .A4(new_n421), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n421), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(G169), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n424), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n360), .A2(G50), .B1(G20), .B2(new_n237), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n347), .B2(new_n262), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n356), .A2(KEYINPUT11), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n273), .A2(new_n237), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT12), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n389), .A2(G68), .A3(new_n354), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT11), .B1(new_n356), .B2(new_n436), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n431), .B2(G200), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n427), .A2(G190), .A3(new_n429), .A4(new_n421), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR4_X1   g0249(.A1(new_n375), .A2(new_n401), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n358), .A2(new_n353), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n325), .A2(new_n451), .B1(new_n273), .B2(new_n358), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G58), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n237), .ZN(new_n455));
  OAI21_X1  g0255(.A(G20), .B1(new_n455), .B2(new_n201), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n360), .A2(G159), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT7), .B1(new_n378), .B2(new_n211), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT7), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  AOI21_X1  g0262(.A(G33), .B1(new_n243), .B2(new_n244), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT3), .B1(new_n248), .B2(new_n249), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT76), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n247), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT73), .A2(G33), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT73), .A2(G33), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n343), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT76), .A3(new_n462), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n460), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n459), .B1(new_n476), .B2(new_n237), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT16), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n322), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n245), .A2(new_n250), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(new_n461), .A3(new_n211), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G68), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(new_n245), .B2(new_n250), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n461), .ZN(new_n484));
  OAI211_X1 g0284(.A(KEYINPUT16), .B(new_n459), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT75), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n237), .B1(new_n483), .B2(new_n461), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n471), .A2(new_n472), .A3(new_n343), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n468), .A2(new_n469), .A3(new_n247), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n211), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n458), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT75), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT16), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n453), .B1(new_n479), .B2(new_n495), .ZN(new_n496));
  MUX2_X1   g0296(.A(G223), .B(G226), .S(G1698), .Z(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(new_n245), .A3(new_n250), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G87), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n288), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n336), .B1(new_n224), .B2(new_n339), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n372), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n383), .B1(new_n500), .B2(new_n501), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT77), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n505), .B(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT18), .B1(new_n496), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n485), .A2(KEYINPUT75), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n493), .B1(new_n492), .B2(KEYINPUT16), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n460), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT76), .B1(new_n474), .B2(new_n462), .ZN(new_n513));
  INV_X1    g0313(.A(new_n462), .ZN(new_n514));
  AOI211_X1 g0314(.A(new_n466), .B(new_n514), .C1(new_n470), .C2(new_n473), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n458), .B1(new_n516), .B2(G68), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n267), .B1(new_n517), .B2(KEYINPUT16), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n452), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT18), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n505), .B(KEYINPUT77), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n508), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n502), .A2(G190), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n368), .B2(new_n502), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n452), .B(new_n526), .C1(new_n511), .C2(new_n518), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n496), .A2(KEYINPUT17), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n450), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n277), .A2(G97), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n326), .B2(new_n263), .ZN(new_n537));
  XNOR2_X1  g0337(.A(G97), .B(G107), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n539), .A2(new_n263), .A3(G107), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(G20), .B1(G77), .B2(new_n360), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n476), .B2(new_n376), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n537), .B1(new_n544), .B2(new_n267), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n245), .A2(new_n250), .A3(G244), .A4(new_n304), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n306), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n549), .A2(new_n304), .A3(new_n342), .A4(new_n344), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n342), .A2(new_n344), .A3(G250), .A4(G1698), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n289), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT5), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT5), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n334), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n271), .B(G45), .C1(new_n334), .C2(KEYINPUT5), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT78), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(G41), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT78), .B1(new_n300), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n562), .B(new_n297), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(G41), .B1(new_n558), .B2(new_n560), .ZN(new_n569));
  OAI211_X1 g0369(.A(G257), .B(new_n288), .C1(new_n569), .C2(new_n563), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT80), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(KEYINPUT80), .A3(new_n570), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n556), .A2(new_n573), .A3(new_n372), .A4(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n288), .B1(new_n548), .B2(new_n554), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n383), .B1(new_n576), .B2(new_n571), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n545), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n556), .A2(new_n574), .A3(new_n573), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(G200), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n580), .A3(G200), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n537), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n540), .A2(new_n541), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n587), .A2(new_n211), .B1(new_n347), .B2(new_n361), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n516), .B2(G107), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n589), .B2(new_n322), .ZN(new_n590));
  INV_X1    g0390(.A(new_n571), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n553), .B1(new_n547), .B2(new_n546), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(G190), .C1(new_n288), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n576), .A2(new_n571), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(KEYINPUT82), .A3(G190), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n590), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n579), .B1(new_n585), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n211), .A2(G116), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n272), .ZN(new_n602));
  INV_X1    g0402(.A(G116), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n279), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n389), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n322), .A2(new_n600), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n551), .B(new_n211), .C1(G33), .C2(new_n263), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT20), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(KEYINPUT20), .A2(new_n607), .A3(new_n601), .A4(new_n267), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G257), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n304), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n304), .A2(G264), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n245), .A2(new_n250), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n378), .A2(G303), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n288), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(G270), .B(new_n288), .C1(new_n569), .C2(new_n563), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n568), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n610), .B(G169), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n610), .ZN(new_n622));
  OAI21_X1  g0422(.A(G200), .B1(new_n618), .B2(new_n616), .ZN(new_n623));
  INV_X1    g0423(.A(new_n618), .ZN(new_n624));
  INV_X1    g0424(.A(new_n616), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n622), .B(new_n623), .C1(new_n626), .C2(new_n398), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(KEYINPUT21), .A3(G169), .A4(new_n610), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n618), .A2(new_n616), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(G179), .A3(new_n610), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n621), .A2(new_n627), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n309), .A2(G294), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n611), .A2(G1698), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G250), .B2(G1698), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n480), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n289), .ZN(new_n637));
  INV_X1    g0437(.A(new_n563), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n289), .B1(new_n562), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n569), .A2(new_n293), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n563), .A2(new_n564), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n300), .A2(KEYINPUT78), .A3(new_n566), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n639), .A2(G264), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n636), .B1(new_n635), .B2(new_n289), .ZN(new_n646));
  OAI21_X1  g0446(.A(G169), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n635), .A2(new_n289), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT89), .B1(new_n649), .B2(new_n372), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n644), .A2(new_n648), .A3(new_n651), .A4(G179), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n647), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n273), .A2(new_n376), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT25), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n326), .B2(new_n376), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT22), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n211), .A2(G87), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n378), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n376), .A2(G20), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT23), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n309), .A2(new_n211), .A3(G116), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n659), .A2(new_n256), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n245), .A2(new_n250), .A3(new_n211), .A4(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n671));
  INV_X1    g0471(.A(new_n669), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT87), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n670), .A2(KEYINPUT24), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n267), .B1(new_n673), .B2(KEYINPUT24), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n658), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n653), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n675), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n670), .A2(KEYINPUT24), .A3(new_n673), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n657), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n649), .A2(new_n368), .ZN(new_n681));
  INV_X1    g0481(.A(new_n646), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n637), .A3(new_n644), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n683), .B2(G190), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n631), .A2(new_n677), .A3(new_n685), .ZN(new_n686));
  AND4_X1   g0486(.A1(new_n333), .A2(new_n534), .A3(new_n599), .A4(new_n686), .ZN(G372));
  NAND2_X1  g0487(.A1(new_n318), .A2(new_n282), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n545), .B2(new_n578), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n590), .A2(KEYINPUT91), .A3(new_n575), .A4(new_n577), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n330), .A2(new_n688), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT26), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n690), .A2(new_n691), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n621), .A2(new_n628), .A3(new_n630), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n677), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n653), .A2(new_n676), .A3(KEYINPUT90), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n595), .A2(new_n597), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n581), .A2(new_n580), .A3(G200), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n700), .B(new_n545), .C1(new_n701), .C2(new_n582), .ZN(new_n702));
  INV_X1    g0502(.A(new_n579), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n703), .A3(new_n685), .A4(new_n692), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n688), .B(new_n694), .C1(new_n699), .C2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n693), .B1(new_n333), .B2(new_n579), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n534), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT92), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n523), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n508), .A2(new_n522), .A3(KEYINPUT92), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n448), .A2(new_n394), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n531), .B1(new_n444), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n371), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n715), .A2(new_n374), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(new_n716), .ZN(G369));
  OR3_X1    g0517(.A1(new_n272), .A2(KEYINPUT27), .A3(G20), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT27), .B1(new_n272), .B2(G20), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G213), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G343), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n610), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT93), .Z(new_n724));
  MUX2_X1   g0524(.A(new_n695), .B(new_n631), .S(new_n724), .Z(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n685), .A2(new_n677), .ZN(new_n728));
  INV_X1    g0528(.A(new_n722), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n680), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n677), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n697), .A2(new_n698), .A3(new_n729), .ZN(new_n733));
  INV_X1    g0533(.A(new_n695), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n722), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n732), .A2(new_n733), .A3(new_n736), .ZN(G399));
  INV_X1    g0537(.A(new_n207), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G41), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n257), .A2(G116), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n739), .A2(new_n271), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n210), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n742), .B1(new_n743), .B2(new_n739), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT28), .Z(new_n745));
  INV_X1    g0545(.A(G330), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n686), .A2(new_n599), .A3(new_n333), .A4(new_n729), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n626), .A2(new_n372), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n635), .A2(new_n289), .B1(new_n639), .B2(G264), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n320), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n748), .A2(new_n750), .A3(KEYINPUT30), .A4(new_n596), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT30), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n320), .A2(new_n629), .A3(G179), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n556), .A2(new_n591), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n320), .A2(G179), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n581), .A2(new_n756), .A3(new_n626), .A4(new_n649), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n722), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT31), .B1(new_n758), .B2(new_n722), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n746), .B1(new_n747), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT94), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n707), .A2(new_n729), .ZN(new_n765));
  XOR2_X1   g0565(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT26), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n319), .A2(new_n330), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT86), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n319), .A2(KEYINPUT86), .A3(new_n330), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n772), .A2(new_n693), .A3(new_n773), .A4(new_n579), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n769), .A2(new_n688), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT96), .ZN(new_n776));
  INV_X1    g0576(.A(new_n704), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n677), .A2(new_n734), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n769), .A2(new_n774), .A3(KEYINPUT96), .A4(new_n688), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n722), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT29), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n764), .B1(new_n767), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n745), .B1(new_n783), .B2(G1), .ZN(G364));
  INV_X1    g0584(.A(new_n739), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n211), .A2(G13), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n271), .B1(new_n786), .B2(G45), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT97), .Z(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n212), .B1(G20), .B2(new_n383), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n211), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(new_n398), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n376), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n211), .A2(new_n372), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n398), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n211), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n799), .A2(new_n454), .B1(new_n263), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n797), .A2(new_n368), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n795), .B(new_n802), .C1(G50), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G190), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n793), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n808));
  NAND3_X1  g0608(.A1(new_n807), .A2(G159), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(new_n807), .B2(G159), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(G87), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n796), .A2(new_n398), .A3(G200), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n345), .B1(new_n814), .B2(new_n237), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n796), .A2(new_n805), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(G77), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n804), .A2(new_n809), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n801), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G294), .B1(new_n812), .B2(G303), .ZN(new_n821));
  INV_X1    g0621(.A(new_n814), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n822), .A2(new_n823), .B1(new_n817), .B2(G311), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n345), .B1(new_n807), .B2(G329), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G322), .A2(new_n798), .B1(new_n803), .B2(G326), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n794), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n792), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(G13), .A2(G33), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT98), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(G20), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n791), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n207), .A2(G355), .A3(new_n345), .ZN(new_n835));
  INV_X1    g0635(.A(new_n480), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n738), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(G45), .B2(new_n210), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n241), .A2(new_n299), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n835), .B1(G116), .B2(new_n207), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n790), .B(new_n830), .C1(new_n834), .C2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  INV_X1    g0642(.A(new_n833), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n725), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n727), .A2(new_n789), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(G330), .B2(new_n725), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  OR2_X1    g0648(.A1(new_n791), .A2(new_n831), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n789), .B1(G77), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT101), .ZN(new_n851));
  INV_X1    g0651(.A(G311), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n816), .A2(new_n603), .B1(new_n806), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n345), .B(new_n853), .C1(G283), .C2(new_n822), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n798), .A2(G294), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n794), .A2(new_n256), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G303), .B2(new_n803), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n820), .A2(G97), .B1(new_n812), .B2(G107), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n854), .A2(new_n855), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n794), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(G68), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n235), .B2(new_n811), .C1(new_n454), .C2(new_n801), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n480), .B(new_n862), .C1(G132), .C2(new_n807), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n822), .A2(G150), .B1(new_n817), .B2(G159), .ZN(new_n865));
  INV_X1    g0665(.A(new_n803), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  INV_X1    g0667(.A(G143), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n865), .B1(new_n866), .B2(new_n867), .C1(new_n868), .C2(new_n799), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT34), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n859), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n791), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n399), .B1(new_n397), .B2(new_n729), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n395), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n394), .A2(new_n729), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n851), .B(new_n874), .C1(new_n878), .C2(new_n832), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n878), .B(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n765), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n729), .B(new_n878), .C1(new_n705), .C2(new_n706), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n764), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n885), .A2(new_n886), .A3(new_n789), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(new_n764), .A3(new_n883), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT104), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n880), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(G384));
  NAND2_X1  g0691(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n212), .A2(new_n211), .A3(new_n603), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n542), .B2(KEYINPUT35), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT106), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  XOR2_X1   g0697(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OR3_X1    g0699(.A1(new_n210), .A2(new_n347), .A3(new_n455), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n271), .B(G13), .C1(new_n900), .C2(new_n236), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n356), .B1(new_n492), .B2(KEYINPUT16), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n494), .B2(new_n486), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n521), .B1(new_n904), .B2(new_n453), .ZN(new_n905));
  INV_X1    g0705(.A(new_n720), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n904), .B2(new_n453), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n527), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n519), .A2(new_n521), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n720), .B(KEYINPUT108), .Z(new_n911));
  NAND2_X1  g0711(.A1(new_n519), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .A4(new_n527), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n907), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n523), .B2(new_n531), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n915), .A2(new_n917), .A3(KEYINPUT38), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n918), .ZN(new_n922));
  INV_X1    g0722(.A(new_n911), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n527), .B(KEYINPUT92), .C1(new_n496), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n910), .A2(new_n912), .A3(new_n527), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n496), .A2(new_n923), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n453), .B(new_n525), .C1(new_n479), .C2(new_n495), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n930), .A2(new_n709), .A3(KEYINPUT37), .A4(new_n910), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n531), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n710), .A2(new_n933), .A3(new_n711), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n922), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n921), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n444), .A2(new_n722), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n883), .A2(new_n877), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n443), .A2(new_n722), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n444), .A2(new_n448), .A3(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n443), .B(new_n722), .C1(new_n449), .C2(new_n434), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n919), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n922), .A2(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n947), .A2(new_n949), .B1(new_n712), .B2(new_n923), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n534), .A2(new_n782), .A3(new_n767), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n716), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n747), .A2(new_n761), .ZN(new_n955));
  AND4_X1   g0755(.A1(KEYINPUT40), .A2(new_n955), .A3(new_n945), .A4(new_n878), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n934), .A2(new_n928), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n930), .A2(new_n910), .B1(new_n924), .B2(KEYINPUT37), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n527), .B1(new_n496), .B2(new_n923), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n496), .A2(new_n507), .ZN(new_n960));
  NOR4_X1   g0760(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT92), .A4(new_n913), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n956), .B1(new_n963), .B2(new_n918), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n955), .A2(new_n945), .A3(new_n878), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n918), .B2(new_n919), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n533), .B1(new_n747), .B2(new_n761), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n746), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n970), .B2(new_n969), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n954), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT110), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n271), .B2(new_n786), .C1(new_n954), .C2(new_n972), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(KEYINPUT110), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n902), .B1(new_n975), .B2(new_n976), .ZN(G367));
  OAI211_X1 g0777(.A(new_n702), .B(new_n703), .C1(new_n545), .C2(new_n729), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n579), .A2(new_n722), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(new_n736), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT42), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n978), .A2(new_n677), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n722), .B1(new_n983), .B2(new_n703), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(KEYINPUT42), .B2(new_n981), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n328), .A2(new_n285), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n692), .B1(new_n986), .B2(new_n729), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n986), .A2(new_n688), .A3(new_n729), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n982), .A2(new_n985), .B1(KEYINPUT43), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n990), .B(new_n991), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n732), .A2(new_n980), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n739), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n736), .B1(new_n731), .B2(new_n735), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n727), .A2(KEYINPUT113), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n726), .B(KEYINPUT113), .Z(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n783), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n736), .A2(new_n733), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n980), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT44), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n980), .A2(new_n1004), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n732), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n732), .B1(new_n1009), .B2(KEYINPUT111), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1006), .A2(new_n1013), .A3(new_n1008), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT112), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1012), .A2(KEYINPUT112), .A3(new_n1014), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1003), .B(new_n1011), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n783), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n997), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n995), .B1(new_n1021), .B2(new_n787), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n837), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n834), .B1(new_n207), .B2(new_n270), .C1(new_n1023), .C2(new_n230), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n789), .A2(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n868), .A2(new_n866), .B1(new_n799), .B2(new_n359), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G58), .B2(new_n812), .ZN(new_n1027));
  INV_X1    g0827(.A(G159), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n814), .A2(new_n1028), .B1(new_n816), .B2(new_n235), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n378), .B(new_n1029), .C1(G137), .C2(new_n807), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n801), .A2(new_n237), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n794), .A2(new_n347), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1027), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(G294), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n814), .A2(new_n1035), .B1(new_n816), .B2(new_n828), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G317), .B2(new_n807), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n836), .B1(G97), .B2(new_n860), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n820), .A2(G107), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G303), .A2(new_n798), .B1(new_n803), .B2(G311), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n811), .A2(new_n603), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT46), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1034), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1025), .B1(new_n1045), .B2(new_n791), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n987), .A2(new_n833), .A3(new_n988), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1022), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G387));
  INV_X1    g0851(.A(new_n787), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1002), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n207), .A2(new_n345), .A3(new_n741), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(G107), .B2(new_n207), .ZN(new_n1055));
  AOI211_X1 g0855(.A(G45), .B(new_n741), .C1(G68), .C2(G77), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1058));
  OR3_X1    g0858(.A1(new_n358), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT50), .B1(new_n358), .B2(G50), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1023), .B1(new_n227), .B2(G45), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n834), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n789), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n799), .A2(new_n235), .B1(new_n811), .B2(new_n347), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G159), .B2(new_n803), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n276), .A2(new_n820), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n822), .A2(new_n386), .B1(new_n807), .B2(G150), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n237), .B2(new_n816), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n480), .B1(G97), .B2(new_n860), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n836), .B1(G326), .B2(new_n807), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n801), .A2(new_n828), .B1(new_n811), .B2(new_n1035), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n822), .A2(G311), .B1(new_n817), .B2(G303), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n798), .A2(G317), .ZN(new_n1077));
  INV_X1    g0877(.A(G322), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1076), .B(new_n1077), .C1(new_n1078), .C2(new_n866), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT48), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1075), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1080), .B2(new_n1079), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT49), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1074), .B1(new_n603), .B2(new_n794), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1073), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1065), .B1(new_n1086), .B2(new_n791), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n731), .B2(new_n843), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1003), .ZN(new_n1089));
  OAI21_X1  g0889(.A(KEYINPUT115), .B1(new_n1089), .B2(new_n785), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n783), .B2(new_n1002), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(KEYINPUT115), .A3(new_n785), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1053), .B(new_n1088), .C1(new_n1091), .C2(new_n1092), .ZN(G393));
  AOI21_X1  g0893(.A(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1089), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1009), .B(new_n1010), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n739), .C1(new_n1089), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n980), .A2(new_n833), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n834), .B1(new_n263), .B2(new_n207), .C1(new_n1023), .C2(new_n234), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n789), .A2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT116), .Z(new_n1102));
  NOR2_X1   g0902(.A1(new_n801), .A2(new_n347), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n856), .B(new_n1103), .C1(G68), .C2(new_n812), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n814), .A2(new_n235), .B1(new_n816), .B2(new_n358), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n480), .B1(G143), .B2(new_n807), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G150), .A2(new_n803), .B1(new_n798), .B2(G159), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT51), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G311), .A2(new_n798), .B1(new_n803), .B2(G317), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT52), .Z(new_n1116));
  OAI22_X1  g0916(.A1(new_n816), .A2(new_n1035), .B1(new_n806), .B2(new_n1078), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n345), .B(new_n1117), .C1(G303), .C2(new_n822), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n811), .A2(new_n828), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n795), .B(new_n1119), .C1(G116), .C2(new_n820), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1113), .A2(new_n1114), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1102), .B1(new_n791), .B2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1097), .A2(new_n1052), .B1(new_n1099), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1098), .A2(new_n1124), .ZN(G390));
  INV_X1    g0925(.A(KEYINPUT120), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n945), .B1(new_n764), .B2(new_n878), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n762), .A2(new_n878), .A3(new_n945), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n940), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n955), .A2(G330), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n763), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n762), .A2(KEYINPUT94), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n878), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1128), .B1(new_n1133), .B2(new_n946), .ZN(new_n1134));
  OAI21_X1  g0934(.A(KEYINPUT120), .B1(new_n1134), .B2(new_n941), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n764), .A2(new_n878), .A3(new_n945), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n877), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n781), .B2(new_n876), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n946), .B1(new_n881), .B2(new_n1130), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n952), .B(new_n716), .C1(new_n533), .C2(new_n1130), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n938), .B1(new_n940), .B2(new_n945), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n920), .B1(new_n963), .B2(new_n918), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n948), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n938), .B(KEYINPUT119), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n963), .B2(new_n918), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n775), .A2(new_n776), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n777), .A2(new_n778), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n780), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n729), .A3(new_n876), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n946), .B1(new_n1156), .B2(new_n877), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1128), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n936), .B(new_n1151), .C1(new_n1139), .C2(new_n946), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n1137), .C1(new_n937), .C2(new_n1147), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1146), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1143), .A2(new_n1145), .A3(new_n1161), .A4(new_n1159), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n739), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n789), .B1(new_n386), .B2(new_n849), .ZN(new_n1166));
  INV_X1    g0966(.A(G132), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n799), .A2(new_n1167), .B1(new_n1028), .B2(new_n801), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n866), .A2(new_n1169), .B1(new_n794), .B2(new_n235), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n811), .A2(new_n359), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT53), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n378), .B1(new_n817), .B2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n822), .A2(G137), .B1(new_n807), .B2(G125), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1171), .A2(new_n1173), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n816), .A2(new_n263), .B1(new_n806), .B2(new_n1035), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n345), .B(new_n1179), .C1(G107), .C2(new_n822), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n861), .C1(new_n256), .C2(new_n811), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1103), .B1(G116), .B2(new_n798), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n828), .B2(new_n866), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1178), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1166), .B1(new_n791), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n937), .B2(new_n832), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n1162), .B2(new_n787), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1165), .B1(new_n1189), .B2(new_n1190), .ZN(G378));
  NAND3_X1  g0991(.A1(new_n964), .A2(new_n968), .A3(G330), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n364), .A2(new_n906), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n375), .B(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n375), .B1(new_n364), .B2(new_n906), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1193), .B1(new_n371), .B2(new_n374), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1192), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n964), .A3(new_n968), .A4(G330), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n951), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n939), .A3(new_n1204), .A4(new_n950), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1201), .A2(new_n832), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n789), .B1(G50), .B2(new_n849), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n480), .B2(new_n334), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G41), .B(new_n836), .C1(G77), .C2(new_n812), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT122), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n860), .A2(G58), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n866), .B2(new_n603), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G107), .B2(new_n798), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n814), .A2(new_n263), .B1(new_n806), .B2(new_n828), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1031), .B(new_n1220), .C1(new_n276), .C2(new_n817), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1215), .A2(new_n1216), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1212), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n798), .A2(G128), .B1(new_n812), .B2(new_n1175), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT123), .Z(new_n1226));
  AOI22_X1  g1026(.A1(G150), .A2(new_n820), .B1(new_n803), .B2(G125), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT124), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n822), .A2(G132), .B1(new_n817), .B2(G137), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n860), .A2(G159), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G33), .B(G41), .C1(new_n807), .C2(G124), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1224), .B1(new_n1223), .B2(new_n1222), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1210), .B1(new_n1236), .B2(new_n791), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1208), .A2(new_n1052), .B1(new_n1209), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1141), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1145), .B1(new_n1162), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n1208), .A3(KEYINPUT57), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1208), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n739), .B(new_n1241), .C1(new_n1242), .C2(KEYINPUT125), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1244), .B(KEYINPUT57), .C1(new_n1240), .C2(new_n1208), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1238), .B1(new_n1243), .B2(new_n1245), .ZN(G375));
  NAND2_X1  g1046(.A1(new_n1239), .A2(new_n1144), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1146), .A2(new_n997), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n946), .A2(new_n831), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n789), .B1(G68), .B2(new_n849), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1217), .B1(new_n866), .B2(new_n1167), .C1(new_n867), .C2(new_n799), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n480), .B(new_n1251), .C1(new_n822), .C2(new_n1175), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n801), .A2(new_n235), .B1(new_n816), .B2(new_n359), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT126), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n811), .A2(new_n1028), .B1(new_n806), .B2(new_n1169), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT127), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n814), .A2(new_n603), .B1(new_n816), .B2(new_n376), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n345), .B(new_n1258), .C1(G303), .C2(new_n807), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1032), .B1(G283), .B2(new_n798), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n803), .A2(G294), .B1(new_n812), .B2(G97), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1259), .A2(new_n1068), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1250), .B1(new_n1263), .B2(new_n791), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1249), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1239), .B2(new_n787), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1248), .A2(new_n1267), .ZN(G381));
  INV_X1    g1068(.A(G390), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1050), .A2(new_n890), .A3(new_n1269), .ZN(new_n1270));
  OR3_X1    g1070(.A1(G381), .A2(G393), .A3(G396), .ZN(new_n1271));
  OR4_X1    g1071(.A1(G378), .A2(new_n1270), .A3(G375), .A4(new_n1271), .ZN(G407));
  INV_X1    g1072(.A(G378), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n721), .A2(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(G375), .C2(new_n1276), .ZN(G409));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1238), .C1(new_n1243), .C2(new_n1245), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1240), .A2(new_n1208), .A3(new_n997), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1238), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1281), .B(new_n1165), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1274), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1239), .A2(KEYINPUT60), .A3(new_n1144), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1285), .A2(new_n739), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1239), .A2(new_n1144), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1247), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1290), .B2(new_n1267), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n890), .B(new_n1266), .C1(new_n1286), .C2(new_n1289), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1278), .B1(new_n1284), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1267), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n890), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1290), .A2(G384), .A3(new_n1267), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1275), .A2(G2897), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1299), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1269), .B1(new_n1022), .B2(new_n1049), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(G393), .B(new_n847), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n996), .B1(new_n1095), .B2(new_n783), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n994), .B1(new_n1307), .B2(new_n1052), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1048), .A3(G390), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1305), .A2(new_n1306), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1306), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1275), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1293), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1295), .A2(new_n1304), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1313), .A2(new_n1316), .A3(new_n1293), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1318), .B1(new_n1313), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1316), .B1(new_n1313), .B2(new_n1293), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1317), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1322), .B2(new_n1312), .ZN(G405));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1273), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1324), .A2(new_n1294), .A3(new_n1279), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1294), .B1(new_n1324), .B2(new_n1279), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(new_n1312), .ZN(G402));
endmodule


