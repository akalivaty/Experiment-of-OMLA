//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G238), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT65), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n218), .B(new_n223), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AND2_X1   g0031(.A1(new_n229), .A2(new_n230), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n208), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n211), .B(new_n216), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT68), .B(G50), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n256), .A2(new_n206), .A3(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n214), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n205), .A2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G50), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n257), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(G50), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT71), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT8), .B(G58), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n206), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G150), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n206), .B1(new_n201), .B2(new_n220), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n259), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT70), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT70), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G222), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n282), .B2(new_n287), .ZN(new_n293));
  AOI22_X1  g0093(.A1(G77), .A2(new_n289), .B1(new_n293), .B2(G223), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n278), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n277), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n278), .A2(new_n296), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n221), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G190), .ZN(new_n305));
  OAI21_X1  g0105(.A(G200), .B1(new_n295), .B2(new_n303), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n276), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT10), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n275), .B1(new_n304), .B2(G169), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n295), .A2(G179), .A3(new_n303), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G68), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT12), .B1(new_n257), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n217), .A2(new_n206), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n256), .A2(G1), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n318), .A2(KEYINPUT12), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n260), .A2(G68), .A3(new_n261), .ZN(new_n321));
  INV_X1    g0121(.A(G77), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n271), .A2(new_n220), .B1(new_n268), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n259), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT11), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n320), .B(new_n321), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n325), .B2(new_n324), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT74), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT75), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n293), .A2(G232), .B1(G33), .B2(G97), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n288), .A2(G226), .A3(new_n292), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n278), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G238), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n301), .B1(new_n335), .B2(new_n302), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT13), .B1(new_n334), .B2(new_n336), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n331), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n339), .A2(KEYINPUT75), .A3(G179), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n339), .B2(new_n340), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n330), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n341), .A2(G200), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n339), .A2(G190), .A3(new_n340), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n329), .A3(new_n355), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n267), .A2(new_n271), .B1(new_n206), .B2(new_n322), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n268), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n259), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n360), .B(KEYINPUT72), .Z(new_n361));
  AOI21_X1  g0161(.A(new_n322), .B1(new_n205), .B2(G20), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n260), .A2(new_n362), .B1(new_n322), .B2(new_n257), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n290), .A2(G232), .ZN(new_n365));
  AOI22_X1  g0165(.A1(G107), .A2(new_n289), .B1(new_n293), .B2(G238), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n277), .ZN(new_n368));
  INV_X1    g0168(.A(new_n302), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(G244), .B1(new_n298), .B2(new_n300), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n364), .B1(new_n372), .B2(G169), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(G179), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g0175(.A(new_n364), .B(KEYINPUT73), .Z(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(G190), .B2(new_n372), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n371), .A2(G200), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n314), .A2(new_n353), .A3(new_n356), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT79), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n267), .B1(new_n205), .B2(G20), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n260), .B1(new_n257), .B2(new_n267), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n385));
  NOR2_X1   g0185(.A1(KEYINPUT7), .A2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n282), .A2(new_n287), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n286), .A2(new_n206), .ZN(new_n388));
  AND2_X1   g0188(.A1(KEYINPUT76), .A2(G33), .ZN(new_n389));
  NOR2_X1   g0189(.A1(KEYINPUT76), .A2(G33), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(new_n283), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n387), .B(new_n217), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(KEYINPUT64), .A2(G68), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT64), .A2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(G58), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n202), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(G20), .B1(G159), .B2(new_n270), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n385), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT78), .ZN(new_n401));
  INV_X1    g0201(.A(new_n259), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n201), .B1(new_n217), .B2(G58), .ZN(new_n403));
  INV_X1    g0203(.A(G159), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n403), .A2(new_n206), .B1(new_n404), .B2(new_n271), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT3), .B1(new_n389), .B2(new_n390), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n406), .A2(new_n393), .A3(new_n206), .A4(new_n285), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n285), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(G20), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n405), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n402), .B1(new_n411), .B2(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n384), .B1(new_n401), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n369), .A2(G232), .B1(new_n298), .B2(new_n300), .ZN(new_n414));
  NOR2_X1   g0214(.A1(G223), .A2(G1698), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n221), .B2(G1698), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n409), .A2(new_n416), .B1(G33), .B2(G87), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n278), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G200), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G190), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n414), .B(new_n421), .C1(new_n278), .C2(new_n417), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n381), .B1(new_n413), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n394), .A2(new_n399), .ZN(new_n425));
  INV_X1    g0225(.A(new_n385), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT78), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n400), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n412), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n431), .A2(new_n423), .A3(new_n381), .A4(new_n383), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT17), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n418), .A2(new_n342), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(G169), .B2(new_n418), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n413), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n383), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n418), .A2(G169), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n342), .B2(new_n418), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n431), .A2(new_n383), .A3(new_n423), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT17), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n434), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n380), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n228), .A2(G1698), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(G250), .B2(G1698), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n285), .B2(new_n406), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT76), .B(G33), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G294), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT85), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT85), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n281), .B1(new_n452), .B2(KEYINPUT3), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n453), .C1(new_n457), .C2(new_n450), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n277), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n277), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G264), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT86), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n300), .A2(new_n461), .A3(new_n462), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n459), .A2(KEYINPUT86), .A3(new_n464), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n467), .A2(G179), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(new_n468), .A3(new_n464), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G169), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n409), .A2(new_n206), .A3(G87), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n225), .A2(KEYINPUT22), .A3(G20), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n474), .A2(KEYINPUT22), .B1(new_n288), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n452), .A2(new_n206), .A3(G116), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n206), .A2(G107), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT23), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT24), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n476), .A2(KEYINPUT24), .A3(new_n480), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n259), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n260), .B1(G1), .B2(new_n284), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT25), .B1(new_n257), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n486), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n473), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n419), .ZN(new_n496));
  INV_X1    g0296(.A(new_n471), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n421), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n492), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(KEYINPUT87), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n495), .A2(new_n419), .B1(new_n421), .B2(new_n497), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n492), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n494), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n387), .B(G107), .C1(new_n392), .C2(new_n393), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n227), .A2(new_n486), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n486), .A2(KEYINPUT6), .A3(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n270), .A2(G77), .ZN(new_n514));
  XOR2_X1   g0314(.A(new_n514), .B(KEYINPUT80), .Z(new_n515));
  NAND3_X1  g0315(.A1(new_n506), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n516), .A2(new_n259), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n257), .A2(new_n227), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n485), .B2(new_n227), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n463), .A2(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n468), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n409), .A2(G244), .A3(new_n292), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n292), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n293), .A2(G250), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n523), .B1(new_n530), .B2(new_n277), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n531), .A2(G179), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n347), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n521), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(G190), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n520), .C1(new_n419), .C2(new_n531), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n462), .A2(new_n461), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(new_n278), .A3(G270), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n468), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n228), .A2(new_n292), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(G264), .B2(new_n292), .ZN(new_n543));
  INV_X1    g0343(.A(G303), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n457), .A2(new_n543), .B1(new_n288), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n541), .B1(new_n277), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n260), .B(G116), .C1(G1), .C2(new_n284), .ZN(new_n547));
  INV_X1    g0347(.A(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n257), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n528), .B(new_n206), .C1(G33), .C2(new_n227), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(new_n259), .C1(new_n206), .C2(G116), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT20), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n547), .B(new_n549), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n546), .A2(G179), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT83), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT83), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n546), .A2(new_n558), .A3(new_n555), .A4(G179), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n545), .A2(new_n277), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n468), .A3(new_n540), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(G169), .A3(new_n555), .ZN(new_n563));
  NOR2_X1   g0363(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n555), .B1(new_n562), .B2(G200), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n421), .B2(new_n562), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n560), .A2(new_n565), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n358), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n263), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n409), .A2(new_n206), .A3(G68), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n206), .B1(new_n284), .B2(new_n227), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n509), .A2(new_n225), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n268), .A2(KEYINPUT19), .A3(new_n227), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n571), .B1(new_n578), .B2(new_n259), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n358), .B2(new_n485), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n335), .A2(G1698), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n409), .A2(new_n581), .B1(G116), .B2(new_n452), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n409), .A2(G244), .A3(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n278), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n461), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n278), .A2(G250), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n300), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(new_n585), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n342), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n347), .B1(new_n584), .B2(new_n588), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n580), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n485), .A2(new_n225), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n579), .B(new_n595), .C1(new_n589), .C2(new_n419), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(KEYINPUT82), .B1(G190), .B2(new_n589), .ZN(new_n597));
  AOI211_X1 g0397(.A(new_n571), .B(new_n594), .C1(new_n259), .C2(new_n578), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT82), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n419), .C2(new_n589), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n593), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n538), .A2(new_n569), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n537), .B1(new_n534), .B2(new_n536), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n448), .A2(new_n505), .A3(new_n604), .ZN(G372));
  INV_X1    g0405(.A(new_n356), .ZN(new_n606));
  INV_X1    g0406(.A(new_n375), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n353), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n434), .A3(new_n446), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n413), .A2(new_n437), .A3(new_n435), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT18), .B1(new_n439), .B2(new_n441), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n438), .A2(KEYINPUT89), .A3(new_n442), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n311), .B1(new_n615), .B2(new_n308), .ZN(new_n616));
  INV_X1    g0416(.A(new_n448), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n589), .A2(G190), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n600), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n531), .A2(G179), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n347), .B2(new_n531), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n620), .A2(new_n521), .A3(new_n622), .A4(new_n592), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT26), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n520), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n598), .B(new_n619), .C1(new_n419), .C2(new_n589), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(new_n592), .ZN(new_n629));
  INV_X1    g0429(.A(new_n533), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(KEYINPUT88), .A3(new_n621), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n626), .A2(new_n627), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n624), .A2(new_n632), .A3(new_n592), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n565), .A2(new_n560), .A3(new_n566), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n493), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n629), .A2(new_n534), .A3(new_n536), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n504), .B2(new_n501), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n616), .B1(new_n617), .B2(new_n638), .ZN(G369));
  NAND2_X1  g0439(.A1(new_n318), .A2(new_n206), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(G213), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n493), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n492), .A2(new_n645), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT87), .B1(new_n499), .B2(new_n500), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n503), .A2(new_n492), .A3(new_n502), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n493), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n494), .A2(new_n645), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT90), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n650), .A2(new_n654), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n634), .A2(new_n645), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n646), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n555), .A2(new_n645), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n569), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n634), .B2(new_n659), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n658), .A2(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n209), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n509), .A2(new_n225), .A3(new_n548), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n668), .A2(G1), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n212), .B2(new_n668), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  INV_X1    g0474(.A(new_n645), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n604), .A2(new_n505), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT91), .B1(new_n562), .B2(new_n342), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n546), .A2(new_n678), .A3(G179), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n677), .A2(new_n589), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n467), .A2(new_n469), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n680), .A2(KEYINPUT30), .A3(new_n682), .A4(new_n531), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n677), .A2(new_n531), .A3(new_n589), .A4(new_n679), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n681), .ZN(new_n686));
  NOR4_X1   g0486(.A1(new_n531), .A2(G179), .A3(new_n589), .A4(new_n546), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n495), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n683), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n645), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT31), .B1(new_n689), .B2(new_n645), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n674), .B1(new_n676), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n592), .B1(new_n623), .B2(KEYINPUT26), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(KEYINPUT26), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n635), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n634), .A2(new_n493), .A3(KEYINPUT92), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n637), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n645), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n638), .B2(new_n645), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n693), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n673), .B1(new_n705), .B2(G1), .ZN(G364));
  NOR2_X1   g0506(.A1(new_n256), .A2(G20), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n205), .B1(new_n707), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n667), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n663), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G330), .B2(new_n661), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n288), .A2(new_n209), .ZN(new_n713));
  INV_X1    g0513(.A(G355), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(G116), .B2(new_n209), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n251), .A2(G45), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n457), .A2(new_n209), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n460), .B2(new_n213), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n715), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n214), .B1(G20), .B2(new_n347), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n710), .B1(new_n719), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n206), .A2(new_n421), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n342), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n206), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(G58), .A2(new_n730), .B1(new_n733), .B2(G77), .ZN(new_n734));
  NAND3_X1  g0534(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n421), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n220), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT93), .Z(new_n739));
  NOR2_X1   g0539(.A1(new_n419), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n727), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n731), .A2(new_n740), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n288), .B1(new_n225), .B2(new_n741), .C1(new_n486), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G159), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n735), .A2(G190), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n747), .A2(KEYINPUT32), .B1(new_n748), .B2(G68), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n206), .B1(new_n744), .B2(G190), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n749), .B1(KEYINPUT32), .B2(new_n747), .C1(new_n227), .C2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n739), .A2(new_n743), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT94), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT94), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT33), .B(G317), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n730), .A2(G322), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  INV_X1    g0557(.A(new_n741), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G303), .A2(new_n758), .B1(new_n733), .B2(G311), .ZN(new_n759));
  INV_X1    g0559(.A(new_n742), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G283), .A2(new_n760), .B1(new_n746), .B2(G329), .ZN(new_n761));
  INV_X1    g0561(.A(G294), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n289), .B1(new_n762), .B2(new_n750), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G326), .B2(new_n736), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n757), .A2(new_n759), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n753), .A2(new_n754), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n726), .B1(new_n766), .B2(new_n723), .ZN(new_n767));
  INV_X1    g0567(.A(new_n722), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n661), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n712), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(G396));
  NOR2_X1   g0571(.A1(new_n638), .A2(new_n645), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n364), .A2(new_n645), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n379), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n375), .A2(new_n645), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT97), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n772), .B(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n693), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT98), .Z(new_n782));
  AOI21_X1  g0582(.A(new_n710), .B1(new_n779), .B2(new_n780), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n723), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n721), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n710), .B1(G77), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT96), .ZN(new_n788));
  INV_X1    g0588(.A(new_n748), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(new_n750), .B2(new_n227), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G303), .B2(new_n736), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n741), .A2(new_n486), .B1(new_n732), .B2(new_n548), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G311), .B2(new_n746), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n742), .A2(new_n225), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G294), .B2(new_n730), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n792), .A2(new_n794), .A3(new_n289), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n742), .A2(new_n315), .B1(new_n745), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G50), .B2(new_n758), .ZN(new_n800));
  INV_X1    g0600(.A(new_n750), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n457), .B1(G58), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n730), .B1(new_n733), .B2(G159), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n737), .B2(new_n804), .C1(new_n269), .C2(new_n789), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n800), .B(new_n802), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n797), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n788), .B1(new_n809), .B2(new_n723), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n778), .B2(new_n721), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n784), .A2(new_n811), .ZN(G384));
  INV_X1    g0612(.A(KEYINPUT40), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n393), .B1(new_n457), .B2(new_n206), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n407), .A2(G68), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n399), .B(KEYINPUT16), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n259), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n410), .A2(G68), .A3(new_n407), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n385), .B1(new_n818), .B2(new_n399), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n383), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT100), .ZN(new_n821));
  INV_X1    g0621(.A(new_n643), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT100), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n823), .B(new_n383), .C1(new_n817), .C2(new_n819), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n447), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT38), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n424), .A2(new_n433), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT102), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n413), .B2(new_n643), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n439), .A2(KEYINPUT102), .A3(new_n822), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT37), .B1(new_n439), .B2(new_n441), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n828), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n444), .A2(KEYINPUT79), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n440), .B(new_n643), .C1(new_n342), .C2(new_n418), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n821), .A2(new_n836), .A3(new_n824), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n835), .A2(new_n432), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n838), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT101), .B1(new_n838), .B2(KEYINPUT37), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n834), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT103), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n834), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n827), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT101), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n838), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n843), .B1(new_n850), .B2(new_n834), .ZN(new_n851));
  INV_X1    g0651(.A(new_n844), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n826), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n845), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n676), .A2(new_n692), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n329), .A2(new_n675), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n353), .A2(new_n356), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n345), .A2(new_n356), .A3(new_n350), .A4(new_n351), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT99), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT99), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n863), .A3(new_n857), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n859), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n856), .A2(new_n865), .A3(new_n778), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n813), .B1(new_n855), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n813), .ZN(new_n868));
  INV_X1    g0668(.A(new_n827), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n851), .B2(new_n852), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n610), .B1(new_n413), .B2(new_n437), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n439), .A2(KEYINPUT89), .A3(new_n441), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n444), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT102), .B1(new_n439), .B2(new_n822), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n829), .B(new_n643), .C1(new_n431), .C2(new_n383), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n833), .A2(new_n835), .A3(new_n432), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT104), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT104), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n828), .A2(new_n832), .A3(new_n880), .A4(new_n833), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n613), .A2(new_n434), .A3(new_n446), .A4(new_n614), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n876), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n854), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n870), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n868), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n867), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n448), .A2(new_n856), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(G330), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT106), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n822), .B1(new_n613), .B2(new_n614), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n607), .A2(new_n645), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n772), .B2(new_n778), .ZN(new_n898));
  INV_X1    g0698(.A(new_n865), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n842), .A2(new_n844), .B1(new_n447), .B2(new_n825), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n870), .B1(new_n901), .B2(KEYINPUT38), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n896), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n886), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT105), .B1(new_n905), .B2(new_n845), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT39), .B1(new_n885), .B2(new_n854), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n870), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n906), .A2(new_n909), .B1(new_n902), .B2(KEYINPUT39), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n353), .A2(new_n645), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n903), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n448), .A2(new_n704), .A3(new_n702), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n616), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n913), .B(new_n915), .Z(new_n916));
  OAI22_X1  g0716(.A1(new_n895), .A2(new_n916), .B1(new_n205), .B2(new_n707), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n916), .B2(new_n895), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(G116), .A3(new_n215), .A4(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT36), .Z(new_n922));
  NAND3_X1  g0722(.A1(new_n213), .A2(G77), .A3(new_n397), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n220), .A2(G68), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n205), .B(G13), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  OR3_X1    g0725(.A1(new_n918), .A2(new_n922), .A3(new_n925), .ZN(G367));
  OAI221_X1 g0726(.A(new_n724), .B1(new_n209), .B2(new_n358), .C1(new_n245), .C2(new_n717), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(new_n710), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n741), .A2(new_n548), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n929), .A2(KEYINPUT46), .B1(new_n762), .B2(new_n789), .ZN(new_n930));
  XOR2_X1   g0730(.A(KEYINPUT111), .B(G311), .Z(new_n931));
  OAI22_X1  g0731(.A1(new_n737), .A2(new_n931), .B1(new_n486), .B2(new_n750), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(G283), .A2(new_n733), .B1(new_n746), .B2(G317), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n742), .A2(new_n227), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G303), .B2(new_n730), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n409), .B1(new_n929), .B2(KEYINPUT46), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n933), .A2(new_n934), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(G143), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n737), .A2(new_n939), .B1(new_n729), .B2(new_n269), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n750), .A2(new_n315), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n220), .A2(new_n732), .B1(new_n742), .B2(new_n322), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n741), .A2(new_n248), .B1(new_n745), .B2(new_n804), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n289), .B1(G159), .B2(new_n748), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n938), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n598), .A2(new_n675), .ZN(new_n952));
  MUX2_X1   g0752(.A(new_n629), .B(new_n593), .S(new_n952), .Z(new_n953));
  OAI221_X1 g0753(.A(new_n928), .B1(new_n785), .B2(new_n951), .C1(new_n953), .C2(new_n768), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n626), .A2(new_n631), .A3(new_n645), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n534), .B(new_n536), .C1(new_n520), .C2(new_n675), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n650), .A2(new_n654), .A3(new_n651), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n654), .B1(new_n650), .B2(new_n651), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n657), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n494), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n645), .B1(new_n962), .B2(new_n534), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n960), .B2(KEYINPUT42), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT107), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT42), .ZN(new_n967));
  INV_X1    g0767(.A(new_n657), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n653), .B2(new_n655), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n969), .B2(new_n957), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT107), .B1(new_n970), .B2(new_n963), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT108), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n966), .A2(new_n971), .A3(KEYINPUT108), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n966), .A2(new_n971), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n953), .B(KEYINPUT43), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n957), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n664), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(KEYINPUT109), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n977), .A2(new_n983), .A3(new_n980), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n667), .B(KEYINPUT41), .Z(new_n987));
  OAI21_X1  g0787(.A(new_n657), .B1(new_n958), .B2(new_n959), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n653), .A2(new_n655), .A3(new_n968), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n662), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n989), .A3(new_n663), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n705), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT110), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n658), .B2(new_n957), .ZN(new_n997));
  INV_X1    g0797(.A(new_n646), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n988), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(KEYINPUT44), .A3(new_n982), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n999), .B2(new_n982), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n658), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n664), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1001), .A2(new_n1005), .A3(new_n664), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n995), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n987), .B1(new_n1010), .B2(new_n705), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n985), .B(new_n986), .C1(new_n1011), .C2(new_n709), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT109), .B1(new_n981), .B2(new_n984), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n954), .B1(new_n1012), .B2(new_n1013), .ZN(G387));
  NOR2_X1   g0814(.A1(new_n241), .A2(new_n460), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1015), .A2(new_n717), .B1(new_n670), .B2(new_n713), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n267), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT50), .B1(new_n267), .B2(G50), .ZN(new_n1018));
  AOI21_X1  g0818(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1017), .A2(new_n670), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1020), .B1(new_n486), .B2(new_n666), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n710), .B1(new_n1021), .B2(new_n725), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n656), .A2(new_n768), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G116), .A2(new_n760), .B1(new_n746), .B2(G326), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n741), .A2(new_n762), .B1(new_n750), .B2(new_n790), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G317), .A2(new_n730), .B1(new_n733), .B2(G303), .ZN(new_n1026));
  INV_X1    g0826(.A(G322), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n737), .B2(new_n1027), .C1(new_n789), .C2(new_n931), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1025), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n457), .B(new_n1024), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n267), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1035), .A2(new_n748), .B1(G159), .B2(new_n736), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n801), .A2(new_n570), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n409), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n935), .B1(G68), .B2(new_n733), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n220), .B2(new_n729), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G77), .A2(new_n758), .B1(new_n746), .B2(G150), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1040), .B1(KEYINPUT113), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT113), .B2(new_n1041), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1033), .A2(new_n1034), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1022), .B(new_n1023), .C1(new_n723), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n991), .A2(new_n992), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1045), .B1(new_n1047), .B2(new_n709), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n667), .B(KEYINPUT114), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n1047), .B2(new_n705), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n995), .B2(new_n1050), .ZN(G393));
  AND3_X1   g0851(.A1(new_n1001), .A2(new_n1005), .A3(new_n664), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n664), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(new_n995), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n1010), .A3(new_n1049), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n982), .A2(new_n722), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n724), .B1(new_n227), .B2(new_n209), .C1(new_n254), .C2(new_n717), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n710), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n732), .A2(new_n267), .B1(new_n745), .B2(new_n939), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n795), .B(new_n1060), .C1(new_n217), .C2(new_n758), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n737), .A2(new_n269), .B1(new_n729), .B2(new_n404), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n750), .A2(new_n322), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1064), .B(new_n457), .C1(G50), .C2(new_n748), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n741), .A2(new_n790), .B1(new_n745), .B2(new_n1027), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT115), .Z(new_n1068));
  OAI221_X1 g0868(.A(new_n289), .B1(new_n486), .B2(new_n742), .C1(new_n762), .C2(new_n732), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n789), .A2(new_n544), .B1(new_n750), .B2(new_n548), .ZN(new_n1070));
  OR3_X1    g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n730), .A2(G311), .B1(G317), .B2(new_n736), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1066), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1059), .B1(new_n1074), .B2(new_n723), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1054), .A2(new_n709), .B1(new_n1057), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1056), .A2(new_n1076), .ZN(G390));
  INV_X1    g0877(.A(KEYINPUT116), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n693), .A2(new_n778), .A3(new_n865), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n865), .B1(new_n693), .B2(new_n778), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1081), .B2(new_n898), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n693), .A2(new_n778), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n899), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n693), .A2(new_n778), .A3(new_n865), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n898), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(KEYINPUT116), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n897), .B1(new_n701), .B2(new_n778), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1081), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1082), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n914), .B(new_n616), .C1(new_n617), .C2(new_n780), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n842), .A2(new_n844), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT38), .B1(new_n1094), .B2(new_n826), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT39), .B1(new_n1095), .B2(new_n845), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n912), .B1(new_n898), .B2(new_n899), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n908), .B1(new_n870), .B2(new_n907), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n870), .A2(new_n907), .A3(new_n908), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n887), .B(new_n912), .C1(new_n899), .C2(new_n1088), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1100), .A2(new_n1085), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1085), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1093), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1079), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1100), .A2(new_n1085), .A3(new_n1101), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1086), .A2(KEYINPUT116), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1091), .B1(new_n1108), .B2(new_n1082), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1104), .A2(new_n1110), .A3(new_n1049), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1064), .B1(new_n736), .B2(G283), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n486), .B2(new_n789), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G97), .A2(new_n733), .B1(new_n746), .B2(G294), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n548), .B2(new_n729), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n741), .A2(new_n225), .B1(new_n742), .B2(new_n315), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1113), .A2(new_n1115), .A3(new_n288), .A4(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n729), .A2(new_n798), .B1(new_n732), .B2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n801), .A2(G159), .B1(G137), .B2(new_n748), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT53), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n741), .A2(new_n269), .ZN(new_n1122));
  INV_X1    g0922(.A(G128), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .C1(new_n1123), .C2(new_n737), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1119), .B(new_n1124), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n288), .B1(new_n220), .B2(new_n742), .C1(new_n1126), .C2(new_n745), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT117), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1117), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n710), .B1(new_n1035), .B2(new_n786), .C1(new_n1129), .C2(new_n785), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n910), .B2(new_n720), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n709), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1111), .A2(new_n1133), .ZN(G378));
  NAND2_X1  g0934(.A1(new_n888), .A2(G330), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n866), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT40), .B1(new_n902), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n275), .A2(new_n822), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT55), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n313), .B(new_n1139), .ZN(new_n1140));
  XOR2_X1   g0940(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1140), .B(new_n1142), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1135), .A2(new_n1137), .A3(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1140), .B(new_n1141), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n674), .B1(new_n868), .B2(new_n887), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n867), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n913), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n911), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n867), .A2(new_n1146), .A3(new_n1145), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1151), .A3(new_n903), .A4(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1148), .A2(new_n1153), .A3(new_n709), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n710), .B1(G50), .B2(new_n786), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n409), .A2(G41), .ZN(new_n1156));
  INV_X1    g0956(.A(G41), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G50), .B(new_n1156), .C1(new_n284), .C2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n729), .A2(new_n486), .B1(new_n732), .B2(new_n358), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n742), .A2(new_n248), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G77), .B2(new_n758), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n227), .B2(new_n789), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1159), .B(new_n1162), .C1(G283), .C2(new_n746), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n941), .B1(new_n736), .B2(G116), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT118), .Z(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1165), .A3(new_n1156), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT58), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1158), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n284), .B(new_n1157), .C1(new_n742), .C2(new_n404), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G124), .B2(new_n746), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n789), .A2(new_n798), .B1(new_n732), .B2(new_n804), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT119), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n737), .A2(new_n1126), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n750), .A2(new_n269), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1123), .A2(new_n729), .B1(new_n741), .B2(new_n1118), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT59), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1170), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1176), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1168), .B1(new_n1167), .B2(new_n1166), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1155), .B1(new_n1181), .B2(new_n723), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1143), .B2(new_n721), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1154), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1091), .B1(new_n1132), .B2(new_n1109), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1148), .A2(new_n1153), .A3(KEYINPUT57), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1049), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1110), .A2(new_n1092), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1187), .B2(new_n1190), .ZN(G375));
  INV_X1    g0991(.A(new_n987), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1108), .A2(new_n1091), .A3(new_n1082), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1093), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n865), .A2(new_n721), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT121), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n289), .B1(new_n322), .B2(new_n742), .C1(new_n790), .C2(new_n729), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G107), .A2(new_n733), .B1(new_n746), .B2(G303), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n227), .B2(new_n741), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1037), .B1(new_n737), .B2(new_n762), .C1(new_n548), .C2(new_n789), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT123), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n457), .B(new_n1160), .C1(G137), .C2(new_n730), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n789), .A2(new_n1118), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n801), .A2(G50), .B1(G132), .B2(new_n736), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n732), .A2(new_n269), .B1(new_n745), .B2(new_n1123), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G159), .B2(new_n758), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n723), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n710), .B1(G68), .B2(new_n786), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT122), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1196), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1090), .B2(new_n709), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1194), .A2(new_n1215), .ZN(G381));
  INV_X1    g1016(.A(G375), .ZN(new_n1217));
  OR3_X1    g1017(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1218), .A2(G390), .A3(G381), .ZN(new_n1219));
  INV_X1    g1019(.A(G378), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(G387), .ZN(G407));
  NAND3_X1  g1022(.A1(new_n1217), .A2(new_n644), .A3(new_n1220), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G407), .A2(G213), .A3(new_n1223), .ZN(G409));
  INV_X1    g1024(.A(G390), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT124), .B1(G387), .B2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(G393), .B(new_n770), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n705), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1054), .B2(new_n995), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n708), .B1(new_n1230), .B2(new_n987), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n981), .A2(new_n984), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT109), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1231), .A2(new_n1234), .A3(new_n985), .A4(new_n986), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1235), .A2(new_n954), .A3(G390), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G390), .B1(new_n1235), .B2(new_n954), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n1226), .A2(new_n1228), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1237), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n954), .A3(G390), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(KEYINPUT124), .A3(new_n1227), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1184), .C1(new_n1187), .C2(new_n1190), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1188), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1184), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1220), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1245), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1193), .A2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1091), .A4(new_n1082), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1049), .A3(new_n1093), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1215), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n784), .A2(new_n811), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G384), .A2(new_n1215), .A3(new_n1254), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1245), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1259), .A2(G2897), .A3(new_n1245), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1245), .A2(G2897), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1257), .A2(new_n1258), .A3(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1243), .A2(new_n1261), .A3(new_n1269), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1250), .A2(new_n1260), .A3(new_n1274), .A4(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1269), .A2(new_n1276), .A3(KEYINPUT126), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1242), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1250), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1274), .B1(new_n1250), .B2(new_n1260), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT126), .B1(new_n1285), .B2(new_n1278), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1273), .B1(new_n1280), .B2(new_n1286), .ZN(G405));
  AND3_X1   g1087(.A1(new_n1238), .A2(new_n1241), .A3(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G375), .A2(new_n1220), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1289), .A2(new_n1259), .A3(new_n1246), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1259), .B1(new_n1289), .B2(new_n1246), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT127), .B1(new_n1238), .B2(new_n1241), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1288), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1242), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1238), .A2(new_n1241), .A3(KEYINPUT127), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1294), .A2(new_n1299), .ZN(G402));
endmodule


