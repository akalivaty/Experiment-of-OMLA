//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT73), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G137), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n193), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G119), .B(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(KEYINPUT72), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n202), .B(new_n204), .C1(G119), .C2(new_n203), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n198), .A2(new_n199), .B1(G110), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT16), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT74), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n198), .A2(new_n199), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n212), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n214), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n205), .A2(G110), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n216), .A2(new_n217), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n217), .B1(new_n216), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n196), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n216), .A2(new_n223), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n195), .B1(new_n227), .B2(KEYINPUT74), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n229), .B2(G902), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n190), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(new_n188), .A3(new_n190), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT0), .A3(G128), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT11), .A2(G134), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT11), .A2(G134), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(KEYINPUT64), .A2(G137), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT64), .A2(G137), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT65), .B1(new_n250), .B2(new_n243), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n245), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT64), .A2(G137), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n243), .A3(KEYINPUT65), .A4(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n247), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G131), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n243), .A3(new_n254), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n246), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n242), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  OR3_X1    g080(.A1(new_n266), .A2(KEYINPUT2), .A3(G113), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(KEYINPUT2), .B2(G113), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n267), .A2(new_n268), .B1(KEYINPUT2), .B2(G113), .ZN(new_n269));
  XNOR2_X1  g083(.A(G116), .B(G119), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n201), .A2(G116), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G119), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT68), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n271), .B1(new_n276), .B2(new_n269), .ZN(new_n277));
  AOI211_X1 g091(.A(G131), .B(new_n246), .C1(new_n261), .C2(new_n255), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n250), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n263), .B1(G134), .B2(G137), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n214), .A2(G143), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n203), .B1(new_n283), .B2(KEYINPUT1), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(new_n239), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n239), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n265), .A2(new_n277), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n277), .ZN(new_n290));
  INV_X1    g104(.A(new_n242), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n262), .A2(new_n263), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(new_n278), .ZN(new_n293));
  INV_X1    g107(.A(G143), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G146), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n283), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n284), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n264), .A2(new_n298), .A3(new_n282), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n290), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT28), .B1(new_n289), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n293), .A2(new_n290), .A3(new_n299), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G237), .A2(G953), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G210), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n307), .B(KEYINPUT27), .Z(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(G101), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n313), .B(new_n316), .C1(new_n265), .C2(new_n288), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n293), .A2(new_n314), .A3(new_n315), .A4(new_n299), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n290), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(new_n289), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n312), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n305), .A2(KEYINPUT29), .A3(new_n311), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n322), .B2(KEYINPUT71), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n321), .B(new_n323), .C1(KEYINPUT71), .C2(new_n322), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n311), .B1(new_n301), .B2(new_n304), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n319), .A2(new_n310), .A3(new_n289), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT69), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n317), .A2(new_n318), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n277), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n311), .A3(new_n302), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT31), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(KEYINPUT32), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n337), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT32), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT70), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n343), .A3(new_n337), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n238), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G210), .B1(G237), .B2(G902), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n201), .A3(G116), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n350), .A2(G113), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n270), .B(KEYINPUT68), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT81), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n355), .B(new_n351), .C1(new_n352), .C2(new_n349), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n357), .B2(G107), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G104), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(G107), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n358), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n357), .A2(G107), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n360), .A2(G104), .ZN(new_n366));
  OAI21_X1  g180(.A(G101), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n354), .A2(new_n356), .A3(new_n271), .A4(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G110), .B(G122), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT8), .Z(new_n371));
  OAI21_X1  g185(.A(new_n351), .B1(new_n349), .B2(new_n275), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n271), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n368), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n369), .A2(KEYINPUT83), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT83), .B1(new_n369), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n291), .A2(G125), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(G125), .B2(new_n297), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n191), .A2(G224), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n354), .A2(new_n356), .A3(new_n271), .A4(new_n374), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n358), .A2(new_n361), .A3(new_n363), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(G101), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(G101), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n364), .A3(KEYINPUT4), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n277), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(new_n370), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n383), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n188), .B1(new_n378), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n384), .A2(new_n391), .ZN(new_n396));
  INV_X1    g210(.A(new_n370), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n392), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n381), .B(KEYINPUT82), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n380), .B(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n396), .A2(new_n402), .A3(new_n397), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT84), .B(new_n348), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n348), .A2(KEYINPUT84), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n395), .A2(KEYINPUT85), .A3(new_n404), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n404), .A3(new_n347), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n406), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n294), .A2(G128), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n203), .A2(G143), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n415), .A2(new_n279), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT13), .B1(new_n294), .B2(G128), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n417), .A2(KEYINPUT93), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(KEYINPUT93), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n294), .A2(KEYINPUT13), .A3(G128), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n418), .A2(new_n414), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n416), .B1(new_n421), .B2(G134), .ZN(new_n422));
  INV_X1    g236(.A(G122), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT91), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G122), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n273), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n273), .A2(G122), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT92), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT91), .B(G122), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n431), .B(new_n428), .C1(new_n432), .C2(new_n273), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n430), .A2(G107), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(G107), .B1(new_n430), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n422), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n430), .A2(new_n433), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n360), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n428), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n424), .A2(new_n426), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G116), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n428), .A2(KEYINPUT14), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT94), .B1(new_n428), .B2(KEYINPUT14), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n439), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G107), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n415), .B(new_n279), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n438), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT9), .B(G234), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n449), .A2(new_n187), .A3(G953), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n436), .A2(new_n447), .A3(new_n450), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n188), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT95), .ZN(new_n456));
  INV_X1    g270(.A(G478), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n208), .A2(new_n210), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G146), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n215), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT18), .A2(G131), .ZN(new_n466));
  INV_X1    g280(.A(G237), .ZN(new_n467));
  AND4_X1   g281(.A1(G143), .A2(new_n467), .A3(new_n191), .A4(G214), .ZN(new_n468));
  AOI21_X1  g282(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n191), .A3(G214), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n294), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(KEYINPUT18), .A3(G131), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n462), .A2(new_n215), .A3(KEYINPUT86), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n465), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(KEYINPUT17), .B(G131), .C1(new_n468), .C2(new_n469), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n220), .A2(new_n213), .A3(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n468), .A2(new_n469), .A3(G131), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n263), .B1(new_n472), .B2(new_n473), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n484));
  AOI22_X1  g298(.A1(KEYINPUT88), .A2(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n220), .A2(new_n479), .A3(new_n486), .A4(new_n213), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n478), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G113), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n357), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n460), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n480), .A2(KEYINPUT88), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n483), .A2(new_n484), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  AND4_X1   g308(.A1(new_n460), .A2(new_n494), .A3(new_n490), .A4(new_n477), .ZN(new_n495));
  INV_X1    g309(.A(new_n483), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT19), .Z(new_n498));
  OAI211_X1 g312(.A(new_n213), .B(new_n496), .C1(new_n498), .C2(G146), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n499), .A2(new_n477), .ZN(new_n500));
  OAI22_X1  g314(.A1(new_n491), .A2(new_n495), .B1(new_n490), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n490), .B1(new_n499), .B2(new_n477), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n494), .A2(new_n477), .ZN(new_n506));
  INV_X1    g320(.A(new_n490), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT89), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n488), .A2(new_n460), .A3(new_n490), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n503), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT20), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n491), .A2(new_n495), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n494), .A2(new_n514), .A3(new_n477), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n494), .B2(new_n477), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(new_n490), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n188), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n504), .A2(new_n512), .B1(new_n518), .B2(G475), .ZN(new_n519));
  NAND2_X1  g333(.A1(G234), .A2(G237), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n520), .A2(G952), .A3(new_n191), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(G902), .A3(G953), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT96), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT21), .B(G898), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n459), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G214), .B1(G237), .B2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n297), .B(new_n374), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n292), .A2(new_n278), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT77), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(KEYINPUT77), .A2(KEYINPUT12), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n531), .C2(new_n532), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n258), .A2(new_n264), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n298), .A2(KEYINPUT10), .A3(new_n374), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT10), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n297), .B2(new_n368), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n291), .A2(new_n390), .A3(new_n388), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G110), .B(G140), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n191), .A2(G227), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n543), .A2(new_n547), .A3(new_n545), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n555), .A2(KEYINPUT78), .A3(new_n541), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT78), .B1(new_n555), .B2(new_n541), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n540), .A2(new_n554), .B1(new_n558), .B2(new_n552), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT80), .B(G469), .Z(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n188), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n549), .A2(new_n536), .A3(new_n539), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n552), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n549), .B(new_n553), .C1(new_n556), .C2(new_n557), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n566), .A3(new_n563), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G221), .B1(new_n449), .B2(G902), .ZN(new_n573));
  AND4_X1   g387(.A1(new_n412), .A2(new_n530), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n346), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(G101), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G3));
  NAND2_X1  g391(.A1(new_n336), .A2(new_n188), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G472), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n341), .A2(new_n579), .A3(new_n344), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n573), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n237), .ZN(new_n583));
  INV_X1    g397(.A(new_n404), .ZN(new_n584));
  OAI211_X1 g398(.A(KEYINPUT98), .B(new_n348), .C1(new_n584), .C2(new_n394), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n410), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT98), .B1(new_n405), .B2(new_n348), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n528), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n515), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n516), .A2(new_n490), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n589), .A2(new_n590), .B1(new_n508), .B2(new_n509), .ZN(new_n591));
  OAI21_X1  g405(.A(G475), .B1(new_n591), .B2(G902), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n510), .A2(KEYINPUT20), .A3(new_n511), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT99), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(KEYINPUT99), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n436), .A2(new_n447), .A3(new_n450), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n450), .B1(new_n436), .B2(new_n447), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n452), .A2(KEYINPUT99), .A3(new_n596), .A4(new_n453), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n457), .A2(G902), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT100), .B(G478), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n454), .B2(new_n188), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n595), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n526), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n583), .A2(new_n588), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(new_n459), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n592), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n235), .A2(new_n236), .A3(new_n526), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n504), .A2(KEYINPUT102), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT103), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(KEYINPUT103), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n512), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n594), .A3(new_n622), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n619), .B(new_n620), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n348), .B1(new_n584), .B2(new_n394), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n410), .A3(new_n585), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n628), .A2(new_n582), .A3(new_n528), .A4(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  INV_X1    g449(.A(new_n580), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n195), .A2(KEYINPUT36), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n227), .B(new_n637), .Z(new_n638));
  NOR3_X1   g452(.A1(new_n638), .A2(G902), .A3(new_n189), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n234), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n574), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  NAND2_X1  g458(.A1(new_n339), .A2(new_n345), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n572), .A2(new_n573), .A3(new_n641), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n588), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT104), .B(G900), .Z(new_n648));
  AOI21_X1  g462(.A(new_n521), .B1(new_n523), .B2(new_n648), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n649), .B(new_n619), .C1(new_n625), .C2(new_n627), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XOR2_X1   g466(.A(new_n649), .B(KEYINPUT39), .Z(new_n653));
  NAND3_X1  g467(.A1(new_n572), .A2(new_n573), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n459), .A2(new_n519), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n640), .A3(new_n528), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n654), .B2(KEYINPUT40), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n412), .B(KEYINPUT38), .ZN(new_n659));
  INV_X1    g473(.A(new_n320), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n311), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n289), .A2(new_n300), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n661), .B(new_n188), .C1(new_n311), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n345), .A2(new_n338), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n655), .A2(new_n658), .A3(new_n659), .A4(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n294), .ZN(G45));
  NOR2_X1   g485(.A1(new_n611), .A2(new_n649), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n645), .A2(new_n647), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  OAI21_X1  g488(.A(G469), .B1(new_n559), .B2(G902), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n562), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n573), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n588), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n238), .A2(new_n613), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n645), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND3_X1  g497(.A1(new_n645), .A2(new_n628), .A3(new_n679), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  NOR2_X1   g499(.A1(new_n527), .A2(new_n640), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n645), .A2(new_n679), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT106), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n645), .A2(new_n689), .A3(new_n679), .A4(new_n686), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  OAI21_X1  g506(.A(new_n329), .B1(new_n328), .B2(new_n327), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n337), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n237), .A2(new_n579), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n656), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n588), .A2(new_n696), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n573), .A2(new_n562), .A3(new_n526), .A4(new_n675), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(new_n697), .A3(KEYINPUT107), .A4(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n698), .A2(new_n528), .A3(new_n632), .A4(new_n656), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n237), .A2(new_n579), .A3(new_n694), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(G122), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G24));
  AND2_X1   g520(.A1(new_n579), .A2(new_n694), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n707), .A2(new_n641), .A3(new_n672), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n679), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  NOR2_X1   g524(.A1(new_n412), .A2(new_n529), .ZN(new_n711));
  INV_X1    g525(.A(new_n573), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n565), .A2(new_n566), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(G902), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n712), .B1(new_n715), .B2(new_n562), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n672), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n325), .A2(new_n338), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT32), .B1(new_n336), .B2(new_n337), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n237), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n346), .A2(new_n717), .A3(new_n726), .A4(new_n672), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT110), .B(G131), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G33));
  NAND3_X1  g545(.A1(new_n346), .A2(new_n650), .A3(new_n717), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(G134), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G36));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n605), .A2(new_n609), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n604), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n601), .B2(new_n602), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT112), .B1(new_n740), .B2(new_n608), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n736), .B1(new_n742), .B2(new_n595), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n736), .B1(new_n605), .B2(new_n609), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n512), .A2(new_n504), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n592), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n744), .B1(new_n519), .B2(new_n745), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n580), .A2(KEYINPUT44), .A3(new_n641), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n711), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n580), .A2(new_n641), .A3(new_n749), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n751), .B1(new_n750), .B2(new_n711), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n735), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n750), .A2(new_n711), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT114), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(KEYINPUT115), .A3(new_n752), .A4(new_n755), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  OAI21_X1  g576(.A(G469), .B1(new_n713), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n568), .A2(new_n569), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(new_n762), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n571), .A2(new_n188), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT46), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n765), .B2(new_n766), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n562), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n573), .A3(new_n653), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n758), .A2(new_n761), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT116), .B(G137), .Z(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G39));
  NAND3_X1  g590(.A1(new_n711), .A2(new_n672), .A3(new_n238), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n645), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n771), .A2(new_n573), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n573), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n207), .ZN(G42));
  AND3_X1   g598(.A1(new_n704), .A2(new_n684), .A3(new_n681), .ZN(new_n785));
  INV_X1    g599(.A(new_n746), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n611), .B1(new_n619), .B2(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n412), .A2(new_n528), .A3(new_n526), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n582), .A2(new_n237), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n575), .A2(new_n642), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n711), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n625), .A2(new_n627), .ZN(new_n792));
  INV_X1    g606(.A(new_n649), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n459), .A2(new_n592), .A3(new_n793), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n791), .A2(new_n792), .A3(new_n646), .A4(new_n794), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n795), .A2(new_n645), .B1(new_n708), .B2(new_n717), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n785), .A2(new_n790), .A3(new_n691), .A4(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n728), .B(new_n732), .C1(new_n725), .C2(new_n726), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n641), .A2(new_n649), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n665), .A2(new_n697), .A3(new_n716), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n651), .A2(new_n709), .A3(new_n673), .A4(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(KEYINPUT119), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(KEYINPUT119), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n805), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n800), .A2(new_n801), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n807), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n804), .A2(KEYINPUT119), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n806), .A2(KEYINPUT52), .A3(new_n807), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n799), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n812), .B(KEYINPUT54), .C1(new_n818), .C2(new_n801), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n801), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n790), .A2(new_n796), .A3(KEYINPUT53), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n798), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n785), .A2(new_n691), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n810), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n659), .A2(new_n528), .A3(new_n678), .ZN(new_n830));
  INV_X1    g644(.A(new_n749), .ZN(new_n831));
  INV_X1    g645(.A(new_n521), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n831), .A2(new_n702), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT50), .Z(new_n835));
  NAND3_X1  g649(.A1(new_n711), .A2(new_n573), .A3(new_n677), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n836), .A2(new_n665), .A3(new_n238), .A4(new_n832), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n595), .A2(new_n610), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n836), .A2(new_n832), .A3(new_n831), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n707), .A2(new_n641), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n837), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n781), .B(new_n782), .C1(new_n573), .C2(new_n676), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n711), .A3(new_n833), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n835), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n723), .A2(new_n724), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n839), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT48), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n833), .A2(new_n679), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(G952), .A3(new_n191), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n612), .B2(new_n837), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n846), .A2(new_n847), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n829), .A2(new_n854), .B1(G952), .B2(G953), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n237), .A2(new_n573), .A3(new_n528), .A4(new_n610), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n676), .A2(KEYINPUT49), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n595), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(KEYINPUT49), .B2(new_n676), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n665), .A3(new_n659), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT117), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n855), .A2(new_n861), .ZN(G75));
  NOR2_X1   g676(.A1(new_n191), .A2(G952), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n188), .B1(new_n820), .B2(new_n826), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT56), .B1(new_n865), .B2(G210), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n866), .B2(KEYINPUT121), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n820), .A2(new_n826), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(G902), .ZN(new_n870));
  INV_X1    g684(.A(G210), .ZN(new_n871));
  OAI211_X1 g685(.A(KEYINPUT121), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n399), .A2(new_n403), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(new_n401), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT55), .Z(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n866), .A2(KEYINPUT121), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n867), .B1(new_n876), .B2(new_n878), .ZN(G51));
  XNOR2_X1  g693(.A(new_n766), .B(KEYINPUT57), .ZN(new_n880));
  INV_X1    g694(.A(new_n828), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n827), .B1(new_n820), .B2(new_n826), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n560), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n865), .A2(new_n765), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n863), .B1(new_n884), .B2(new_n885), .ZN(G54));
  NAND2_X1  g700(.A1(KEYINPUT58), .A2(G475), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT122), .Z(new_n888));
  NOR2_X1   g702(.A1(new_n870), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n864), .B1(new_n889), .B2(new_n501), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n870), .A2(new_n510), .A3(new_n888), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n603), .B1(new_n829), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n603), .B(new_n895), .C1(new_n881), .C2(new_n882), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n864), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT60), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n869), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n863), .B1(new_n903), .B2(new_n229), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n904), .B(KEYINPUT61), .C1(new_n638), .C2(new_n903), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n638), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n901), .B1(new_n820), .B2(new_n826), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n864), .B1(new_n908), .B2(new_n230), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n910), .ZN(G66));
  INV_X1    g725(.A(new_n524), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n191), .B1(new_n912), .B2(G224), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n785), .A2(new_n790), .A3(new_n691), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n913), .B1(new_n915), .B2(new_n191), .ZN(new_n916));
  INV_X1    g730(.A(G898), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n873), .B1(new_n917), .B2(G953), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n916), .B(new_n918), .ZN(G69));
  XOR2_X1   g733(.A(new_n331), .B(new_n498), .Z(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(G953), .ZN(new_n921));
  INV_X1    g735(.A(new_n654), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n346), .A2(new_n922), .A3(new_n711), .A4(new_n787), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n783), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n709), .A2(new_n651), .A3(new_n673), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n668), .A2(new_n669), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n668), .A2(KEYINPUT62), .A3(new_n925), .A4(new_n669), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(KEYINPUT123), .A3(new_n774), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT123), .B1(new_n930), .B2(new_n774), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n921), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(KEYINPUT124), .B(KEYINPUT127), .Z(new_n935));
  AOI21_X1  g749(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n191), .A2(G900), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n771), .A2(new_n573), .A3(new_n653), .A4(new_n697), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n724), .B2(new_n723), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n798), .A2(new_n783), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n774), .A2(KEYINPUT125), .A3(new_n925), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT125), .B1(new_n774), .B2(new_n925), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n944), .B2(new_n191), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n920), .B1(new_n945), .B2(KEYINPUT126), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n947), .B(new_n938), .C1(new_n944), .C2(new_n191), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n934), .B(new_n937), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n938), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n783), .A2(new_n940), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n727), .A3(new_n728), .A4(new_n732), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n774), .A2(new_n925), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n774), .A2(KEYINPUT125), .A3(new_n925), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n958), .B2(G953), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n947), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n920), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n937), .B1(new_n962), .B2(new_n934), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n950), .A2(new_n963), .ZN(G72));
  OAI21_X1  g778(.A(new_n812), .B1(new_n818), .B2(new_n801), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  NOR2_X1   g781(.A1(new_n320), .A2(new_n311), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n327), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n864), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n933), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n914), .A3(new_n931), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n661), .B1(new_n972), .B2(new_n967), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n958), .A2(new_n914), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n311), .B(new_n660), .C1(new_n974), .C2(new_n967), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(G57));
endmodule


