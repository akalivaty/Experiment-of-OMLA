//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT69), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT2), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(G261));
  INV_X1    g035(.A(G261), .ZN(G325));
  INV_X1    g036(.A(new_n459), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n456), .A2(G567), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT70), .A3(G137), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n479), .A2(new_n474), .ZN(new_n480));
  INV_X1    g055(.A(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT71), .Z(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n478), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NOR2_X1   g061(.A1(new_n469), .A2(new_n474), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n470), .A2(G136), .ZN(new_n489));
  NOR2_X1   g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n488), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n469), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n496), .A2(G2105), .B1(G102), .B2(new_n482), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n467), .B2(new_n468), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n502), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n473), .A2(new_n504), .A3(new_n499), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT73), .B(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT76), .A3(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT73), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT73), .A2(G651), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n519), .B(KEYINPUT6), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n525), .A2(G88), .A3(new_n515), .A4(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT6), .B1(new_n521), .B2(new_n522), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n530));
  AND2_X1   g105(.A1(G50), .A2(G543), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n530), .A2(new_n527), .A3(new_n523), .A4(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT77), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n537), .B(new_n528), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n518), .B1(new_n536), .B2(new_n538), .ZN(G166));
  NAND2_X1  g114(.A1(G63), .A2(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n530), .A2(new_n527), .A3(new_n523), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n530), .A2(KEYINPUT78), .A3(new_n527), .A4(new_n523), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G543), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G51), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n544), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  AND4_X1   g128(.A1(new_n515), .A2(new_n530), .A3(new_n527), .A4(new_n523), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n556));
  INV_X1    g131(.A(new_n514), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT76), .B1(new_n513), .B2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G64), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n509), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n554), .A2(G90), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n548), .A2(G52), .A3(G543), .A4(new_n549), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(G301));
  INV_X1    g140(.A(G301), .ZN(G171));
  NAND4_X1  g141(.A1(new_n548), .A2(G43), .A3(G543), .A4(new_n549), .ZN(new_n567));
  OAI211_X1 g142(.A(G56), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n568));
  NAND2_X1  g143(.A1(G68), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n509), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n554), .B2(G81), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT80), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(new_n580), .ZN(G188));
  NAND4_X1  g156(.A1(new_n530), .A2(new_n515), .A3(new_n527), .A4(new_n523), .ZN(new_n582));
  INV_X1    g157(.A(G91), .ZN(new_n583));
  OR3_X1    g158(.A1(new_n582), .A2(KEYINPUT81), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT81), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G65), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n559), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n584), .A2(new_n585), .B1(G651), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n548), .A2(G53), .A3(G543), .A4(new_n549), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n590), .A2(KEYINPUT9), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(KEYINPUT9), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(G299));
  INV_X1    g168(.A(new_n518), .ZN(new_n594));
  INV_X1    g169(.A(new_n538), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n525), .A2(new_n596), .A3(new_n527), .A4(new_n531), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n537), .B1(new_n599), .B2(new_n528), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(new_n595), .B2(new_n600), .ZN(G303));
  OAI21_X1  g176(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT82), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n554), .A2(G87), .ZN(new_n604));
  INV_X1    g179(.A(G49), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n550), .C2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT83), .ZN(G288));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n608));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n559), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G73), .A2(G543), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n515), .A2(KEYINPUT84), .A3(G61), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n562), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n515), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(new_n541), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(G305));
  NAND2_X1  g192(.A1(G72), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G60), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n559), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n554), .A2(G85), .B1(new_n620), .B2(new_n562), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n548), .A2(G47), .A3(G543), .A4(new_n549), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(G290));
  NAND2_X1  g198(.A1(G301), .A2(G868), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n554), .A2(KEYINPUT10), .A3(G92), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n582), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n548), .A2(G54), .A3(G543), .A4(new_n549), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(new_n526), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n624), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n624), .B1(new_n634), .B2(G868), .ZN(G321));
  NAND2_X1  g211(.A1(G286), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(G299), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G280));
  XNOR2_X1  g214(.A(G280), .B(KEYINPUT85), .ZN(G297));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n634), .B1(new_n641), .B2(G860), .ZN(G148));
  NAND2_X1  g217(.A1(new_n634), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G868), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n483), .A2(new_n473), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT13), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n487), .A2(G123), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n470), .A2(G135), .ZN(new_n652));
  NOR2_X1   g227(.A1(G99), .A2(G2105), .ZN(new_n653));
  OAI21_X1  g228(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n651), .B(new_n652), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(G2096), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1341), .B(G1348), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2427), .B(G2430), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT86), .B(KEYINPUT14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n663), .B(new_n669), .Z(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(G14), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT87), .ZN(new_n673));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(KEYINPUT17), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(G2072), .A2(G2078), .ZN(new_n681));
  OAI22_X1  g256(.A1(new_n675), .A2(new_n679), .B1(new_n444), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n686), .A2(new_n687), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n692), .B1(KEYINPUT20), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n689), .A2(new_n691), .A3(new_n693), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n695), .B(new_n696), .C1(KEYINPUT20), .C2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  AND2_X1   g279(.A1(KEYINPUT89), .A2(G29), .ZN(new_n705));
  NOR2_X1   g280(.A1(KEYINPUT89), .A2(G29), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G35), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G162), .B2(new_n708), .ZN(new_n710));
  MUX2_X1   g285(.A(new_n709), .B(new_n710), .S(KEYINPUT98), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT29), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G2090), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n483), .A2(G105), .ZN(new_n714));
  AOI22_X1  g289(.A1(G129), .A2(new_n487), .B1(new_n470), .B2(G141), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G29), .B2(G32), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n655), .A2(new_n708), .ZN(new_n725));
  INV_X1    g300(.A(G28), .ZN(new_n726));
  OR3_X1    g301(.A1(new_n726), .A2(KEYINPUT96), .A3(KEYINPUT30), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(KEYINPUT30), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT96), .B1(new_n726), .B2(KEYINPUT30), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n723), .A2(new_n724), .A3(new_n725), .A4(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(G29), .A2(G33), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n482), .A2(G103), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT25), .ZN(new_n736));
  NAND2_X1  g311(.A1(G115), .A2(G2104), .ZN(new_n737));
  INV_X1    g312(.A(G127), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n469), .B2(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n739), .A2(G2105), .B1(new_n470), .B2(G139), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(new_n728), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(new_n442), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n442), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n732), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G1961), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n708), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n708), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2078), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G34), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n708), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n485), .B2(new_n728), .ZN(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n746), .A2(new_n750), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G11), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n747), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n747), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n749), .A2(G1961), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n762), .A2(new_n763), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT97), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n747), .A2(G20), .ZN(new_n771));
  OAI211_X1 g346(.A(KEYINPUT23), .B(new_n771), .C1(new_n638), .C2(new_n747), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT23), .B2(new_n771), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  AND4_X1   g349(.A1(new_n768), .A2(new_n746), .A3(new_n750), .A4(new_n761), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n775), .A2(new_n776), .A3(new_n763), .A4(new_n767), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n573), .A2(new_n747), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n747), .B2(G19), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(G1341), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n747), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n634), .B2(new_n747), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1348), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n780), .A2(G1341), .ZN(new_n785));
  AOI21_X1  g360(.A(KEYINPUT28), .B1(new_n708), .B2(G26), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n708), .A2(KEYINPUT28), .A3(G26), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n487), .A2(G128), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n470), .A2(G140), .ZN(new_n790));
  NOR2_X1   g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(new_n474), .B2(G116), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n786), .B(new_n788), .C1(new_n793), .C2(G29), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n781), .A2(new_n784), .A3(new_n785), .A4(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n770), .A2(new_n774), .A3(new_n777), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n747), .A2(G23), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n799), .B1(new_n802), .B2(new_n747), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT33), .B(G1976), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n807));
  NOR2_X1   g382(.A1(G166), .A2(new_n747), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n747), .B2(G22), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT93), .B(G1971), .Z(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n747), .A2(G6), .ZN(new_n812));
  INV_X1    g387(.A(G305), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n747), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT32), .B(G1981), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n809), .B2(new_n810), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n806), .A2(new_n807), .A3(new_n811), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n811), .A2(new_n817), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT34), .B1(new_n819), .B2(new_n805), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n487), .A2(G119), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n470), .A2(G131), .ZN(new_n822));
  NOR2_X1   g397(.A1(G95), .A2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(new_n474), .B2(G107), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G25), .B(new_n825), .S(new_n707), .Z(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT90), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G16), .A2(G24), .ZN(new_n830));
  XOR2_X1   g405(.A(G290), .B(KEYINPUT91), .Z(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(G16), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(G1986), .Z(new_n833));
  NAND4_X1  g408(.A1(new_n818), .A2(new_n820), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n836));
  AOI211_X1 g411(.A(new_n713), .B(new_n798), .C1(new_n835), .C2(new_n836), .ZN(G311));
  AOI21_X1  g412(.A(new_n798), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  INV_X1    g413(.A(new_n713), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(G150));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n559), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n554), .A2(G93), .B1(new_n843), .B2(new_n562), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n548), .A2(G55), .A3(G543), .A4(new_n549), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n567), .A3(new_n571), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n572), .A2(new_n845), .A3(new_n844), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n633), .A2(new_n641), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n856), .A2(KEYINPUT99), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(KEYINPUT99), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n854), .A2(new_n855), .ZN(new_n859));
  NOR4_X1   g434(.A1(new_n857), .A2(new_n858), .A3(G860), .A4(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n848), .B1(new_n862), .B2(new_n863), .ZN(G145));
  AND3_X1   g439(.A1(new_n503), .A2(KEYINPUT101), .A3(new_n505), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT101), .B1(new_n503), .B2(new_n505), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n497), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n793), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n718), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n648), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n487), .A2(G130), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT102), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n470), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n741), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n825), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n870), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n485), .B(G162), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(new_n655), .Z(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OR3_X1    g457(.A1(new_n879), .A2(KEYINPUT103), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT103), .B1(new_n879), .B2(new_n882), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n879), .A2(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g463(.A1(G299), .A2(new_n634), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n590), .B(KEYINPUT9), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n589), .A3(new_n633), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT41), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n643), .B(new_n851), .Z(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n889), .A2(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n889), .A2(KEYINPUT104), .A3(new_n891), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n895), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n896), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n897), .B1(new_n896), .B2(new_n902), .ZN(new_n904));
  INV_X1    g479(.A(G290), .ZN(new_n905));
  NAND2_X1  g480(.A1(G303), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n536), .A2(new_n538), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n594), .A3(G290), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n906), .A2(G305), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(G305), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n909), .A2(new_n910), .A3(new_n802), .ZN(new_n911));
  INV_X1    g486(.A(new_n802), .ZN(new_n912));
  INV_X1    g487(.A(new_n908), .ZN(new_n913));
  NOR2_X1   g488(.A1(G166), .A2(G290), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n813), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n906), .A2(G305), .A3(new_n908), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n903), .A2(new_n904), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n903), .B2(new_n904), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(G868), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G868), .B1(new_n844), .B2(new_n845), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(KEYINPUT105), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(KEYINPUT105), .B2(new_n921), .ZN(G295));
  OAI21_X1  g499(.A(new_n923), .B1(KEYINPUT105), .B2(new_n921), .ZN(G331));
  INV_X1    g500(.A(new_n893), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n849), .A2(new_n850), .A3(G301), .ZN(new_n928));
  AOI21_X1  g503(.A(G301), .B1(new_n849), .B2(new_n850), .ZN(new_n929));
  OAI21_X1  g504(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n851), .A2(G171), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n849), .A2(new_n850), .A3(G301), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G168), .A3(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n926), .A2(new_n927), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n930), .A2(new_n933), .A3(new_n898), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n918), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n928), .A2(new_n929), .A3(G286), .ZN(new_n939));
  AOI21_X1  g514(.A(G168), .B1(new_n931), .B2(new_n932), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n939), .A2(new_n940), .B1(new_n892), .B2(new_n893), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n802), .B1(new_n909), .B2(new_n910), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n915), .A2(new_n912), .A3(new_n916), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n930), .A2(new_n933), .A3(new_n898), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n938), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  AND4_X1   g525(.A1(new_n900), .A2(new_n930), .A3(new_n933), .A4(new_n901), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n951), .A2(new_n934), .B1(new_n911), .B2(new_n917), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n934), .B2(new_n935), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n941), .A2(new_n955), .A3(new_n944), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n954), .B(new_n956), .C1(new_n911), .C2(new_n917), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(new_n947), .A3(new_n938), .A4(new_n946), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n938), .A2(new_n946), .A3(new_n947), .A4(new_n952), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT108), .B1(new_n960), .B2(KEYINPUT43), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n953), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n960), .B2(KEYINPUT43), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n945), .B(new_n937), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(new_n950), .A3(new_n947), .A4(new_n957), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n964), .B2(new_n966), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n962), .A2(KEYINPUT44), .B1(new_n968), .B2(new_n969), .ZN(G397));
  NAND2_X1  g545(.A1(new_n482), .A2(G102), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n473), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(new_n474), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n506), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT101), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(G1384), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n478), .A2(new_n480), .A3(new_n484), .A4(G40), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n793), .B(new_n795), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n719), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT125), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n982), .B2(G1996), .ZN(new_n987));
  INV_X1    g562(.A(new_n982), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(KEYINPUT46), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n985), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT126), .Z(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT48), .Z(new_n996));
  XNOR2_X1  g571(.A(new_n825), .B(new_n827), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT110), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n718), .B(new_n989), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n983), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n988), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n825), .A2(new_n827), .ZN(new_n1003));
  OAI22_X1  g578(.A1(new_n1000), .A2(new_n1003), .B1(G2067), .B2(new_n793), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n988), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n993), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT112), .B1(new_n977), .B2(G1384), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n867), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n980), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1015), .B1(KEYINPUT115), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1016), .A2(new_n1023), .A3(KEYINPUT49), .A4(new_n1017), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1019), .A2(KEYINPUT116), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(KEYINPUT115), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(new_n1022), .A3(new_n1027), .A4(new_n1024), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n800), .B2(new_n801), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1032), .B2(new_n1015), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n1032), .C2(new_n1015), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1025), .A2(new_n1030), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(G166), .B2(new_n1014), .ZN(new_n1039));
  NAND3_X1  g614(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT113), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n977), .A2(KEYINPUT112), .A3(G1384), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1010), .B1(new_n867), .B2(new_n1011), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n497), .B2(new_n506), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n981), .B1(new_n1047), .B2(new_n1043), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(G2090), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1052));
  INV_X1    g627(.A(new_n506), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1011), .B1(new_n1053), .B2(new_n973), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1052), .A2(new_n981), .A3(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(G1971), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1014), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1042), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(new_n1027), .C1(new_n1031), .C2(new_n912), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1037), .A2(new_n1060), .A3(KEYINPUT63), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT50), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1064), .A2(G2084), .A3(new_n1048), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1009), .A2(new_n1055), .A3(new_n1012), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n980), .B1(new_n1047), .B2(KEYINPUT45), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1966), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G286), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1059), .B2(new_n1041), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1008), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1037), .A2(new_n1059), .A3(new_n1062), .A4(new_n1042), .ZN(new_n1073));
  AOI211_X1 g648(.A(G1976), .B(G288), .C1(new_n1025), .C2(new_n1030), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1016), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1027), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1009), .A2(KEYINPUT50), .A3(new_n1012), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT117), .B1(new_n1054), .B2(KEYINPUT50), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1047), .A2(new_n1080), .A3(new_n1043), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1082), .A3(new_n981), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1057), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G299), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n890), .A2(KEYINPUT57), .A3(new_n589), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT58), .B(G1341), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1052), .A2(new_n981), .A3(new_n1056), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1013), .A2(new_n1098), .B1(new_n1099), .B2(G1996), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n573), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1096), .A2(new_n1097), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1013), .A2(new_n795), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1348), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1112), .B2(new_n634), .ZN(new_n1113));
  INV_X1    g688(.A(G1348), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1064), .B2(new_n1048), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1105), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1116), .A2(KEYINPUT120), .A3(new_n633), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1109), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1112), .A2(new_n1110), .A3(new_n634), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT120), .B1(new_n1116), .B2(new_n633), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(KEYINPUT60), .A4(new_n1108), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1092), .A2(KEYINPUT119), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1088), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1095), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1104), .A2(new_n1118), .A3(new_n1121), .A4(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1095), .B(new_n634), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1128), .A2(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n766), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1046), .A2(new_n1049), .A3(new_n759), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1014), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(G286), .A2(G8), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT121), .Z(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT51), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT122), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1069), .A2(new_n1141), .A3(new_n1138), .A4(new_n1135), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(G8), .B(G286), .C1(new_n1065), .C2(new_n1068), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n1146));
  INV_X1    g721(.A(G1961), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1057), .A2(new_n443), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1050), .A2(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(G2078), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1066), .A2(new_n1067), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(G301), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1146), .B1(new_n1153), .B2(KEYINPUT124), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n981), .B1(new_n978), .B2(KEYINPUT45), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1155), .A2(KEYINPUT123), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(KEYINPUT123), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1052), .A3(new_n1151), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1150), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(G171), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1150), .A2(new_n1161), .A3(G301), .A4(new_n1152), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1154), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(G171), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1158), .A2(new_n1150), .A3(G301), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1146), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1145), .A2(new_n1163), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1130), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1070), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1145), .A2(KEYINPUT62), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1143), .A2(new_n1173), .A3(new_n1144), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1172), .A2(G171), .A3(new_n1164), .A4(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1170), .A2(new_n1171), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1037), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1058), .B1(new_n1083), .B2(G2090), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1041), .B1(G8), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1077), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(G290), .B(G1986), .Z(new_n1182));
  OAI21_X1  g757(.A(new_n1001), .B1(new_n982), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT111), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1007), .B1(new_n1181), .B2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g760(.A1(G229), .A2(G401), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n885), .B2(new_n886), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n953), .A2(new_n959), .A3(new_n961), .ZN(new_n1189));
  NOR2_X1   g763(.A1(G227), .A2(new_n465), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(G225));
  INV_X1    g765(.A(G225), .ZN(G308));
endmodule


