//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  OR2_X1    g004(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n204), .B(new_n211), .C1(new_n208), .C2(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G226gat), .A2(G233gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n217), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n220), .A2(new_n221), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(new_n223), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT65), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n229), .A2(new_n233), .A3(new_n234), .A4(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT27), .B(G183gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT28), .B1(new_n243), .B2(new_n219), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT27), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G183gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n245), .B2(new_n247), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(G190gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n244), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n256), .A2(new_n237), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT70), .B1(new_n235), .B2(new_n255), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n259), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n225), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n242), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n225), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n266), .A2(new_n267), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n230), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n240), .B1(new_n272), .B2(KEYINPUT68), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n230), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n234), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT75), .B1(new_n264), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n236), .A2(new_n234), .A3(new_n239), .A4(new_n237), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n224), .A2(new_n228), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(KEYINPUT65), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n246), .A2(G183gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT69), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n253), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n243), .A2(new_n219), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n252), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n257), .A2(new_n261), .B1(G183gat), .B2(G190gat), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n280), .A2(new_n229), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n272), .A2(KEYINPUT68), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n275), .A3(new_n241), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT25), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n216), .B1(new_n277), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n216), .ZN(new_n297));
  AOI211_X1 g096(.A(KEYINPUT29), .B(new_n297), .C1(new_n290), .C2(new_n293), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n215), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(new_n297), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n277), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n215), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n290), .A2(new_n293), .A3(new_n297), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G8gat), .B(G36gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(G64gat), .B(G92gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  NAND3_X1  g108(.A1(new_n299), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n299), .A2(KEYINPUT77), .A3(new_n306), .A4(new_n309), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT79), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n312), .A2(new_n317), .A3(new_n313), .A4(new_n314), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n309), .B1(new_n299), .B2(new_n306), .ZN(new_n319));
  INV_X1    g118(.A(new_n310), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT30), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n316), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G127gat), .ZN(new_n324));
  INV_X1    g123(.A(G127gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(KEYINPUT1), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n331), .B(new_n333), .C1(new_n332), .C2(G120gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n332), .A2(G120gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n330), .A2(G113gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n328), .A2(new_n334), .B1(new_n338), .B2(new_n327), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n264), .B2(new_n276), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n328), .A2(new_n334), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n327), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n290), .A2(new_n293), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G227gat), .ZN(new_n345));
  INV_X1    g144(.A(G233gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n349));
  XOR2_X1   g148(.A(G15gat), .B(G43gat), .Z(new_n350));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT34), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n344), .ZN(new_n357));
  INV_X1    g156(.A(new_n347), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI211_X1 g158(.A(KEYINPUT34), .B(new_n347), .C1(new_n340), .C2(new_n344), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n349), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(new_n358), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT34), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n357), .A2(new_n356), .A3(new_n358), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n348), .A2(new_n354), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n353), .ZN(new_n369));
  INV_X1    g168(.A(new_n349), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n361), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT81), .ZN(new_n379));
  INV_X1    g178(.A(new_n374), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  INV_X1    g180(.A(G155gat), .ZN(new_n382));
  INV_X1    g181(.A(G162gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n380), .B1(new_n384), .B2(new_n375), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n374), .A3(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(G141gat), .A2(G148gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n387), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n389), .A2(new_n382), .A3(new_n383), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n374), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n301), .B1(new_n213), .B2(new_n214), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n396), .B1(new_n386), .B2(new_n385), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n378), .A2(KEYINPUT81), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n404), .B(new_n400), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n215), .B1(new_n407), .B2(new_n300), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n408), .B2(KEYINPUT86), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n410), .B(new_n215), .C1(new_n300), .C2(new_n407), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n373), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n400), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n378), .A2(KEYINPUT81), .B1(new_n395), .B2(new_n392), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n387), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n215), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n417), .B2(new_n404), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n373), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n407), .A2(new_n300), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n304), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT87), .B1(new_n412), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT85), .ZN(new_n426));
  XOR2_X1   g225(.A(G78gat), .B(G106gat), .Z(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(G22gat), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n418), .A2(new_n373), .A3(new_n408), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n301), .B1(new_n415), .B2(new_n404), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n410), .B1(new_n433), .B2(new_n215), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n408), .A2(KEYINPUT86), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n403), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n432), .B1(new_n436), .B2(new_n373), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n431), .B(new_n428), .C1(new_n437), .C2(KEYINPUT87), .ZN(new_n438));
  INV_X1    g237(.A(new_n214), .ZN(new_n439));
  AND2_X1   g238(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n441));
  OAI21_X1  g240(.A(G211gat), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n443));
  NOR2_X1   g242(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n211), .B1(new_n446), .B2(new_n204), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n300), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n415), .B1(new_n448), .B2(new_n404), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n422), .B2(new_n410), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n420), .B1(new_n450), .B2(new_n435), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n451), .A2(new_n452), .A3(new_n432), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n430), .A2(new_n438), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n430), .B2(new_n438), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n372), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n343), .A2(KEYINPUT83), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n339), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n401), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n397), .A2(new_n339), .A3(new_n400), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT84), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n415), .A2(new_n464), .A3(new_n339), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n457), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT4), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n401), .A2(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n472), .A2(new_n407), .A3(new_n458), .A4(new_n460), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n339), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n471), .A2(new_n473), .A3(new_n474), .A4(new_n467), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n407), .A2(new_n458), .A3(new_n460), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n415), .A2(new_n404), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n457), .B(new_n467), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n470), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT0), .ZN(new_n487));
  XNOR2_X1  g286(.A(G57gat), .B(G85gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n484), .A3(new_n489), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n485), .A2(KEYINPUT6), .A3(new_n490), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n322), .A2(new_n456), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n202), .B(new_n203), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n322), .A2(new_n456), .A3(KEYINPUT92), .A4(new_n496), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n316), .A2(new_n496), .A3(new_n318), .A4(new_n321), .ZN(new_n501));
  INV_X1    g300(.A(new_n453), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n452), .B1(new_n451), .B2(new_n432), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n431), .B1(new_n503), .B2(new_n428), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n424), .A2(G22gat), .A3(new_n429), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n430), .A2(new_n438), .A3(new_n453), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n506), .A2(new_n371), .A3(new_n364), .A4(new_n507), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n501), .A2(new_n508), .A3(new_n498), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT35), .B(new_n500), .C1(new_n509), .C2(KEYINPUT92), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n312), .A2(new_n313), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n309), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n319), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n303), .A2(new_n305), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n215), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n296), .A2(new_n298), .ZN(new_n518));
  OAI211_X1 g317(.A(KEYINPUT90), .B(new_n517), .C1(new_n518), .C2(new_n215), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n296), .A2(new_n215), .A3(new_n298), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n513), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT38), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n319), .A2(new_n514), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n513), .B1(new_n299), .B2(new_n306), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n511), .B(new_n512), .C1(new_n524), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n454), .A2(new_n455), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n482), .A2(new_n473), .A3(new_n483), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n468), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(KEYINPUT39), .C1(new_n468), .C2(new_n466), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n534), .A3(new_n468), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n535), .A2(new_n536), .A3(new_n489), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n535), .B2(new_n489), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT40), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n533), .B(KEYINPUT40), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n491), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n529), .B(new_n530), .C1(new_n322), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n369), .A2(new_n370), .A3(new_n361), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n370), .B1(new_n369), .B2(new_n361), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n364), .A2(new_n545), .A3(new_n546), .A4(new_n371), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n530), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(new_n501), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n544), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT88), .B(new_n553), .C1(new_n554), .C2(new_n501), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n499), .B(new_n510), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G197gat), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT11), .B(G169gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT12), .Z(new_n564));
  INV_X1    g363(.A(G29gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT14), .B(G29gat), .Z(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(G36gat), .ZN(new_n568));
  AND2_X1   g367(.A1(G43gat), .A2(G50gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(G43gat), .A2(G50gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT15), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT94), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT93), .B(G43gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(G50gat), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n568), .A2(new_n576), .A3(new_n571), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT16), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(G1gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(G1gat), .B2(new_n582), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(G8gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n578), .A2(new_n586), .A3(new_n580), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(KEYINPUT95), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT13), .Z(new_n592));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n593), .A3(new_n586), .A4(new_n580), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT96), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n590), .A2(new_n597), .A3(new_n592), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n578), .A2(KEYINPUT17), .A3(new_n580), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n586), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n604), .A2(new_n588), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(KEYINPUT18), .A3(new_n591), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n591), .A3(new_n588), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n564), .B1(new_n600), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n564), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n599), .A2(new_n612), .A3(new_n609), .A4(new_n606), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(KEYINPUT97), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n615), .B(new_n564), .C1(new_n600), .C2(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n559), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G230gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n346), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT8), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(KEYINPUT101), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(KEYINPUT101), .B2(new_n623), .ZN(new_n625));
  NAND2_X1  g424(.A1(G85gat), .A2(G92gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT7), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT102), .B(G85gat), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n625), .B(new_n627), .C1(G92gat), .C2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT107), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G99gat), .B(G106gat), .Z(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G64gat), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(G57gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(G57gat), .ZN(new_n636));
  AND2_X1   g435(.A1(G71gat), .A2(G78gat), .ZN(new_n637));
  OAI22_X1  g436(.A1(new_n635), .A2(new_n636), .B1(KEYINPUT9), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G71gat), .B(G78gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n629), .B1(KEYINPUT103), .B2(new_n632), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n632), .A2(KEYINPUT103), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n640), .B(KEYINPUT98), .Z(new_n647));
  OAI211_X1 g446(.A(new_n642), .B(new_n643), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT10), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n621), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n651), .A2(new_n621), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT108), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n657), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n647), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT21), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G231gat), .A2(G233gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G127gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G183gat), .B(G211gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n587), .B1(new_n647), .B2(KEYINPUT21), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G155gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n671), .B(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n669), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n646), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n602), .A2(new_n603), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(G232gat), .A2(G233gat), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n581), .A2(new_n646), .B1(KEYINPUT41), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(G190gat), .B(G218gat), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n682), .A2(KEYINPUT105), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT105), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n680), .A2(KEYINPUT41), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT100), .ZN(new_n687));
  XOR2_X1   g486(.A(G134gat), .B(G162gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OAI22_X1  g488(.A1(new_n684), .A2(new_n685), .B1(KEYINPUT106), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n683), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n679), .A2(new_n691), .A3(new_n681), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT104), .Z(new_n693));
  INV_X1    g492(.A(new_n689), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n690), .B2(new_n693), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AND4_X1   g499(.A1(new_n619), .A2(new_n661), .A3(new_n677), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n496), .B(KEYINPUT109), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  INV_X1    g504(.A(new_n322), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n707), .A2(G8gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT16), .B(G8gat), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT42), .B2(new_n710), .ZN(G1325gat));
  INV_X1    g511(.A(G15gat), .ZN(new_n713));
  INV_X1    g512(.A(new_n372), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n701), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n701), .A2(new_n553), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n713), .ZN(G1326gat));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n554), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(new_n677), .ZN(new_n721));
  AND4_X1   g520(.A1(new_n619), .A2(new_n661), .A3(new_n721), .A4(new_n699), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n565), .A3(new_n703), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n544), .A2(new_n555), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n510), .A2(new_n499), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n699), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n559), .A2(KEYINPUT44), .A3(new_n699), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n660), .B(KEYINPUT110), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n721), .A2(new_n618), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT111), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(new_n703), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n724), .B1(new_n739), .B2(new_n565), .ZN(G1328gat));
  INV_X1    g539(.A(G36gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n722), .A2(new_n741), .A3(new_n706), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT46), .Z(new_n743));
  AND2_X1   g542(.A1(new_n738), .A2(new_n706), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n741), .ZN(G1329gat));
  INV_X1    g544(.A(new_n553), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n575), .B1(new_n734), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n372), .A2(new_n575), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n722), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(KEYINPUT47), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n553), .A3(new_n737), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n751), .A2(new_n575), .B1(new_n722), .B2(new_n748), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g552(.A(KEYINPUT48), .B(G50gat), .C1(new_n734), .C2(new_n530), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n530), .A2(G50gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT112), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n722), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n754), .B(new_n757), .C1(new_n758), .C2(KEYINPUT48), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n735), .A2(new_n554), .A3(new_n737), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n677), .A2(new_n700), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n764), .A2(new_n618), .A3(new_n732), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(new_n726), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n703), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT114), .B(G57gat), .Z(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1332gat));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n706), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT49), .B(G64gat), .Z(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(G71gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n766), .A2(new_n774), .A3(new_n714), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n766), .A2(new_n553), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(new_n774), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g577(.A1(new_n766), .A2(new_n554), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g579(.A1(new_n721), .A2(new_n617), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n661), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n729), .A2(new_n730), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT115), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n729), .A2(new_n730), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n628), .B1(new_n787), .B2(new_n702), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n727), .A2(new_n781), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  OR3_X1    g589(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n781), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OR3_X1    g591(.A1(new_n702), .A2(new_n661), .A3(new_n628), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n788), .B1(new_n792), .B2(new_n793), .ZN(G1336gat));
  OAI21_X1  g593(.A(G92gat), .B1(new_n783), .B2(new_n322), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n732), .A2(G92gat), .A3(new_n322), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n795), .B(new_n796), .C1(new_n792), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n789), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n798), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n706), .A3(new_n786), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(G92gat), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n799), .B1(new_n805), .B2(new_n796), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n787), .B2(new_n746), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n661), .A2(G99gat), .A3(new_n372), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n792), .B2(new_n808), .ZN(G1338gat));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n783), .B2(new_n530), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n732), .A2(G106gat), .A3(new_n530), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n810), .B(new_n811), .C1(new_n792), .C2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n784), .A2(new_n554), .A3(new_n786), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n817), .A2(new_n818), .A3(G106gat), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n817), .B2(G106gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n802), .A2(new_n813), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n816), .B1(new_n822), .B2(new_n810), .ZN(G1339gat));
  INV_X1    g622(.A(new_n650), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n648), .A2(new_n621), .A3(new_n649), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n656), .B1(new_n650), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT55), .B1(new_n826), .B2(new_n828), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n650), .A2(new_n652), .A3(new_n657), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n614), .A2(new_n832), .A3(new_n616), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n605), .A2(new_n591), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n592), .B1(new_n590), .B2(new_n594), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n563), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n660), .A2(new_n613), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n699), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n613), .A2(new_n836), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT119), .Z(new_n840));
  NAND3_X1  g639(.A1(new_n697), .A2(new_n832), .A3(new_n698), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n721), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n677), .A2(new_n617), .A3(new_n661), .A4(new_n700), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(KEYINPUT120), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n706), .A2(new_n702), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n849), .A2(new_n508), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n618), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g653(.A(G120gat), .B1(new_n852), .B2(new_n660), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n732), .A2(new_n330), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n852), .B2(new_n856), .ZN(G1341gat));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n677), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(G127gat), .ZN(G1342gat));
  AND2_X1   g658(.A1(new_n852), .A2(new_n699), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n843), .A2(KEYINPUT120), .A3(new_n844), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT120), .B1(new_n843), .B2(new_n844), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n699), .A2(new_n322), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(G134gat), .A3(new_n702), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n456), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n860), .A2(new_n323), .B1(new_n868), .B2(new_n869), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n553), .A2(new_n530), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n861), .A2(new_n862), .A3(new_n702), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT122), .B1(new_n849), .B2(new_n702), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n617), .A2(G141gat), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT123), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n875), .A2(new_n322), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n847), .A2(new_n880), .A3(new_n554), .A4(new_n848), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n833), .A2(new_n837), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT121), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n700), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n842), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n677), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n844), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n554), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT57), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n851), .A2(new_n553), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n881), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n617), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT58), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT57), .B1(new_n849), .B2(new_n530), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n844), .B(KEYINPUT124), .Z(new_n902));
  OAI211_X1 g701(.A(new_n880), .B(new_n554), .C1(new_n902), .C2(new_n888), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n901), .A2(new_n660), .A3(new_n903), .A4(new_n892), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n900), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n893), .A2(new_n661), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n900), .A2(G148gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n875), .A2(new_n322), .A3(new_n876), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n661), .A2(G148gat), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n905), .A2(new_n908), .B1(new_n909), .B2(new_n910), .ZN(G1345gat));
  NOR2_X1   g710(.A1(new_n721), .A2(G155gat), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n875), .A2(new_n322), .A3(new_n876), .A4(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G155gat), .B1(new_n893), .B2(new_n721), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT125), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n893), .B2(new_n700), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n864), .A2(G162gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n875), .A2(new_n876), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n703), .A2(new_n322), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n508), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n863), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n617), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(G169gat), .Z(G1348gat));
  OAI21_X1  g728(.A(G176gat), .B1(new_n927), .B2(new_n732), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n661), .A2(G176gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n927), .B2(new_n931), .ZN(G1349gat));
  OR3_X1    g731(.A1(new_n927), .A2(new_n251), .A3(new_n721), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n218), .B1(new_n927), .B2(new_n721), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1350gat));
  OAI22_X1  g737(.A1(new_n927), .A2(new_n700), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n553), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n901), .A2(new_n903), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(G197gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n617), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n863), .A2(new_n554), .A3(new_n942), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(new_n617), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(G1352gat));
  OAI21_X1  g748(.A(G204gat), .B1(new_n944), .B2(new_n732), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n661), .A2(G204gat), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n947), .A2(KEYINPUT62), .A3(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(G1353gat));
  NAND4_X1  g754(.A1(new_n901), .A2(new_n677), .A3(new_n903), .A4(new_n942), .ZN(new_n956));
  AND2_X1   g755(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n957));
  OAI21_X1  g756(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n957), .B1(new_n956), .B2(new_n959), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n677), .A2(new_n205), .ZN(new_n962));
  OAI22_X1  g761(.A1(new_n960), .A2(new_n961), .B1(new_n947), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(new_n699), .B1(new_n441), .B2(new_n440), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n944), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n947), .A2(new_n700), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n966), .A2(G218gat), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n965), .A2(new_n967), .ZN(G1355gat));
endmodule


