

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(G651), .A2(n635), .ZN(n648) );
  XNOR2_X1 U553 ( .A(n721), .B(n720), .ZN(n726) );
  XNOR2_X1 U554 ( .A(n761), .B(KEYINPUT97), .ZN(n762) );
  NAND2_X1 U555 ( .A1(n813), .A2(n812), .ZN(n815) );
  XNOR2_X1 U556 ( .A(n522), .B(KEYINPUT23), .ZN(n523) );
  AND2_X1 U557 ( .A1(G2104), .A2(G101), .ZN(n521) );
  NOR2_X2 U558 ( .A1(G543), .A2(G651), .ZN(n580) );
  OR2_X1 U559 ( .A1(KEYINPUT33), .A2(n765), .ZN(n518) );
  OR2_X1 U560 ( .A1(n799), .A2(n738), .ZN(n519) );
  NOR2_X1 U561 ( .A1(n699), .A2(n698), .ZN(n700) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n720) );
  NOR2_X1 U563 ( .A1(n732), .A2(n731), .ZN(n733) );
  INV_X1 U564 ( .A(KEYINPUT95), .ZN(n736) );
  NOR2_X1 U565 ( .A1(G1966), .A2(n738), .ZN(n750) );
  INV_X1 U566 ( .A(KEYINPUT64), .ZN(n763) );
  XNOR2_X1 U567 ( .A(n764), .B(n763), .ZN(n765) );
  AND2_X1 U568 ( .A1(n800), .A2(n519), .ZN(n801) );
  INV_X1 U569 ( .A(KEYINPUT99), .ZN(n814) );
  INV_X1 U570 ( .A(KEYINPUT66), .ZN(n522) );
  XNOR2_X1 U571 ( .A(n815), .B(n814), .ZN(n817) );
  NAND2_X1 U572 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U573 ( .A1(n530), .A2(n529), .ZN(G160) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n520), .Z(n686) );
  NAND2_X1 U576 ( .A1(G137), .A2(n686), .ZN(n526) );
  INV_X1 U577 ( .A(G2105), .ZN(n543) );
  NAND2_X1 U578 ( .A1(n543), .A2(n521), .ZN(n524) );
  XNOR2_X1 U579 ( .A(n524), .B(n523), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n526), .A2(n525), .ZN(n530) );
  NOR2_X2 U581 ( .A1(G2104), .A2(n543), .ZN(n889) );
  NAND2_X1 U582 ( .A1(G125), .A2(n889), .ZN(n528) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U584 ( .A1(G113), .A2(n890), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U586 ( .A(G2427), .B(KEYINPUT102), .ZN(n540) );
  XOR2_X1 U587 ( .A(G2430), .B(G2446), .Z(n532) );
  XNOR2_X1 U588 ( .A(KEYINPUT103), .B(G2438), .ZN(n531) );
  XNOR2_X1 U589 ( .A(n532), .B(n531), .ZN(n536) );
  XOR2_X1 U590 ( .A(G2435), .B(G2454), .Z(n534) );
  XNOR2_X1 U591 ( .A(G1348), .B(G1341), .ZN(n533) );
  XNOR2_X1 U592 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U593 ( .A(n536), .B(n535), .Z(n538) );
  XNOR2_X1 U594 ( .A(G2451), .B(G2443), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n540), .B(n539), .ZN(n541) );
  AND2_X1 U597 ( .A1(n541), .A2(G14), .ZN(G401) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U599 ( .A1(G123), .A2(n889), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n542), .B(KEYINPUT18), .ZN(n551) );
  AND2_X1 U601 ( .A1(n543), .A2(G2104), .ZN(n885) );
  NAND2_X1 U602 ( .A1(G99), .A2(n885), .ZN(n546) );
  INV_X1 U603 ( .A(n686), .ZN(n544) );
  INV_X1 U604 ( .A(n544), .ZN(n886) );
  NAND2_X1 U605 ( .A1(G135), .A2(n886), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G111), .A2(n890), .ZN(n547) );
  XNOR2_X1 U608 ( .A(KEYINPUT79), .B(n547), .ZN(n548) );
  NOR2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U610 ( .A1(n551), .A2(n550), .ZN(n922) );
  XNOR2_X1 U611 ( .A(G2096), .B(n922), .ZN(n552) );
  OR2_X1 U612 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  XOR2_X1 U614 ( .A(G543), .B(KEYINPUT0), .Z(n635) );
  NAND2_X1 U615 ( .A1(G52), .A2(n648), .ZN(n556) );
  INV_X1 U616 ( .A(G651), .ZN(n557) );
  NOR2_X1 U617 ( .A1(G543), .A2(n557), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n553) );
  XNOR2_X2 U619 ( .A(n554), .B(n553), .ZN(n651) );
  NAND2_X1 U620 ( .A1(G64), .A2(n651), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G90), .A2(n580), .ZN(n559) );
  NOR2_X2 U623 ( .A1(n635), .A2(n557), .ZN(n646) );
  NAND2_X1 U624 ( .A1(G77), .A2(n646), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U628 ( .A1(n580), .A2(G89), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT4), .B(n563), .Z(n566) );
  NAND2_X1 U630 ( .A1(n646), .A2(G76), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT74), .B(n564), .Z(n565) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT75), .B(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT5), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G51), .A2(n648), .ZN(n570) );
  NAND2_X1 U636 ( .A1(G63), .A2(n651), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT76), .B(KEYINPUT6), .Z(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT7), .B(n575), .ZN(G168) );
  XOR2_X1 U642 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n577) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n835) );
  NAND2_X1 U646 ( .A1(n835), .A2(G567), .ZN(n578) );
  XOR2_X1 U647 ( .A(KEYINPUT11), .B(n578), .Z(G234) );
  NAND2_X1 U648 ( .A1(n651), .A2(G56), .ZN(n579) );
  XNOR2_X1 U649 ( .A(n579), .B(KEYINPUT14), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G81), .A2(n580), .ZN(n581) );
  XNOR2_X1 U651 ( .A(n581), .B(KEYINPUT12), .ZN(n582) );
  XNOR2_X1 U652 ( .A(n582), .B(KEYINPUT72), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G68), .A2(n646), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U655 ( .A(n585), .B(KEYINPUT13), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT73), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G43), .A2(n648), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n982) );
  INV_X1 U659 ( .A(G860), .ZN(n609) );
  OR2_X1 U660 ( .A1(n982), .A2(n609), .ZN(G153) );
  INV_X1 U661 ( .A(G171), .ZN(G301) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G92), .A2(n580), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G66), .A2(n651), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G79), .A2(n646), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G54), .A2(n648), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n597), .Z(n977) );
  INV_X1 U671 ( .A(n977), .ZN(n706) );
  INV_X1 U672 ( .A(G868), .ZN(n666) );
  NAND2_X1 U673 ( .A1(n706), .A2(n666), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(G284) );
  XOR2_X1 U675 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U676 ( .A1(G91), .A2(n580), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G78), .A2(n646), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n648), .A2(G53), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT70), .B(n602), .Z(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n651), .A2(G65), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n606), .A2(n605), .ZN(G299) );
  NOR2_X1 U684 ( .A1(G286), .A2(n666), .ZN(n608) );
  NOR2_X1 U685 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n610), .A2(n977), .ZN(n611) );
  XNOR2_X1 U689 ( .A(n611), .B(KEYINPUT16), .ZN(n612) );
  XOR2_X1 U690 ( .A(KEYINPUT77), .B(n612), .Z(G148) );
  NOR2_X1 U691 ( .A1(n706), .A2(n666), .ZN(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT78), .B(n613), .Z(n614) );
  NOR2_X1 U693 ( .A1(G559), .A2(n614), .ZN(n616) );
  NOR2_X1 U694 ( .A1(G868), .A2(n982), .ZN(n615) );
  NOR2_X1 U695 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U696 ( .A1(n977), .A2(G559), .ZN(n664) );
  XNOR2_X1 U697 ( .A(n982), .B(n664), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n617), .A2(G860), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G93), .A2(n580), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G80), .A2(n646), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G67), .A2(n651), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT80), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n648), .A2(G55), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  OR2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n667) );
  XOR2_X1 U707 ( .A(n625), .B(n667), .Z(G145) );
  NAND2_X1 U708 ( .A1(G88), .A2(n580), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G75), .A2(n646), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G50), .A2(n648), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G62), .A2(n651), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G49), .A2(n648), .ZN(n633) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U718 ( .A1(n651), .A2(n634), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U721 ( .A1(n651), .A2(G60), .ZN(n638) );
  XNOR2_X1 U722 ( .A(n638), .B(KEYINPUT68), .ZN(n645) );
  NAND2_X1 U723 ( .A1(G85), .A2(n580), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G72), .A2(n646), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U726 ( .A1(G47), .A2(n648), .ZN(n641) );
  XNOR2_X1 U727 ( .A(KEYINPUT69), .B(n641), .ZN(n642) );
  NOR2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U730 ( .A1(G73), .A2(n646), .ZN(n647) );
  XNOR2_X1 U731 ( .A(n647), .B(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U732 ( .A1(G86), .A2(n580), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G48), .A2(n648), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U735 ( .A1(G61), .A2(n651), .ZN(n652) );
  XNOR2_X1 U736 ( .A(KEYINPUT81), .B(n652), .ZN(n653) );
  NOR2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(G305) );
  XOR2_X1 U739 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n657) );
  XNOR2_X1 U740 ( .A(G288), .B(n657), .ZN(n658) );
  XNOR2_X1 U741 ( .A(G166), .B(n658), .ZN(n660) );
  INV_X1 U742 ( .A(G299), .ZN(n714) );
  XNOR2_X1 U743 ( .A(G290), .B(n714), .ZN(n659) );
  XNOR2_X1 U744 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U745 ( .A(n667), .B(n661), .Z(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(G305), .ZN(n663) );
  XNOR2_X1 U747 ( .A(n982), .B(n663), .ZN(n907) );
  XOR2_X1 U748 ( .A(n907), .B(n664), .Z(n665) );
  NOR2_X1 U749 ( .A1(n666), .A2(n665), .ZN(n669) );
  NOR2_X1 U750 ( .A1(G868), .A2(n667), .ZN(n668) );
  NOR2_X1 U751 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n671), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n672) );
  XNOR2_X1 U756 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G2072), .ZN(n675) );
  XNOR2_X1 U758 ( .A(n675), .B(KEYINPUT84), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n677) );
  NAND2_X1 U761 ( .A1(G132), .A2(G82), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U763 ( .A1(n678), .A2(G218), .ZN(n679) );
  NAND2_X1 U764 ( .A1(G96), .A2(n679), .ZN(n839) );
  NAND2_X1 U765 ( .A1(n839), .A2(G2106), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U767 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U768 ( .A1(G108), .A2(n681), .ZN(n840) );
  NAND2_X1 U769 ( .A1(n840), .A2(G567), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n841) );
  NAND2_X1 U771 ( .A1(G661), .A2(G483), .ZN(n684) );
  XNOR2_X1 U772 ( .A(KEYINPUT86), .B(n684), .ZN(n685) );
  NOR2_X1 U773 ( .A1(n841), .A2(n685), .ZN(n838) );
  NAND2_X1 U774 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U775 ( .A1(G102), .A2(n885), .ZN(n688) );
  NAND2_X1 U776 ( .A1(G138), .A2(n686), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U778 ( .A1(G126), .A2(n889), .ZN(n690) );
  NAND2_X1 U779 ( .A1(G114), .A2(n890), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U781 ( .A1(n692), .A2(n691), .ZN(G164) );
  INV_X1 U782 ( .A(G166), .ZN(G303) );
  NOR2_X1 U783 ( .A1(G164), .A2(G1384), .ZN(n768) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n767) );
  INV_X1 U785 ( .A(KEYINPUT92), .ZN(n693) );
  XNOR2_X1 U786 ( .A(n767), .B(n693), .ZN(n694) );
  NAND2_X2 U787 ( .A1(n768), .A2(n694), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(G1341), .ZN(n696) );
  INV_X1 U789 ( .A(n982), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n699) );
  INV_X1 U791 ( .A(G1996), .ZN(n944) );
  NOR2_X1 U792 ( .A1(n740), .A2(n944), .ZN(n697) );
  XNOR2_X1 U793 ( .A(n697), .B(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U794 ( .A(n700), .B(KEYINPUT65), .ZN(n704) );
  INV_X1 U795 ( .A(n740), .ZN(n722) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n722), .ZN(n702) );
  NAND2_X1 U797 ( .A1(G1348), .A2(n740), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n705) );
  OR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n722), .A2(G2072), .ZN(n709) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT27), .ZN(n711) );
  AND2_X1 U805 ( .A1(G1956), .A2(n740), .ZN(n710) );
  NOR2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n719) );
  NOR2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n717) );
  INV_X1 U810 ( .A(KEYINPUT28), .ZN(n716) );
  XNOR2_X1 U811 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U813 ( .A(KEYINPUT93), .B(G1961), .ZN(n993) );
  NAND2_X1 U814 ( .A1(n740), .A2(n993), .ZN(n724) );
  XNOR2_X1 U815 ( .A(G2078), .B(KEYINPUT25), .ZN(n949) );
  NAND2_X1 U816 ( .A1(n722), .A2(n949), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n730) );
  NAND2_X1 U818 ( .A1(n730), .A2(G171), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n735) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n740), .ZN(n752) );
  NAND2_X1 U821 ( .A1(G8), .A2(n740), .ZN(n738) );
  NOR2_X1 U822 ( .A1(n752), .A2(n750), .ZN(n727) );
  NAND2_X1 U823 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U824 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U825 ( .A1(n729), .A2(G168), .ZN(n732) );
  NOR2_X1 U826 ( .A1(G171), .A2(n730), .ZN(n731) );
  XOR2_X1 U827 ( .A(KEYINPUT31), .B(n733), .Z(n734) );
  NAND2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n748) );
  NAND2_X1 U829 ( .A1(G286), .A2(n748), .ZN(n737) );
  XNOR2_X1 U830 ( .A(n737), .B(n736), .ZN(n745) );
  INV_X1 U831 ( .A(n738), .ZN(n739) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n738), .ZN(n742) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U835 ( .A1(G303), .A2(n743), .ZN(n744) );
  NAND2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n746), .A2(G8), .ZN(n747) );
  XNOR2_X1 U838 ( .A(n747), .B(KEYINPUT32), .ZN(n756) );
  INV_X1 U839 ( .A(n748), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U841 ( .A(n751), .B(KEYINPUT94), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n752), .A2(G8), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n802) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n757) );
  XNOR2_X1 U847 ( .A(KEYINPUT96), .B(n757), .ZN(n758) );
  NOR2_X1 U848 ( .A1(n976), .A2(n758), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n802), .A2(n759), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NAND2_X1 U851 ( .A1(n760), .A2(n973), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n739), .ZN(n764) );
  XOR2_X1 U853 ( .A(G1981), .B(KEYINPUT98), .Z(n766) );
  XNOR2_X1 U854 ( .A(G305), .B(n766), .ZN(n967) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n829) );
  XNOR2_X1 U856 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  NAND2_X1 U857 ( .A1(G104), .A2(n885), .ZN(n770) );
  NAND2_X1 U858 ( .A1(G140), .A2(n886), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n771), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n890), .A2(G116), .ZN(n772) );
  XOR2_X1 U862 ( .A(KEYINPUT87), .B(n772), .Z(n774) );
  NAND2_X1 U863 ( .A1(n889), .A2(G128), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  NOR2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n778), .ZN(n896) );
  NOR2_X1 U868 ( .A1(n827), .A2(n896), .ZN(n937) );
  NAND2_X1 U869 ( .A1(n829), .A2(n937), .ZN(n779) );
  XNOR2_X1 U870 ( .A(KEYINPUT88), .B(n779), .ZN(n825) );
  AND2_X1 U871 ( .A1(n967), .A2(n825), .ZN(n798) );
  NAND2_X1 U872 ( .A1(G95), .A2(n885), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G131), .A2(n886), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G119), .A2(n889), .ZN(n782) );
  XNOR2_X1 U876 ( .A(KEYINPUT89), .B(n782), .ZN(n783) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n890), .A2(G107), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n899) );
  XNOR2_X1 U880 ( .A(KEYINPUT90), .B(G1991), .ZN(n955) );
  NAND2_X1 U881 ( .A1(n899), .A2(n955), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G141), .A2(n886), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G129), .A2(n889), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n885), .A2(G105), .ZN(n789) );
  XOR2_X1 U886 ( .A(KEYINPUT38), .B(n789), .Z(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n890), .A2(G117), .ZN(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n900) );
  NAND2_X1 U890 ( .A1(G1996), .A2(n900), .ZN(n794) );
  NAND2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U892 ( .A(KEYINPUT91), .B(n796), .ZN(n927) );
  INV_X1 U893 ( .A(n927), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n797), .A2(n829), .ZN(n818) );
  AND2_X1 U895 ( .A1(n798), .A2(n818), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n976), .A2(KEYINPUT33), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n518), .A2(n801), .ZN(n813) );
  NOR2_X1 U898 ( .A1(G2090), .A2(G303), .ZN(n803) );
  NAND2_X1 U899 ( .A1(G8), .A2(n803), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n802), .A2(n804), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n805), .A2(n738), .ZN(n809) );
  NOR2_X1 U902 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XOR2_X1 U903 ( .A(n806), .B(KEYINPUT24), .Z(n807) );
  OR2_X1 U904 ( .A1(n738), .A2(n807), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  AND2_X1 U906 ( .A1(n825), .A2(n810), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n818), .A2(n811), .ZN(n812) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U909 ( .A1(n979), .A2(n829), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n832) );
  XNOR2_X1 U911 ( .A(KEYINPUT39), .B(KEYINPUT100), .ZN(n824) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n900), .ZN(n929) );
  INV_X1 U913 ( .A(n818), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n955), .A2(n899), .ZN(n925) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n925), .A2(n819), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n929), .A2(n822), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n824), .B(n823), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n827), .A2(n896), .ZN(n934) );
  NAND2_X1 U922 ( .A1(n828), .A2(n934), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n834) );
  XOR2_X1 U925 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n833) );
  XNOR2_X1 U926 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U929 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U933 ( .A(G132), .ZN(G219) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G82), .ZN(G220) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n841), .ZN(G319) );
  XOR2_X1 U941 ( .A(G2100), .B(G2096), .Z(n843) );
  XNOR2_X1 U942 ( .A(KEYINPUT42), .B(G2678), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2090), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2084), .B(G2078), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1961), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n864) );
  XOR2_X1 U953 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n853) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n854), .B(KEYINPUT104), .Z(n862) );
  XOR2_X1 U957 ( .A(KEYINPUT105), .B(G1981), .Z(n856) );
  XNOR2_X1 U958 ( .A(G1966), .B(G1956), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U960 ( .A(G2474), .B(KEYINPUT109), .Z(n858) );
  XNOR2_X1 U961 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(n864), .B(n863), .Z(G229) );
  NAND2_X1 U966 ( .A1(G100), .A2(n885), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G112), .A2(n890), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G124), .A2(n889), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G136), .A2(n886), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n868), .B(KEYINPUT110), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G130), .A2(n889), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G118), .A2(n890), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G106), .A2(n885), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G142), .A2(n886), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n877), .ZN(n878) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n878), .ZN(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(n881), .B(KEYINPUT46), .Z(n883) );
  XNOR2_X1 U985 ( .A(G164), .B(KEYINPUT48), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U987 ( .A(G162), .B(n884), .ZN(n898) );
  NAND2_X1 U988 ( .A1(G103), .A2(n885), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G139), .A2(n886), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G127), .A2(n889), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G115), .A2(n890), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n917) );
  XNOR2_X1 U996 ( .A(n896), .B(n917), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n904) );
  XOR2_X1 U998 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U999 ( .A(n922), .B(n901), .ZN(n902) );
  XOR2_X1 U1000 ( .A(G160), .B(n902), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(G171), .B(n977), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n906), .B(G286), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G397) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT113), .B(n914), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1017 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(G2072), .B(n917), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(G164), .B(G2078), .ZN(n918) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n940) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT114), .B(n930), .Z(n931) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n931), .Z(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(n938), .B(KEYINPUT115), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n1021), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n960) );
  XNOR2_X1 U1040 ( .A(G32), .B(n944), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G27), .B(n949), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(KEYINPUT117), .B(n950), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(KEYINPUT118), .B(n953), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n954), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G25), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n1022) );
  NOR2_X1 U1057 ( .A1(G29), .A2(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n1022), .A2(n964), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n965), .ZN(n1028) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XOR2_X1 U1061 ( .A(G1966), .B(G168), .Z(n966) );
  XNOR2_X1 U1062 ( .A(KEYINPUT119), .B(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(n970), .B(n969), .ZN(n989) );
  XNOR2_X1 U1066 ( .A(G301), .B(G1961), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G299), .B(G1956), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n986) );
  XNOR2_X1 U1071 ( .A(n977), .B(G1348), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G1971), .B(G303), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(KEYINPUT122), .ZN(n1026) );
  XNOR2_X1 U1082 ( .A(G5), .B(n993), .ZN(n1010) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G21), .ZN(n1008) );
  INV_X1 U1084 ( .A(G1956), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n994), .B(G20), .ZN(n1004) );
  XOR2_X1 U1086 ( .A(G1341), .B(G19), .Z(n999) );
  XOR2_X1 U1087 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT59), .B(G4), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n996), .B(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n997), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(KEYINPUT123), .B(G1981), .Z(n1000) );
  XNOR2_X1 U1093 ( .A(G6), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT60), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1103 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(n1018), .B(KEYINPUT61), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT127), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(G16), .A2(n1020), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

