//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(new_n190), .A3(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT67), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT11), .B1(new_n204), .B2(G134), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G134), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n203), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(G131), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n202), .B1(new_n209), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT64), .B(G143), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G146), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n221), .B2(G146), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n222), .A2(new_n225), .B1(new_n228), .B2(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(G131), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT65), .A2(G131), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT65), .A2(G131), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n208), .A3(new_n212), .A4(new_n213), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n234), .A3(KEYINPUT68), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n217), .A2(new_n229), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n237));
  OAI21_X1  g051(.A(G128), .B1(new_n227), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  AOI21_X1  g055(.A(G146), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n238), .B1(new_n242), .B2(new_n219), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n241), .A3(G146), .ZN(new_n244));
  INV_X1    g058(.A(new_n227), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n237), .A3(G128), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n204), .A3(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT66), .B1(new_n211), .B2(G137), .ZN(new_n250));
  OAI211_X1 g064(.A(G131), .B(new_n249), .C1(new_n250), .C2(new_n206), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n247), .A2(new_n234), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n236), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n201), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n234), .A2(new_n251), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n243), .B2(new_n246), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n230), .A2(new_n234), .A3(KEYINPUT68), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT68), .B1(new_n230), .B2(new_n234), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n257), .B1(new_n260), .B2(new_n229), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT28), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n200), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n230), .A2(new_n234), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n225), .B1(new_n242), .B2(new_n219), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n244), .A2(new_n223), .A3(new_n245), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n201), .B1(new_n271), .B2(new_n257), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n265), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  XOR2_X1   g088(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n275), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n264), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n236), .A2(KEYINPUT30), .A3(new_n252), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n271), .B2(new_n257), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n287), .A3(new_n201), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n266), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n281), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n253), .A2(new_n201), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n265), .B1(new_n266), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n281), .A2(new_n284), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n264), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n264), .A2(new_n294), .A3(KEYINPUT72), .A4(new_n295), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G902), .Z(new_n300));
  NAND4_X1  g114(.A1(new_n291), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G472), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n281), .B1(new_n263), .B2(new_n273), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT31), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n266), .A3(new_n282), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n288), .A2(new_n266), .A3(KEYINPUT70), .A4(new_n282), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n305), .A2(new_n304), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  NOR2_X1   g126(.A1(G472), .A2(G902), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n311), .B2(new_n313), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n302), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT9), .B(G234), .ZN(new_n317));
  OAI21_X1  g131(.A(G221), .B1(new_n317), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT80), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n277), .A2(G227), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G107), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G104), .ZN(new_n327));
  INV_X1    g141(.A(G104), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G107), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G101), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT3), .B1(new_n328), .B2(G107), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n326), .A3(G104), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n334), .A3(new_n329), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT83), .B(G101), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n339), .A2(G128), .B1(new_n245), .B2(new_n244), .ZN(new_n340));
  INV_X1    g154(.A(new_n246), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n243), .B2(new_n246), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n342), .A2(new_n343), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n346));
  INV_X1    g160(.A(new_n335), .ZN(new_n347));
  INV_X1    g161(.A(new_n336), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n335), .A2(G101), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n335), .A2(KEYINPUT82), .A3(G101), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT84), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n335), .A2(new_n346), .A3(G101), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n268), .A2(new_n356), .A3(new_n269), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n335), .A2(KEYINPUT82), .A3(G101), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT4), .B1(new_n335), .B2(new_n336), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT82), .B1(new_n335), .B2(G101), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n268), .A2(new_n356), .A3(new_n269), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT84), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n345), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n260), .ZN(new_n366));
  INV_X1    g180(.A(new_n260), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n345), .A2(new_n367), .A3(new_n364), .A4(new_n358), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n325), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n267), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n244), .A2(new_n245), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n239), .A2(new_n241), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n237), .B1(new_n372), .B2(new_n218), .ZN(new_n373));
  INV_X1    g187(.A(G128), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n337), .B1(new_n375), .B2(new_n246), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n337), .A2(new_n243), .A3(new_n246), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n370), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n337), .A2(new_n243), .A3(new_n246), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n342), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT12), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n378), .A2(KEYINPUT12), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT81), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n369), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n325), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n320), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n300), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n366), .A2(new_n368), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n368), .A2(new_n382), .A3(new_n324), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n391), .A2(new_n325), .B1(new_n392), .B2(KEYINPUT85), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n368), .A2(new_n382), .A3(new_n394), .A4(new_n324), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n390), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n389), .B1(new_n396), .B2(new_n320), .ZN(new_n397));
  NAND2_X1  g211(.A1(G469), .A2(G902), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n319), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT93), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n401));
  XOR2_X1   g215(.A(G113), .B(G122), .Z(new_n402));
  XOR2_X1   g216(.A(KEYINPUT90), .B(G104), .Z(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT90), .B(G104), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n276), .A2(new_n277), .A3(G143), .A4(G214), .ZN(new_n409));
  INV_X1    g223(.A(G214), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n410), .A2(G237), .A3(G953), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n233), .B(new_n409), .C1(new_n372), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT89), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n276), .A2(new_n277), .A3(G214), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n239), .A3(new_n241), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n409), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n215), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n415), .A2(new_n418), .A3(new_n233), .A4(new_n409), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G125), .ZN(new_n422));
  INV_X1    g236(.A(G125), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G140), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n424), .A3(KEYINPUT76), .ZN(new_n425));
  OR3_X1    g239(.A1(new_n423), .A2(KEYINPUT76), .A3(G140), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT16), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n423), .A2(G140), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n428), .A2(KEYINPUT16), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G146), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT19), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n421), .A2(G125), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n422), .A2(new_n424), .A3(KEYINPUT77), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n437), .B2(KEYINPUT19), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n420), .B(new_n431), .C1(G146), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n218), .A3(new_n436), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n425), .A2(new_n426), .A3(G146), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT18), .A2(G131), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n415), .A2(new_n409), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n416), .A2(KEYINPUT18), .A3(G131), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n408), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n408), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n413), .A2(new_n417), .A3(new_n450), .A4(new_n419), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n427), .A2(new_n218), .A3(new_n429), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n215), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n431), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n449), .B(new_n446), .C1(new_n452), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n451), .A2(new_n453), .A3(new_n431), .A4(new_n454), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(KEYINPUT92), .A3(new_n446), .A4(new_n449), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n447), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(G475), .A2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n400), .B(new_n401), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n427), .A2(new_n218), .A3(new_n429), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n218), .B1(new_n427), .B2(new_n429), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n450), .B(new_n233), .C1(new_n415), .C2(new_n409), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n465), .B1(new_n469), .B2(new_n451), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n408), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n458), .A2(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G475), .B1(new_n473), .B2(G902), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n277), .A2(G952), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(G234), .B2(G237), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n277), .B(new_n300), .C1(G234), .C2(G237), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n239), .A2(new_n241), .A3(G128), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n374), .A2(G143), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n211), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n193), .A2(G122), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n193), .A2(G122), .ZN(new_n486));
  OAI21_X1  g300(.A(G107), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G116), .B(G122), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n326), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT13), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT94), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT94), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT13), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n482), .A2(new_n483), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G134), .B1(new_n482), .B2(new_n495), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n484), .B(new_n490), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT95), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n482), .A2(new_n483), .A3(new_n495), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(G134), .C1(new_n482), .C2(new_n495), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(KEYINPUT95), .A3(new_n484), .A4(new_n490), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n482), .A2(new_n483), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G134), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n484), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n326), .B1(new_n485), .B2(KEYINPUT14), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n488), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n507), .A2(new_n509), .B1(new_n326), .B2(new_n488), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G217), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n317), .A2(new_n512), .A3(G953), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n500), .A2(new_n503), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n498), .A2(new_n499), .B1(new_n506), .B2(new_n510), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n513), .B1(new_n516), .B2(new_n503), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n300), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G478), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n518), .B(new_n520), .Z(new_n521));
  INV_X1    g335(.A(new_n447), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT92), .B1(new_n470), .B2(new_n449), .ZN(new_n523));
  INV_X1    g337(.A(new_n460), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT93), .A3(new_n462), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n400), .B1(new_n461), .B2(new_n463), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT20), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n475), .A2(new_n481), .A3(new_n521), .A4(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G210), .B1(G237), .B2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT5), .ZN(new_n532));
  OAI21_X1  g346(.A(G113), .B1(new_n192), .B2(KEYINPUT5), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n195), .A2(new_n196), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n338), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n198), .A2(new_n199), .A3(new_n356), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n362), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G122), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n537), .B(new_n540), .C1(new_n362), .C2(new_n538), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT6), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G224), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n270), .A2(new_n423), .ZN(new_n547));
  AOI21_X1  g361(.A(G125), .B1(new_n243), .B2(new_n246), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n229), .A2(G125), .ZN(new_n550));
  INV_X1    g364(.A(new_n546), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n247), .A2(new_n423), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT6), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n539), .A2(new_n555), .A3(new_n541), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n544), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n549), .A2(new_n553), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n540), .B(KEYINPUT8), .Z(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n536), .B2(new_n337), .ZN(new_n562));
  INV_X1    g376(.A(new_n532), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n563), .A2(KEYINPUT87), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n533), .B1(new_n563), .B2(KEYINPUT87), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n535), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n562), .B1(new_n566), .B2(new_n337), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n550), .A2(new_n558), .A3(new_n551), .A4(new_n552), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n560), .A2(new_n543), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n531), .B1(new_n557), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n544), .A2(new_n554), .A3(new_n556), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(new_n570), .A3(new_n530), .A4(new_n569), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(KEYINPUT88), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(G214), .B1(G237), .B2(G902), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT86), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n579), .B(new_n531), .C1(new_n557), .C2(new_n571), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n529), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n191), .A2(G128), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n583), .A2(KEYINPUT23), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n374), .A2(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT23), .ZN(new_n588));
  OAI22_X1  g402(.A1(new_n584), .A2(new_n586), .B1(new_n588), .B2(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G110), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n585), .A2(new_n583), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT24), .B(G110), .Z(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n593), .A2(KEYINPUT74), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(KEYINPUT74), .ZN(new_n595));
  OAI221_X1 g409(.A(new_n590), .B1(new_n594), .B2(new_n595), .C1(new_n466), .C2(new_n467), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n589), .A2(G110), .B1(new_n591), .B2(new_n592), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n431), .A3(new_n440), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT78), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT22), .B(G137), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n596), .A2(new_n598), .A3(new_n603), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT25), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT79), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n300), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n300), .A3(new_n606), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(KEYINPUT79), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n512), .B1(new_n300), .B2(G234), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(G902), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(new_n607), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n316), .A2(new_n399), .A3(new_n582), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT96), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n336), .ZN(G3));
  NAND2_X1  g433(.A1(new_n311), .A2(new_n300), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(G472), .B1(new_n311), .B2(new_n313), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n385), .A2(new_n388), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G469), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n344), .A2(new_n338), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n376), .B2(KEYINPUT10), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n355), .B1(new_n354), .B2(new_n357), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n367), .B1(new_n627), .B2(new_n358), .ZN(new_n628));
  INV_X1    g442(.A(new_n368), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n325), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n392), .A2(KEYINPUT85), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n395), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n320), .A3(new_n300), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n623), .A2(new_n633), .A3(new_n398), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n621), .A2(new_n616), .A3(new_n318), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n514), .A2(KEYINPUT99), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(KEYINPUT33), .C1(new_n515), .C2(new_n517), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n500), .A2(new_n503), .A3(new_n511), .ZN(new_n638));
  INV_X1    g452(.A(new_n513), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n640), .B(new_n514), .C1(KEYINPUT99), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n390), .A2(new_n519), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n518), .A2(new_n519), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT20), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n464), .A2(new_n474), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n572), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(KEYINPUT98), .B(new_n531), .C1(new_n557), .C2(new_n571), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n574), .A2(KEYINPUT97), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n569), .A2(new_n570), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n530), .A4(new_n573), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n578), .ZN(new_n659));
  NOR4_X1   g473(.A1(new_n635), .A2(new_n480), .A3(new_n650), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NAND2_X1  g477(.A1(new_n475), .A2(new_n528), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n664), .A2(new_n480), .A3(new_n521), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n635), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G107), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  NAND2_X1  g484(.A1(new_n613), .A2(new_n614), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n604), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n599), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n615), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n399), .A2(new_n582), .A3(new_n621), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT102), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  AND3_X1   g493(.A1(new_n658), .A2(new_n675), .A3(new_n578), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n477), .B1(new_n478), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n664), .A2(new_n521), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n316), .A2(new_n680), .A3(new_n399), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XOR2_X1   g499(.A(new_n682), .B(KEYINPUT39), .Z(new_n686));
  NAND3_X1  g500(.A1(new_n634), .A2(new_n318), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n690));
  AND3_X1   g504(.A1(new_n575), .A2(new_n580), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n690), .B1(new_n575), .B2(new_n580), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n521), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n664), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n577), .A3(new_n675), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n688), .A2(new_n689), .A3(new_n693), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n307), .A2(new_n308), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n282), .B1(new_n266), .B2(new_n292), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n570), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G472), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n314), .B2(new_n315), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT104), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(new_n701), .C1(new_n314), .C2(new_n315), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n221), .ZN(G45));
  NOR2_X1   g522(.A1(new_n650), .A2(new_n682), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n316), .A2(new_n680), .A3(new_n399), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  NAND2_X1  g525(.A1(new_n632), .A2(new_n300), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n318), .A3(new_n633), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n659), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n650), .A2(new_n480), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n316), .A3(new_n616), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n316), .A3(new_n616), .A4(new_n665), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  AOI21_X1  g535(.A(new_n529), .B1(new_n671), .B2(new_n674), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n316), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  OAI21_X1  g538(.A(new_n281), .B1(new_n263), .B2(new_n293), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n309), .B2(new_n310), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(KEYINPUT105), .A3(new_n313), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(G472), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n311), .B2(new_n300), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT105), .B1(new_n726), .B2(new_n313), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n659), .A2(new_n695), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n714), .A2(new_n480), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n733), .A3(new_n616), .A4(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT106), .B(G122), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G24));
  NAND4_X1  g551(.A1(new_n732), .A2(new_n715), .A3(new_n675), .A4(new_n709), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n314), .B2(new_n315), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n311), .A2(new_n313), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT32), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(KEYINPUT108), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(new_n745), .A3(new_n302), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n577), .B1(new_n575), .B2(new_n580), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n398), .B(KEYINPUT107), .Z(new_n748));
  NAND3_X1  g562(.A1(new_n623), .A2(new_n633), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n749), .A3(new_n318), .ZN(new_n750));
  INV_X1    g564(.A(new_n682), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n664), .A2(new_n647), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n616), .A4(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n747), .A2(new_n749), .A3(new_n318), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n316), .A3(new_n616), .A4(new_n709), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT109), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n754), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n203), .ZN(G33));
  NAND2_X1  g578(.A1(new_n316), .A2(new_n616), .ZN(new_n765));
  INV_X1    g579(.A(new_n664), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n694), .A3(new_n751), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n765), .A2(new_n767), .A3(new_n750), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n211), .ZN(G36));
  INV_X1    g583(.A(new_n621), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n528), .A2(new_n647), .A3(new_n464), .A4(new_n474), .ZN(new_n771));
  NAND2_X1  g585(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n475), .A2(new_n528), .A3(new_n647), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n777), .A4(new_n675), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n747), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n384), .A2(new_n369), .B1(new_n387), .B2(new_n325), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  OAI21_X1  g596(.A(G469), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n385), .A2(new_n388), .A3(new_n782), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT46), .B(new_n748), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT110), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n748), .B1(new_n783), .B2(new_n785), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n622), .A2(KEYINPUT45), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(G469), .A3(new_n784), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT110), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n793), .A3(KEYINPUT46), .A4(new_n748), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n787), .A2(new_n790), .A3(new_n794), .A4(new_n633), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n318), .A3(new_n686), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n778), .A2(new_n797), .A3(new_n747), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n770), .A2(new_n675), .A3(new_n777), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n780), .A2(new_n796), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  INV_X1    g617(.A(new_n747), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n316), .A2(new_n616), .A3(new_n752), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n318), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT47), .B1(new_n795), .B2(new_n318), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND2_X1  g624(.A1(new_n713), .A2(new_n633), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n771), .B1(new_n811), .B2(KEYINPUT49), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(KEYINPUT49), .B2(new_n811), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n813), .A2(new_n319), .A3(new_n577), .A4(new_n693), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n706), .A3(new_n616), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n747), .A2(new_n477), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n714), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n777), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n732), .A2(new_n675), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n777), .A2(new_n477), .ZN(new_n821));
  INV_X1    g635(.A(new_n730), .ZN(new_n822));
  INV_X1    g636(.A(new_n731), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n616), .A4(new_n727), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n577), .B1(new_n691), .B2(new_n692), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(KEYINPUT119), .A3(new_n714), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n828));
  INV_X1    g642(.A(new_n690), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n530), .B1(new_n655), .B2(new_n573), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n580), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n575), .A2(new_n580), .A3(new_n690), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n578), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n714), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n828), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n825), .B1(new_n827), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n825), .B(KEYINPUT50), .C1(new_n827), .C2(new_n838), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n820), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n795), .A2(new_n318), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT47), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n713), .A2(new_n319), .A3(new_n633), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n806), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n821), .A2(new_n824), .A3(new_n804), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n703), .A2(new_n616), .A3(new_n705), .A4(new_n817), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n664), .A2(new_n647), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n843), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n841), .A2(new_n842), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n859));
  INV_X1    g673(.A(new_n820), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n855), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n856), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n820), .B(new_n854), .C1(new_n841), .C2(new_n842), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(new_n850), .C1(new_n859), .C2(KEYINPUT51), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n746), .A2(new_n616), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n818), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT48), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n825), .A2(new_n715), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT120), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n851), .A2(new_n650), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n476), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n862), .A2(new_n864), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n399), .A2(new_n582), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n650), .A2(KEYINPUT113), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n664), .A2(new_n876), .A3(new_n647), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n481), .A2(new_n575), .A3(new_n578), .A4(new_n580), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n765), .A2(new_n874), .B1(new_n635), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT114), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n617), .B(new_n882), .C1(new_n635), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n634), .A2(new_n616), .A3(new_n318), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n621), .A3(new_n665), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n717), .B(new_n676), .C1(new_n581), .C2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n735), .A2(new_n720), .A3(new_n723), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n766), .A2(new_n521), .A3(new_n751), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT115), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n316), .A2(new_n399), .A3(new_n675), .A4(new_n747), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n891), .A2(new_n892), .B1(new_n819), .B2(new_n753), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n884), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n754), .A2(new_n758), .A3(new_n761), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n761), .B1(new_n754), .B2(new_n758), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n896), .A3(new_n768), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n319), .B1(new_n397), .B2(new_n748), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n682), .B(KEYINPUT116), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n675), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n733), .A2(new_n702), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n738), .A2(new_n901), .A3(new_n684), .A4(new_n710), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n634), .A2(new_n318), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n767), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n752), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n316), .B(new_n680), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(KEYINPUT52), .A3(new_n738), .A4(new_n901), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n894), .A2(new_n897), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT53), .ZN(new_n912));
  INV_X1    g726(.A(new_n768), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n760), .A2(new_n762), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n884), .A2(new_n889), .A3(new_n893), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n902), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n902), .A2(new_n917), .A3(KEYINPUT52), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n912), .A2(new_n923), .A3(KEYINPUT54), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n911), .A2(new_n922), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n759), .A2(KEYINPUT53), .A3(new_n913), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n873), .A2(new_n924), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n873), .A2(new_n924), .A3(new_n930), .A4(KEYINPUT121), .ZN(new_n934));
  OR2_X1    g748(.A1(G952), .A2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n815), .B1(new_n933), .B2(new_n936), .ZN(G75));
  NAND2_X1  g751(.A1(new_n925), .A2(new_n929), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n390), .A3(new_n531), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n544), .A2(new_n556), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n554), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n939), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n939), .B2(new_n940), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n277), .A2(G952), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G51));
  XOR2_X1   g761(.A(new_n748), .B(KEYINPUT57), .Z(new_n948));
  AND3_X1   g762(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n926), .B1(new_n925), .B2(new_n929), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n632), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n300), .B1(new_n925), .B2(new_n929), .ZN(new_n954));
  INV_X1    g768(.A(new_n792), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n911), .A2(new_n922), .B1(new_n921), .B2(new_n928), .ZN(new_n957));
  NOR4_X1   g771(.A1(new_n957), .A2(KEYINPUT122), .A3(new_n300), .A4(new_n792), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n946), .B1(new_n952), .B2(new_n959), .ZN(G54));
  NAND3_X1  g774(.A1(new_n954), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n946), .B1(new_n961), .B2(new_n461), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n954), .A2(KEYINPUT58), .A3(G475), .A4(new_n525), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G60));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n643), .B(new_n967), .C1(new_n949), .C2(new_n950), .ZN(new_n968));
  INV_X1    g782(.A(new_n946), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n924), .A2(new_n930), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n643), .B1(new_n971), .B2(new_n967), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n938), .A2(new_n673), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n607), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n957), .B2(new_n975), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n979), .A3(new_n969), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n977), .A2(new_n979), .A3(KEYINPUT61), .A4(new_n969), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(G66));
  INV_X1    g798(.A(new_n479), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n277), .B1(new_n985), .B2(G224), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n884), .A2(new_n889), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n277), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n941), .B1(G898), .B2(new_n277), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n988), .B(new_n989), .Z(G69));
  NAND2_X1  g804(.A1(new_n908), .A2(new_n738), .ZN(new_n991));
  AND2_X1   g805(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n992));
  NOR2_X1   g806(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n993));
  OAI22_X1  g807(.A1(new_n707), .A2(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n908), .A2(new_n738), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n706), .B2(new_n697), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n996), .B2(new_n992), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n875), .A2(new_n877), .B1(new_n694), .B2(new_n766), .ZN(new_n998));
  OR4_X1    g812(.A1(new_n765), .A2(new_n998), .A3(new_n687), .A4(new_n804), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n809), .A2(new_n802), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n277), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n285), .A2(new_n287), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(new_n438), .Z(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n277), .B1(G227), .B2(G900), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n796), .A2(new_n733), .A3(new_n865), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n809), .A2(new_n802), .A3(new_n995), .A4(new_n1007), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1008), .A2(new_n914), .A3(G953), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n681), .A2(new_n277), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1003), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1004), .B(new_n1006), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(KEYINPUT124), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n809), .A2(new_n995), .A3(new_n1007), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n277), .A3(new_n897), .A4(new_n802), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT124), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n1017), .A3(new_n1011), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1014), .A2(new_n1004), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT125), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1019), .A2(new_n1020), .A3(new_n1005), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1020), .B1(new_n1019), .B2(new_n1005), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1013), .B1(new_n1021), .B2(new_n1022), .ZN(G72));
  NOR3_X1   g837(.A1(new_n997), .A2(new_n987), .A3(new_n1000), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT63), .Z(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n282), .B(new_n289), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n290), .B(KEYINPUT127), .ZN(new_n1029));
  INV_X1    g843(.A(new_n698), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n912), .A2(new_n923), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  OR3_X1    g847(.A1(new_n1008), .A2(new_n914), .A3(new_n987), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n1026), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n289), .A2(new_n282), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n969), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1037), .A2(KEYINPUT126), .A3(new_n969), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1033), .B1(new_n1040), .B2(new_n1041), .ZN(G57));
endmodule


