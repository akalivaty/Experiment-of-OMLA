

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  NOR2_X1 U321 ( .A1(n498), .A2(n582), .ZN(n420) );
  INV_X1 U322 ( .A(n354), .ZN(n353) );
  INV_X1 U323 ( .A(KEYINPUT41), .ZN(n289) );
  NOR2_X1 U324 ( .A1(n525), .A2(n431), .ZN(n569) );
  NOR2_X1 U325 ( .A1(n425), .A2(n424), .ZN(n426) );
  XNOR2_X1 U326 ( .A(n428), .B(KEYINPUT54), .ZN(n429) );
  XOR2_X1 U327 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n384) );
  XNOR2_X1 U328 ( .A(G204GAT), .B(G92GAT), .ZN(n316) );
  XNOR2_X1 U329 ( .A(n419), .B(n289), .ZN(n556) );
  XNOR2_X2 U330 ( .A(KEYINPUT122), .B(n290), .ZN(n566) );
  AND2_X1 U331 ( .A1(n462), .A2(n541), .ZN(n290) );
  XOR2_X1 U332 ( .A(n461), .B(n460), .Z(n541) );
  XNOR2_X2 U333 ( .A(n376), .B(n375), .ZN(n419) );
  XOR2_X1 U334 ( .A(KEYINPUT45), .B(n420), .Z(n291) );
  INV_X1 U335 ( .A(G162GAT), .ZN(n406) );
  XNOR2_X1 U336 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U337 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U338 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U339 ( .A(n414), .B(n413), .Z(n469) );
  XOR2_X1 U340 ( .A(n480), .B(KEYINPUT28), .Z(n532) );
  XNOR2_X1 U341 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n463) );
  XNOR2_X1 U342 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n449) );
  XOR2_X1 U344 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n293) );
  XNOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT83), .ZN(n292) );
  XNOR2_X1 U346 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U347 ( .A(n294), .B(G127GAT), .Z(n296) );
  XNOR2_X1 U348 ( .A(G113GAT), .B(G120GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n461) );
  XOR2_X1 U350 ( .A(G85GAT), .B(G57GAT), .Z(n359) );
  XOR2_X1 U351 ( .A(KEYINPUT95), .B(n359), .Z(n298) );
  XOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT78), .Z(n409) );
  XNOR2_X1 U353 ( .A(G148GAT), .B(n409), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U355 ( .A(n461), .B(n299), .Z(n301) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(KEYINPUT98), .Z(n303) );
  XNOR2_X1 U359 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U361 ( .A(n305), .B(n304), .Z(n313) );
  XOR2_X1 U362 ( .A(KEYINPUT3), .B(G162GAT), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U365 ( .A(G141GAT), .B(n308), .Z(n441) );
  XOR2_X1 U366 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n310) );
  XNOR2_X1 U367 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n441), .B(n311), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n479) );
  XOR2_X1 U371 ( .A(KEYINPUT99), .B(n479), .Z(n525) );
  XOR2_X1 U372 ( .A(G36GAT), .B(G8GAT), .Z(n315) );
  NAND2_X1 U373 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n316), .B(G64GAT), .ZN(n354) );
  INV_X1 U376 ( .A(n353), .ZN(n317) );
  XOR2_X1 U377 ( .A(n318), .B(n317), .Z(n330) );
  XOR2_X1 U378 ( .A(G176GAT), .B(G183GAT), .Z(n320) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U381 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n322) );
  XNOR2_X1 U382 ( .A(G190GAT), .B(KEYINPUT86), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U384 ( .A(n324), .B(n323), .Z(n457) );
  XNOR2_X1 U385 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n325), .B(KEYINPUT21), .ZN(n326) );
  XOR2_X1 U387 ( .A(n326), .B(KEYINPUT91), .Z(n328) );
  XNOR2_X1 U388 ( .A(G197GAT), .B(G218GAT), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n443) );
  XNOR2_X1 U390 ( .A(n457), .B(n443), .ZN(n329) );
  XOR2_X1 U391 ( .A(n330), .B(n329), .Z(n527) );
  INV_X1 U392 ( .A(n527), .ZN(n427) );
  XOR2_X1 U393 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n378) );
  XOR2_X1 U394 ( .A(KEYINPUT29), .B(G141GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G197GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U397 ( .A(G29GAT), .B(G113GAT), .Z(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n347) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n335), .B(G36GAT), .ZN(n336) );
  XOR2_X1 U401 ( .A(n336), .B(KEYINPUT8), .Z(n338) );
  XNOR2_X1 U402 ( .A(G50GAT), .B(KEYINPUT67), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n399) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G15GAT), .Z(n340) );
  XNOR2_X1 U405 ( .A(G8GAT), .B(KEYINPUT68), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U407 ( .A(G1GAT), .B(n341), .Z(n391) );
  XNOR2_X1 U408 ( .A(n399), .B(n391), .ZN(n345) );
  XOR2_X1 U409 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n343) );
  XNOR2_X1 U410 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U412 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n347), .B(n346), .ZN(n349) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XOR2_X1 U415 ( .A(n349), .B(n348), .Z(n511) );
  INV_X1 U416 ( .A(n511), .ZN(n570) );
  XOR2_X1 U417 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n351) );
  XNOR2_X1 U418 ( .A(KEYINPUT76), .B(KEYINPUT71), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n376) );
  XOR2_X1 U420 ( .A(G99GAT), .B(G71GAT), .Z(n450) );
  INV_X1 U421 ( .A(n450), .ZN(n352) );
  NAND2_X1 U422 ( .A1(n353), .A2(n352), .ZN(n356) );
  NAND2_X1 U423 ( .A1(n354), .A2(n450), .ZN(n355) );
  NAND2_X1 U424 ( .A1(n356), .A2(n355), .ZN(n358) );
  AND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U427 ( .A(KEYINPUT33), .B(n384), .Z(n361) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U429 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n367) );
  INV_X1 U431 ( .A(n367), .ZN(n365) );
  XOR2_X1 U432 ( .A(G120GAT), .B(KEYINPUT73), .Z(n366) );
  INV_X1 U433 ( .A(n366), .ZN(n364) );
  NAND2_X1 U434 ( .A1(n365), .A2(n364), .ZN(n369) );
  NAND2_X1 U435 ( .A1(n367), .A2(n366), .ZN(n368) );
  NAND2_X1 U436 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n370), .B(KEYINPUT75), .ZN(n374) );
  XOR2_X1 U438 ( .A(G78GAT), .B(G148GAT), .Z(n372) );
  XNOR2_X1 U439 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n438) );
  XOR2_X1 U441 ( .A(n438), .B(KEYINPUT32), .Z(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n375) );
  NAND2_X1 U443 ( .A1(n570), .A2(n556), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n416) );
  XOR2_X1 U445 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n380) );
  XNOR2_X1 U446 ( .A(G57GAT), .B(G64GAT), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n395) );
  XOR2_X1 U448 ( .A(G78GAT), .B(G155GAT), .Z(n382) );
  XNOR2_X1 U449 ( .A(G71GAT), .B(G211GAT), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U451 ( .A(n384), .B(n383), .Z(n386) );
  XNOR2_X1 U452 ( .A(G127GAT), .B(G183GAT), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U454 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n388) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U457 ( .A(n390), .B(n389), .Z(n393) );
  XNOR2_X1 U458 ( .A(n391), .B(KEYINPUT15), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U460 ( .A(n395), .B(n394), .Z(n498) );
  INV_X1 U461 ( .A(n498), .ZN(n579) );
  XOR2_X1 U462 ( .A(KEYINPUT73), .B(KEYINPUT77), .Z(n397) );
  XNOR2_X1 U463 ( .A(KEYINPUT64), .B(KEYINPUT9), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n414) );
  XOR2_X1 U466 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n401) );
  XNOR2_X1 U467 ( .A(G190GAT), .B(G218GAT), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U469 ( .A(G92GAT), .B(G85GAT), .Z(n403) );
  XNOR2_X1 U470 ( .A(G99GAT), .B(G106GAT), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U472 ( .A(n405), .B(n404), .Z(n412) );
  NAND2_X1 U473 ( .A1(G232GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U474 ( .A(G134GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  INV_X1 U476 ( .A(n469), .ZN(n562) );
  NOR2_X1 U477 ( .A1(n579), .A2(n562), .ZN(n415) );
  NAND2_X1 U478 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n417), .B(KEYINPUT47), .ZN(n418) );
  XNOR2_X1 U480 ( .A(KEYINPUT112), .B(n418), .ZN(n425) );
  XNOR2_X1 U481 ( .A(KEYINPUT36), .B(n469), .ZN(n582) );
  NOR2_X1 U482 ( .A1(n419), .A2(n291), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n421), .B(KEYINPUT113), .ZN(n422) );
  NOR2_X1 U484 ( .A1(n570), .A2(n422), .ZN(n423) );
  XNOR2_X1 U485 ( .A(KEYINPUT114), .B(n423), .ZN(n424) );
  XNOR2_X1 U486 ( .A(KEYINPUT48), .B(n426), .ZN(n537) );
  NOR2_X1 U487 ( .A1(n427), .A2(n537), .ZN(n430) );
  XNOR2_X1 U488 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n428) );
  XOR2_X1 U489 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U490 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U492 ( .A(KEYINPUT89), .B(KEYINPUT94), .Z(n435) );
  XNOR2_X1 U493 ( .A(G204GAT), .B(KEYINPUT92), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n447) );
  XOR2_X1 U496 ( .A(KEYINPUT22), .B(n438), .Z(n440) );
  NAND2_X1 U497 ( .A1(G228GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U499 ( .A(n442), .B(n441), .Z(n445) );
  XNOR2_X1 U500 ( .A(G50GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n480) );
  NAND2_X1 U503 ( .A1(n569), .A2(n480), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n462) );
  XOR2_X1 U505 ( .A(KEYINPUT87), .B(n450), .Z(n452) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U508 ( .A(n453), .B(KEYINPUT20), .Z(n459) );
  XOR2_X1 U509 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n455) );
  XNOR2_X1 U510 ( .A(G43GAT), .B(G15GAT), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U514 ( .A1(n566), .A2(n562), .ZN(n464) );
  NAND2_X1 U515 ( .A1(n566), .A2(n556), .ZN(n468) );
  XOR2_X1 U516 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n466) );
  XOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT56), .Z(n465) );
  XNOR2_X1 U518 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U519 ( .A(n468), .B(n467), .ZN(G1349GAT) );
  OR2_X1 U520 ( .A1(n511), .A2(n419), .ZN(n501) );
  XOR2_X1 U521 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n471) );
  NAND2_X1 U522 ( .A1(n579), .A2(n469), .ZN(n470) );
  XNOR2_X1 U523 ( .A(n471), .B(n470), .ZN(n486) );
  NAND2_X1 U524 ( .A1(n541), .A2(n527), .ZN(n472) );
  NAND2_X1 U525 ( .A1(n480), .A2(n472), .ZN(n473) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n473), .Z(n476) );
  XNOR2_X1 U527 ( .A(n527), .B(KEYINPUT27), .ZN(n482) );
  NOR2_X1 U528 ( .A1(n480), .A2(n541), .ZN(n474) );
  XOR2_X1 U529 ( .A(n474), .B(KEYINPUT26), .Z(n553) );
  INV_X1 U530 ( .A(n553), .ZN(n568) );
  NAND2_X1 U531 ( .A1(n482), .A2(n568), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT100), .B(n477), .Z(n478) );
  NOR2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n485) );
  XOR2_X1 U535 ( .A(n541), .B(KEYINPUT88), .Z(n481) );
  INV_X1 U536 ( .A(n532), .ZN(n540) );
  NAND2_X1 U537 ( .A1(n481), .A2(n540), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n525), .A2(n482), .ZN(n538) );
  NOR2_X1 U539 ( .A1(n483), .A2(n538), .ZN(n484) );
  NOR2_X1 U540 ( .A1(n485), .A2(n484), .ZN(n497) );
  NOR2_X1 U541 ( .A1(n486), .A2(n497), .ZN(n487) );
  XNOR2_X1 U542 ( .A(n487), .B(KEYINPUT101), .ZN(n512) );
  NOR2_X1 U543 ( .A1(n501), .A2(n512), .ZN(n495) );
  NAND2_X1 U544 ( .A1(n495), .A2(n525), .ZN(n488) );
  XNOR2_X1 U545 ( .A(n488), .B(KEYINPUT34), .ZN(n489) );
  XOR2_X1 U546 ( .A(n489), .B(KEYINPUT102), .Z(n491) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(KEYINPUT103), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n527), .A2(n495), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U552 ( .A1(n495), .A2(n541), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n532), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NOR2_X1 U557 ( .A1(n582), .A2(n497), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n499), .A2(n498), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT37), .B(n500), .Z(n524) );
  NOR2_X1 U560 ( .A1(n524), .A2(n501), .ZN(n502) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(n502), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n525), .A2(n509), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U564 ( .A(KEYINPUT104), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U565 ( .A1(n509), .A2(n527), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n509), .A2(n541), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n507), .B(KEYINPUT40), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U570 ( .A1(n532), .A2(n509), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n514) );
  NAND2_X1 U573 ( .A1(n511), .A2(n556), .ZN(n523) );
  NOR2_X1 U574 ( .A1(n512), .A2(n523), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n520), .A2(n525), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n527), .A2(n520), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n517), .ZN(G1333GAT) );
  XOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U582 ( .A1(n520), .A2(n541), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n522) );
  NAND2_X1 U585 ( .A1(n520), .A2(n532), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NOR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n525), .A2(n533), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n533), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n530) );
  NAND2_X1 U593 ( .A1(n533), .A2(n541), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n535) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  NOR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n539), .B(KEYINPUT115), .ZN(n552) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U603 ( .A1(n552), .A2(n542), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n548), .A2(n570), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U607 ( .A1(n548), .A2(n556), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n579), .A2(n548), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n550) );
  NAND2_X1 U613 ( .A1(n548), .A2(n562), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  XOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT117), .Z(n555) );
  NOR2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n563), .A2(n570), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(G1344GAT) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n560) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  NAND2_X1 U622 ( .A1(n563), .A2(n556), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n579), .A2(n563), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n570), .A2(n566), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n579), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n581) );
  INV_X1 U634 ( .A(n581), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n578), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n576) );
  NAND2_X1 U641 ( .A1(n578), .A2(n419), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(G218GAT), .B(n585), .Z(G1355GAT) );
endmodule

