//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n211), .B1(new_n214), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n225), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n218), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n244), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n212), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n205), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G68), .ZN(new_n258));
  OR3_X1    g0058(.A1(new_n256), .A2(KEYINPUT72), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT72), .B1(new_n256), .B2(new_n258), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n255), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n218), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT12), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n267), .A2(new_n268), .B1(new_n206), .B2(G68), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n269), .A2(KEYINPUT71), .B1(new_n245), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n253), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT11), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n261), .B(new_n264), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n274), .A2(new_n275), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT14), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  AND2_X1   g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n212), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n219), .B1(new_n290), .B2(KEYINPUT70), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n285), .B1(new_n212), .B2(new_n282), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n286), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT3), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G33), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n296), .A2(new_n298), .A3(G232), .A4(G1698), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n296), .A2(new_n298), .A3(G226), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n283), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n281), .B1(new_n295), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(G1), .B(G13), .C1(new_n265), .C2(new_n287), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(KEYINPUT70), .A3(new_n285), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n294), .A2(new_n307), .A3(G238), .ZN(new_n308));
  INV_X1    g0108(.A(new_n286), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n280), .B(G169), .C1(new_n305), .C2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n295), .A2(new_n281), .A3(new_n304), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G179), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n314), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n280), .B1(new_n317), .B2(G169), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n279), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(G200), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n313), .A2(G190), .A3(new_n314), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n278), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g0123(.A(new_n323), .B(KEYINPUT73), .Z(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT8), .B(G58), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n325), .A2(new_n267), .B1(new_n326), .B2(new_n271), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n206), .B1(new_n201), .B2(new_n245), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n253), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT66), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT66), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n257), .A2(G50), .ZN(new_n332));
  XOR2_X1   g0132(.A(new_n332), .B(KEYINPUT67), .Z(new_n333));
  INV_X1    g0133(.A(new_n256), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n333), .A2(new_n334), .B1(new_n245), .B2(new_n262), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT9), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT68), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT3), .B(G33), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(G222), .A3(new_n300), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(G1698), .ZN(new_n342));
  INV_X1    g0142(.A(G223), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n341), .B1(new_n268), .B2(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n283), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n286), .B1(G226), .B2(new_n290), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n337), .A2(new_n336), .B1(new_n348), .B2(G190), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(G200), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT10), .B1(new_n339), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n350), .A2(KEYINPUT69), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT10), .B1(new_n350), .B2(KEYINPUT69), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n352), .B1(new_n339), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n336), .C1(G179), .C2(new_n347), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n325), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n257), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n362), .A2(new_n256), .B1(new_n255), .B2(new_n361), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT77), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  INV_X1    g0166(.A(G159), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n271), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n270), .A2(KEYINPUT75), .A3(G159), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n224), .A2(new_n218), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n201), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n265), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n379), .B2(new_n298), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n296), .A2(new_n298), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n381), .B2(new_n206), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT76), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n373), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT76), .B(G68), .C1(new_n380), .C2(new_n382), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n370), .A2(new_n372), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n297), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(G33), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n296), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n393), .B2(new_n374), .ZN(new_n394));
  INV_X1    g0194(.A(new_n296), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n377), .A2(new_n378), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(G33), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n397), .A2(KEYINPUT7), .A3(G20), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT16), .B(new_n388), .C1(new_n394), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n253), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n365), .B1(new_n387), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n309), .B1(new_n225), .B2(new_n292), .ZN(new_n403));
  MUX2_X1   g0203(.A(G223), .B(G226), .S(G1698), .Z(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n392), .A3(new_n296), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n306), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G179), .ZN(new_n409));
  OAI21_X1  g0209(.A(G169), .B1(new_n403), .B2(new_n407), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n401), .A2(new_n402), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n402), .B1(new_n401), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n286), .B1(G232), .B2(new_n290), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n405), .A2(new_n406), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(new_n306), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n408), .B2(G200), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n365), .B(new_n419), .C1(new_n387), .C2(new_n400), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n257), .A2(G77), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n256), .A2(new_n423), .B1(G77), .B2(new_n255), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n361), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n425), .B1(new_n267), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n424), .B1(new_n430), .B2(new_n253), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n342), .A2(new_n219), .B1(new_n432), .B2(new_n340), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n381), .A2(new_n225), .A3(G1698), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n283), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n286), .B1(G244), .B2(new_n290), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n431), .B1(new_n437), .B2(new_n357), .ZN(new_n438));
  INV_X1    g0238(.A(new_n437), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G200), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n431), .B1(new_n437), .B2(new_n416), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n324), .A2(new_n360), .A3(new_n422), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT83), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n205), .A2(G33), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n255), .A2(new_n450), .A3(new_n212), .A4(new_n252), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n220), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT82), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT81), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT19), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n266), .A2(new_n455), .A3(G97), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G97), .A2(G107), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n457), .A2(new_n220), .B1(new_n302), .B2(new_n206), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n455), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n392), .A2(new_n206), .A3(G68), .A4(new_n296), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n253), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n428), .A2(new_n255), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n454), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n254), .B1(new_n459), .B2(new_n460), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n466), .A2(KEYINPUT81), .A3(new_n463), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n453), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n283), .A2(new_n284), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n288), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n205), .A2(G45), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n306), .A2(G250), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n219), .A2(G1698), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n392), .A2(new_n296), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n392), .A2(G244), .A3(G1698), .A4(new_n296), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n392), .A2(new_n480), .A3(new_n296), .A4(new_n475), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n474), .B1(new_n482), .B2(new_n283), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n443), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n416), .B(new_n474), .C1(new_n482), .C2(new_n283), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n468), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n462), .A2(new_n454), .A3(new_n464), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT81), .B1(new_n466), .B2(new_n463), .ZN(new_n488));
  INV_X1    g0288(.A(new_n451), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n487), .A2(new_n488), .B1(new_n428), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n482), .A2(new_n283), .ZN(new_n491));
  INV_X1    g0291(.A(new_n474), .ZN(new_n492));
  AOI21_X1  g0292(.A(G169), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI211_X1 g0293(.A(G179), .B(new_n474), .C1(new_n482), .C2(new_n283), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n449), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  INV_X1    g0297(.A(new_n490), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n453), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n487), .B2(new_n488), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n483), .A2(G190), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(new_n443), .C2(new_n483), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT83), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G257), .A2(G1698), .ZN(new_n506));
  INV_X1    g0306(.A(G264), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n392), .A3(new_n296), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n381), .A2(G303), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n306), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n472), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(G274), .A3(new_n306), .ZN(new_n515));
  INV_X1    g0315(.A(new_n513), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n470), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(G270), .A3(new_n306), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(G169), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n255), .A2(G116), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n451), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(G20), .B1(new_n265), .B2(G97), .ZN(new_n526));
  NAND3_X1  g0326(.A1(KEYINPUT78), .A2(G33), .A3(G283), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT78), .B1(G33), .B2(G283), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n252), .A2(new_n212), .B1(G20), .B2(new_n524), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(KEYINPUT20), .A3(new_n531), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n525), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n521), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n522), .B1(new_n489), .B2(G116), .ZN(new_n538));
  INV_X1    g0338(.A(new_n535), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT20), .B1(new_n530), .B2(new_n531), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n511), .A2(new_n520), .A3(new_n440), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n537), .A2(KEYINPUT21), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT84), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT21), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n521), .B2(new_n536), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n515), .A2(new_n519), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n509), .A2(new_n510), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(G190), .C1(new_n548), .C2(new_n306), .ZN(new_n549));
  OAI21_X1  g0349(.A(G200), .B1(new_n511), .B2(new_n520), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n536), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n543), .A2(new_n544), .A3(new_n546), .A4(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n547), .B1(new_n548), .B2(new_n306), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(KEYINPUT21), .A3(G169), .A4(new_n541), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n542), .A2(new_n541), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n551), .A2(new_n554), .A3(new_n546), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT84), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(new_n432), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n432), .A3(G20), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n561), .A2(KEYINPUT86), .B1(new_n562), .B2(G20), .ZN(new_n563));
  AOI211_X1 g0363(.A(new_n560), .B(new_n563), .C1(KEYINPUT86), .C2(new_n561), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n220), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n392), .A2(new_n206), .A3(new_n296), .A4(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT85), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n206), .A2(G87), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n565), .B1(new_n381), .B2(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n567), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n564), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT24), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n564), .B(new_n575), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n253), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n255), .A2(G107), .ZN(new_n579));
  XNOR2_X1  g0379(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n579), .B(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n432), .B2(new_n451), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G250), .A2(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n227), .B2(G1698), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n397), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G294), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n306), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n518), .A2(G264), .A3(new_n306), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n515), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G190), .ZN(new_n592));
  OAI21_X1  g0392(.A(G200), .B1(new_n588), .B2(new_n590), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n578), .A2(new_n583), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n591), .A2(G169), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n440), .B2(new_n591), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n254), .B1(new_n574), .B2(new_n576), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(new_n582), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n255), .A2(G97), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n489), .B2(G97), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT6), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n603), .A2(new_n226), .A3(G107), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(G20), .B1(G77), .B2(new_n270), .ZN(new_n608));
  OAI21_X1  g0408(.A(G107), .B1(new_n380), .B2(new_n382), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n254), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n518), .A2(G257), .A3(new_n306), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n296), .A2(new_n298), .A3(G250), .A4(G1698), .ZN(new_n612));
  AND2_X1   g0412(.A1(KEYINPUT4), .A2(G244), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n296), .A2(new_n298), .A3(new_n613), .A4(new_n300), .ZN(new_n614));
  NAND2_X1  g0414(.A1(G33), .A2(G283), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT78), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n527), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n612), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT4), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n392), .A2(G244), .A3(new_n300), .A4(new_n296), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n515), .B(new_n611), .C1(new_n622), .C2(new_n306), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n601), .B(new_n610), .C1(new_n623), .C2(G200), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n623), .A2(new_n416), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT79), .B1(new_n610), .B2(new_n601), .ZN(new_n626));
  AOI21_X1  g0426(.A(G33), .B1(new_n390), .B2(new_n391), .ZN(new_n627));
  INV_X1    g0427(.A(new_n298), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n375), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n374), .B1(new_n340), .B2(G20), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n432), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n605), .B1(new_n603), .B2(new_n602), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n632), .A2(new_n206), .B1(new_n268), .B2(new_n271), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n253), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT79), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n600), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n626), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(G169), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n621), .A2(new_n620), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n283), .B1(new_n639), .B2(new_n619), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(G179), .A3(new_n515), .A4(new_n611), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n624), .A2(new_n625), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n558), .A2(new_n594), .A3(new_n598), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n448), .A2(new_n505), .A3(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n318), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n315), .A3(new_n312), .ZN(new_n647));
  INV_X1    g0447(.A(new_n442), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n279), .B1(new_n648), .B2(new_n322), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n421), .B1(new_n649), .B2(KEYINPUT90), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(KEYINPUT90), .B2(new_n649), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n412), .B2(new_n413), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n401), .A2(new_n411), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT18), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n401), .A2(new_n402), .A3(new_n411), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(KEYINPUT89), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n356), .B1(new_n651), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n359), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n637), .A2(new_n642), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT26), .B1(new_n505), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n483), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(KEYINPUT88), .A3(G200), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n483), .B2(new_n443), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n667), .A3(new_n502), .A4(new_n501), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n499), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n543), .A2(new_n546), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n598), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n669), .A2(new_n671), .A3(new_n594), .A4(new_n643), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n610), .A2(new_n601), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n638), .B2(new_n641), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n668), .A2(new_n499), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n499), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n663), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n661), .B1(new_n448), .B2(new_n680), .ZN(G369));
  NAND3_X1  g0481(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n536), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT91), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n558), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n552), .A2(new_n557), .A3(KEYINPUT91), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n691), .A2(new_n692), .B1(new_n670), .B2(new_n689), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n578), .A2(new_n583), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n596), .A3(new_n688), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n687), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n594), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n598), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n670), .A2(new_n687), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n697), .A3(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n209), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR4_X1   g0508(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n215), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n496), .A2(new_n504), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n643), .A2(new_n594), .A3(new_n598), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(new_n558), .A4(new_n688), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n591), .A2(new_n542), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n640), .A2(new_n611), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n483), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n591), .A2(new_n542), .A3(new_n640), .A4(new_n611), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n664), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n591), .A2(G179), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n664), .A3(new_n553), .A4(new_n623), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n687), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n713), .B1(new_n716), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT92), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(KEYINPUT92), .B(new_n713), .C1(new_n716), .C2(new_n730), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n499), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n495), .A2(KEYINPUT93), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n668), .A2(new_n499), .A3(new_n675), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(KEYINPUT26), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n662), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n496), .A2(new_n504), .A3(new_n673), .A4(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(new_n672), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT29), .A3(new_n688), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n680), .A2(new_n687), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n746), .B1(new_n747), .B2(KEYINPUT29), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n736), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n712), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(G13), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n205), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n707), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n695), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n693), .A2(G330), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n693), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n212), .B1(G20), .B2(new_n357), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n206), .A2(G179), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n367), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n206), .A2(new_n440), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n218), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n220), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n767), .A2(new_n416), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n432), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n416), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n206), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n226), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n775), .A2(G190), .A3(new_n443), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n776), .A2(new_n416), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n340), .B1(new_n224), .B2(new_n788), .C1(new_n790), .C2(new_n245), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n775), .A2(new_n768), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(KEYINPUT95), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n791), .B1(G77), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n774), .A2(new_n787), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n785), .ZN(new_n799));
  INV_X1    g0599(.A(new_n792), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(G294), .B1(new_n800), .B2(G311), .ZN(new_n801));
  INV_X1    g0601(.A(G326), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n790), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT97), .ZN(new_n804));
  INV_X1    g0604(.A(new_n772), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G329), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n381), .B1(new_n788), .B2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(KEYINPUT33), .B(G317), .Z(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n778), .A2(new_n809), .B1(new_n782), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n780), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n808), .B(new_n811), .C1(G303), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n804), .A2(new_n806), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n766), .B1(new_n798), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n756), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n209), .A2(G355), .A3(new_n340), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n706), .A2(new_n397), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n216), .B2(G45), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n250), .A2(new_n288), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n817), .B1(G116), .B2(new_n209), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n762), .A2(new_n765), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT94), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n815), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n757), .A2(new_n759), .B1(new_n764), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NOR2_X1   g0629(.A1(new_n442), .A2(new_n687), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n444), .A2(new_n445), .B1(new_n431), .B2(new_n688), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n442), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n446), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n688), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n747), .A2(new_n835), .B1(new_n680), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n756), .B1(new_n736), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n736), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n782), .A2(new_n220), .ZN(new_n841));
  INV_X1    g0641(.A(G303), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n810), .A2(new_n778), .B1(new_n790), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(G107), .C2(new_n812), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n805), .A2(G311), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n796), .A2(G116), .ZN(new_n846));
  INV_X1    g0646(.A(new_n788), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n340), .B(new_n786), .C1(G294), .C2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n397), .B1(new_n224), .B2(new_n785), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n805), .B2(G132), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n245), .A2(new_n780), .B1(new_n782), .B2(new_n218), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT98), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G137), .A2(new_n789), .B1(new_n847), .B2(G143), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n854), .B1(new_n326), .B2(new_n778), .C1(new_n795), .C2(new_n367), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT34), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n851), .B(new_n853), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n855), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT34), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n849), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n765), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n765), .A2(new_n760), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n816), .B1(new_n268), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n835), .C2(new_n761), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n840), .A2(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n753), .A2(new_n205), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT102), .ZN(new_n867));
  INV_X1    g0667(.A(new_n322), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n279), .B(new_n687), .C1(new_n647), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n279), .A2(new_n687), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n319), .A2(new_n322), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n834), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n644), .A2(new_n505), .A3(new_n687), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n728), .A2(new_n729), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n377), .A2(new_n378), .A3(new_n265), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n206), .B1(new_n878), .B2(new_n395), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n218), .B1(new_n879), .B2(KEYINPUT7), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n393), .A2(new_n374), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n373), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n254), .B1(new_n882), .B2(KEYINPUT16), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT16), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n218), .B1(new_n629), .B2(new_n630), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n388), .B1(new_n885), .B2(KEYINPUT76), .ZN(new_n886));
  INV_X1    g0686(.A(new_n386), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n364), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n411), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n420), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n889), .B2(new_n685), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n877), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n685), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT37), .B1(new_n401), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n896), .A2(KEYINPUT99), .A3(new_n654), .A4(new_n420), .ZN(new_n897));
  INV_X1    g0697(.A(new_n363), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n882), .A2(KEYINPUT16), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n400), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n411), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n895), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(new_n420), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n894), .A2(new_n897), .B1(KEYINPUT37), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n902), .B1(new_n414), .B2(new_n421), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n876), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n894), .A2(new_n897), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n905), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n875), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n867), .B1(new_n912), .B2(KEYINPUT40), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n319), .A2(new_n322), .A3(new_n870), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n870), .B1(new_n319), .B2(new_n322), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n835), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n716), .B2(new_n730), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n909), .B2(new_n910), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n904), .A2(new_n905), .A3(new_n876), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(KEYINPUT102), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n401), .A2(new_n895), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n658), .B2(new_n421), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n654), .A2(new_n924), .A3(new_n420), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n894), .A2(new_n897), .B1(new_n926), .B2(KEYINPUT37), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n876), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n911), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n875), .A2(new_n921), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n923), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT103), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n716), .A2(new_n730), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n447), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n713), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n933), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n911), .A2(new_n906), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT39), .ZN(new_n940));
  XNOR2_X1  g0740(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n928), .A2(new_n911), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n647), .A2(new_n279), .A3(new_n688), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n837), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n830), .B1(new_n679), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n914), .A2(new_n915), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n950), .A2(new_n939), .B1(new_n659), .B2(new_n685), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n946), .A2(new_n951), .A3(KEYINPUT101), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT101), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n944), .B1(new_n940), .B2(new_n942), .ZN(new_n954));
  INV_X1    g0754(.A(new_n949), .ZN(new_n955));
  AND4_X1   g0755(.A1(new_n499), .A2(new_n643), .A3(new_n594), .A4(new_n668), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n677), .B1(new_n956), .B2(new_n671), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n837), .B1(new_n957), .B2(new_n663), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n955), .B1(new_n958), .B2(new_n830), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n918), .A2(new_n919), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n959), .A2(new_n960), .B1(new_n658), .B2(new_n895), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n953), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n447), .B(new_n746), .C1(KEYINPUT29), .C2(new_n747), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n661), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n963), .B(new_n965), .Z(new_n966));
  AOI21_X1  g0766(.A(new_n866), .B1(new_n938), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n938), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n524), .B(new_n214), .C1(new_n607), .C2(KEYINPUT35), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(KEYINPUT35), .B2(new_n607), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT36), .ZN(new_n971));
  OAI21_X1  g0771(.A(G77), .B1(new_n224), .B2(new_n218), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n246), .B1(new_n215), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(G1), .A3(new_n752), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n968), .A2(new_n971), .A3(new_n974), .ZN(G367));
  OAI21_X1  g0775(.A(new_n643), .B1(new_n674), .B2(new_n688), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n675), .A2(new_n687), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n701), .A2(new_n703), .A3(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  INV_X1    g0780(.A(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n662), .B1(new_n981), .B2(new_n598), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n688), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n468), .A2(new_n687), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n669), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n499), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT104), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n990), .A2(KEYINPUT104), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n994), .B1(new_n992), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n702), .A2(new_n981), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT105), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT105), .B2(new_n1000), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1000), .A2(KEYINPUT105), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n704), .A2(new_n697), .A3(new_n978), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT45), .Z(new_n1007));
  AOI21_X1  g0807(.A(new_n978), .B1(new_n704), .B2(new_n697), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT44), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(new_n702), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n701), .B(new_n703), .Z(new_n1012));
  INV_X1    g0812(.A(KEYINPUT106), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n695), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n694), .B(KEYINPUT106), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n1012), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n749), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n707), .B(KEYINPUT41), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n754), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1003), .A2(new_n1005), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n818), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n822), .B1(new_n209), .B2(new_n429), .C1(new_n1021), .C2(new_n240), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1022), .A2(new_n756), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n397), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n432), .B2(new_n785), .ZN(new_n1025));
  INV_X1    g0825(.A(G294), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n778), .A2(new_n1026), .B1(new_n782), .B2(new_n226), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n789), .A2(G311), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n842), .B2(new_n788), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1025), .B(new_n1027), .C1(KEYINPUT107), .C2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT107), .B2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n805), .A2(G317), .B1(new_n796), .B2(G283), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n812), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT46), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n780), .B2(new_n524), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n785), .A2(new_n218), .B1(new_n788), .B2(new_n326), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT108), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n778), .A2(new_n367), .B1(new_n782), .B2(new_n268), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G143), .B2(new_n789), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n796), .A2(G50), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n805), .A2(G137), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n381), .B1(new_n812), .B2(G58), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1031), .A2(new_n1036), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT47), .Z(new_n1046));
  OAI221_X1 g0846(.A(new_n1023), .B1(new_n988), .B2(new_n763), .C1(new_n766), .C2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT109), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1020), .A2(new_n1049), .ZN(G387));
  NAND2_X1  g0850(.A1(new_n237), .A2(G45), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT110), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1053));
  NOR3_X1   g0853(.A1(new_n1053), .A2(G50), .A3(new_n325), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n709), .B(new_n288), .C1(new_n218), .C2(new_n268), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1053), .B1(G50), .B2(new_n325), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1021), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1052), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n209), .A2(new_n340), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(G107), .B2(new_n209), .C1(new_n709), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n822), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n756), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n701), .A2(new_n763), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n367), .A2(new_n790), .B1(new_n778), .B2(new_n325), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G77), .B2(new_n812), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n805), .A2(G150), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n788), .A2(new_n245), .B1(new_n792), .B2(new_n218), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1024), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n782), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n799), .A2(new_n428), .B1(new_n1070), .B2(G97), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n397), .B1(G116), .B2(new_n1070), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n785), .A2(new_n810), .B1(new_n780), .B2(new_n1026), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G311), .A2(new_n777), .B1(new_n847), .B2(G317), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n807), .B2(new_n790), .C1(new_n795), .C2(new_n842), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1073), .B1(new_n802), .B2(new_n772), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1072), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1063), .B(new_n1064), .C1(new_n765), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1016), .B2(new_n755), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n750), .A2(new_n1016), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n707), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n750), .A2(new_n1016), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(G393));
  OAI221_X1 g0889(.A(new_n822), .B1(new_n226), .B2(new_n209), .C1(new_n1021), .C2(new_n244), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n756), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1024), .B(new_n841), .C1(new_n796), .C2(new_n361), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n780), .A2(new_n218), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n785), .A2(new_n268), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G50), .C2(new_n777), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n805), .A2(G143), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G150), .A2(new_n789), .B1(new_n847), .B2(G159), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n778), .A2(new_n842), .B1(new_n780), .B2(new_n810), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G116), .B2(new_n799), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n340), .B(new_n783), .C1(G294), .C2(new_n800), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n807), .C2(new_n772), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G317), .A2(new_n789), .B1(new_n847), .B2(G311), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1097), .A2(new_n1099), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1091), .B1(new_n1106), .B2(new_n765), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n978), .B2(new_n763), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1011), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n707), .B1(new_n1109), .B2(new_n1086), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1011), .B1(new_n750), .B2(new_n1016), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1108), .B1(new_n754), .B2(new_n1109), .C1(new_n1110), .C2(new_n1111), .ZN(G390));
  NAND3_X1  g0912(.A1(new_n745), .A2(new_n688), .A3(new_n833), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n831), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n955), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n944), .A3(new_n929), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n940), .A3(new_n942), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n934), .A2(G330), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n916), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(KEYINPUT92), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n731), .A2(new_n732), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n835), .A4(new_n955), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1116), .A2(new_n1118), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n447), .A2(new_n731), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n964), .A2(new_n661), .A3(new_n1129), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n733), .A2(new_n734), .A3(new_n834), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1131), .A2(new_n955), .B1(new_n1120), .B2(new_n916), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n948), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n955), .B1(new_n731), .B2(new_n835), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n1114), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1125), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1130), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n708), .B1(new_n1128), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1138), .B(KEYINPUT112), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n1128), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n432), .A2(new_n778), .B1(new_n790), .B2(new_n810), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1094), .B(new_n1142), .C1(G68), .C2(new_n1070), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n805), .A2(G294), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n796), .A2(G97), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n340), .B(new_n781), .C1(G116), .C2(new_n847), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(G128), .ZN(new_n1148));
  INV_X1    g0948(.A(G132), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n790), .A2(new_n1148), .B1(new_n1149), .B2(new_n788), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT113), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n780), .A2(new_n326), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n782), .A2(new_n245), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n340), .B1(new_n785), .B2(new_n367), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(G137), .C2(new_n777), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n805), .A2(G125), .B1(new_n796), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1151), .A2(new_n1153), .A3(new_n1156), .A4(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n766), .B1(new_n1147), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n816), .B(new_n1161), .C1(new_n325), .C2(new_n862), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT114), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n943), .B2(new_n761), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1127), .B2(new_n754), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1141), .A2(new_n1166), .ZN(G378));
  AOI21_X1  g0967(.A(new_n713), .B1(new_n929), .B2(new_n930), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n336), .A2(new_n895), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n356), .A2(new_n359), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n356), .B2(new_n359), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR3_X1    g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n867), .B(KEYINPUT40), .C1(new_n939), .C2(new_n917), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT102), .B1(new_n920), .B2(new_n921), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1168), .B(new_n1177), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1177), .B1(new_n923), .B2(new_n1168), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n963), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1168), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1177), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(new_n962), .A3(new_n952), .A4(new_n1180), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1183), .A2(new_n1187), .A3(KEYINPUT57), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1130), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1123), .A2(new_n1124), .A3(new_n835), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1121), .B1(new_n1190), .B2(new_n949), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1137), .B1(new_n1191), .B2(new_n948), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1189), .B1(new_n1127), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n708), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1183), .A2(new_n1187), .A3(KEYINPUT118), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT118), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1130), .B1(new_n1128), .B2(new_n1192), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1195), .B1(new_n1199), .B2(KEYINPUT57), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT118), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n963), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1186), .A2(new_n1180), .B1(new_n962), .B2(new_n952), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1183), .A2(new_n1187), .A3(KEYINPUT118), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n755), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n862), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n756), .B1(G50), .B2(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT117), .Z(new_n1209));
  OAI21_X1  g1009(.A(G33), .B1(new_n377), .B2(new_n378), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G50), .B1(new_n1210), .B2(new_n287), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT115), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n782), .A2(new_n224), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n785), .A2(new_n218), .B1(new_n780), .B2(new_n268), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G116), .C2(new_n789), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G41), .B(new_n397), .C1(G107), .C2(new_n847), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n810), .C2(new_n772), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n777), .A2(G97), .B1(new_n800), .B2(new_n428), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT116), .Z(new_n1219));
  NOR2_X1   g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1212), .B1(new_n1220), .B2(KEYINPUT58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n789), .A2(G125), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n778), .B2(new_n1149), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n847), .A2(G128), .B1(new_n800), .B2(G137), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n780), .B2(new_n1157), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G150), .C2(new_n799), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n805), .A2(G124), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n1070), .C2(G159), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT59), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1229), .B(new_n1230), .C1(new_n1226), .C2(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1221), .B1(KEYINPUT58), .B2(new_n1220), .C1(new_n1228), .C2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1209), .B1(new_n1233), .B2(new_n765), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1177), .B2(new_n761), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1206), .A2(KEYINPUT119), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT119), .B1(new_n1206), .B2(new_n1235), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1200), .B1(new_n1236), .B2(new_n1237), .ZN(G375));
  AOI211_X1 g1038(.A(new_n1018), .B(new_n1140), .C1(new_n1130), .C2(new_n1193), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n754), .B(KEYINPUT120), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT121), .B1(new_n1192), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n756), .B1(G68), .B2(new_n1207), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n955), .A2(new_n761), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n381), .B1(new_n268), .B2(new_n782), .C1(new_n772), .C2(new_n842), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G107), .B2(new_n796), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n799), .A2(new_n428), .B1(new_n847), .B2(G283), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n778), .A2(new_n524), .B1(new_n780), .B2(new_n226), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G294), .B2(new_n789), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n772), .A2(new_n1148), .B1(new_n367), .B2(new_n780), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT123), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n397), .B1(new_n326), .B2(new_n792), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1213), .B(new_n1253), .C1(G50), .C2(new_n799), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(KEYINPUT124), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n777), .A2(new_n1158), .B1(new_n847), .B2(G137), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n1149), .C2(new_n790), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT124), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1250), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1242), .B(new_n1243), .C1(new_n765), .C2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1241), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1192), .A2(KEYINPUT121), .A3(new_n1240), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1239), .A2(new_n1263), .ZN(G381));
  OR2_X1    g1064(.A1(G375), .A2(G378), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  INV_X1    g1067(.A(G384), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OR2_X1    g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(G381), .A2(G387), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(new_n1271), .ZN(G407));
  INV_X1    g1072(.A(G213), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(G343), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1266), .A2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT125), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1267), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(new_n828), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1020), .A2(G390), .A3(new_n1049), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1280), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1200), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1183), .A2(new_n1187), .A3(new_n1240), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1204), .A2(new_n1194), .A3(new_n1205), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1235), .B(new_n1287), .C1(new_n1288), .C2(new_n1018), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n1141), .A3(new_n1166), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1274), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1134), .A2(KEYINPUT60), .A3(new_n1130), .A4(new_n1137), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n707), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1134), .A2(new_n1130), .A3(new_n1137), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT60), .B1(new_n1193), .B2(new_n1130), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1268), .B1(new_n1296), .B2(new_n1263), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1294), .B1(new_n1138), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n707), .A3(new_n1292), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1262), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1301), .A2(new_n1241), .A3(new_n1260), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1302), .A3(G384), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1297), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1274), .A2(G2897), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT126), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1307), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1285), .B1(new_n1291), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1309), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1291), .B2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  AOI211_X1 g1116(.A(new_n1274), .B(new_n1309), .C1(new_n1286), .C2(new_n1290), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1313), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1284), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1314), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1320), .B(new_n1285), .C1(new_n1291), .C2(new_n1311), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1284), .B1(KEYINPUT63), .B2(new_n1317), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1278), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1312), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1291), .A2(new_n1314), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1325), .A2(new_n1328), .A3(new_n1284), .A4(new_n1320), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1326), .A2(KEYINPUT62), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1330), .A2(new_n1312), .A3(new_n1315), .ZN(new_n1331));
  OAI211_X1 g1131(.A(KEYINPUT127), .B(new_n1329), .C1(new_n1331), .C2(new_n1284), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1324), .A2(new_n1332), .ZN(G405));
  XNOR2_X1  g1133(.A(G375), .B(G378), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1314), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1335), .B(new_n1284), .ZN(G402));
endmodule


