//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G13), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(G1), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  OR3_X1    g0047(.A1(new_n247), .A2(KEYINPUT12), .A3(G68), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT12), .B1(new_n247), .B2(G68), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n245), .A2(new_n215), .A3(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n214), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n219), .B1(new_n254), .B2(G20), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n248), .A2(new_n249), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n215), .B2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(KEYINPUT67), .A3(G20), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT11), .B1(new_n265), .B2(new_n252), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT64), .B1(new_n271), .B2(new_n214), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT64), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(G1), .A4(G13), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n272), .A2(G274), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT65), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n281), .A2(new_n283), .A3(G232), .A4(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n281), .A2(new_n283), .A3(G226), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n271), .A2(new_n214), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n278), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(new_n272), .A3(new_n275), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n290), .B1(new_n220), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT13), .B1(new_n280), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT65), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n279), .B(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT13), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n291), .A2(new_n272), .A3(new_n275), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n299));
  AOI22_X1  g0099(.A1(G238), .A2(new_n298), .B1(new_n299), .B2(new_n289), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT14), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(G169), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n294), .A2(G179), .A3(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n303), .B1(new_n302), .B2(G169), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n270), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n294), .A2(G190), .A3(new_n301), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n269), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n294), .B2(new_n301), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT70), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n302), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(new_n269), .A4(new_n309), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT3), .B(G33), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(G222), .A3(new_n285), .ZN(new_n320));
  XOR2_X1   g0120(.A(new_n320), .B(KEYINPUT66), .Z(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n281), .A2(new_n283), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n323), .A2(G223), .B1(G77), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n290), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G226), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n296), .B1(new_n327), .B2(new_n292), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G190), .ZN(new_n330));
  OAI21_X1  g0130(.A(G200), .B1(new_n326), .B2(new_n328), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n263), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n252), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n202), .B1(new_n254), .B2(G20), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n253), .A2(new_n336), .B1(new_n202), .B2(new_n250), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(KEYINPUT9), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT9), .B1(new_n335), .B2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT10), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(KEYINPUT69), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n330), .A2(new_n331), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(KEYINPUT69), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(KEYINPUT69), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n330), .A2(new_n345), .A3(new_n331), .A4(new_n342), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n319), .A2(G232), .A3(new_n285), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n324), .A2(G107), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n348), .B(new_n349), .C1(new_n322), .C2(new_n220), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n289), .B1(G244), .B2(new_n298), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n296), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n263), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n257), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n333), .A2(new_n357), .B1(new_n215), .B2(new_n264), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n252), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n264), .B1(new_n254), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n253), .A2(new_n360), .B1(new_n264), .B2(new_n250), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n351), .A2(new_n296), .A3(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n354), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n352), .B2(G200), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(KEYINPUT68), .ZN(new_n367));
  INV_X1    g0167(.A(G190), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n352), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n366), .B2(KEYINPUT68), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n365), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n329), .A2(new_n363), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n335), .A2(new_n337), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n353), .B1(new_n326), .B2(new_n328), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n318), .A2(new_n347), .A3(new_n371), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n333), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G1), .B2(new_n215), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(new_n253), .B1(new_n250), .B2(new_n333), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G58), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(new_n219), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n201), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n257), .A2(G159), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT73), .B1(new_n257), .B2(G159), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT16), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n282), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT7), .B(new_n215), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n319), .B2(G20), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n324), .A2(KEYINPUT71), .A3(KEYINPUT7), .A4(new_n215), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n401), .A2(KEYINPUT72), .A3(G68), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT72), .B1(new_n401), .B2(G68), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n399), .A2(new_n395), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n389), .B1(new_n405), .B2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n252), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n381), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n319), .A2(G226), .A3(G1698), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n319), .A2(G223), .A3(new_n285), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n289), .B1(new_n298), .B2(G232), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n311), .B1(new_n296), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n296), .A2(new_n414), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n417), .B2(G190), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n353), .B1(new_n296), .B2(new_n414), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n417), .B2(G179), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT18), .B1(new_n409), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(G169), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n363), .B2(new_n416), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n401), .A2(G68), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n401), .A2(KEYINPUT72), .A3(G68), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n407), .B1(new_n432), .B2(new_n392), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n425), .B(new_n427), .C1(new_n433), .C2(new_n381), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n418), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n421), .A2(new_n424), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n376), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n281), .A2(new_n283), .A3(G238), .A4(new_n285), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n281), .A2(new_n283), .A3(G244), .A4(G1698), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G116), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n289), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n277), .A2(G1), .A3(G274), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n222), .B1(new_n277), .B2(G1), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n272), .A2(new_n444), .A3(new_n275), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n368), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(G200), .B2(new_n447), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n251), .A2(new_n214), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n254), .A2(G33), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n247), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G87), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT78), .ZN(new_n455));
  OAI21_X1  g0255(.A(G97), .B1(new_n260), .B2(new_n262), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT19), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT67), .B1(new_n261), .B2(G20), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n259), .A2(new_n215), .A3(G33), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT77), .B1(new_n463), .B2(KEYINPUT19), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n319), .A2(new_n215), .A3(G68), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n215), .B1(new_n287), .B2(new_n458), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(G87), .B2(new_n206), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n459), .A2(new_n464), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n252), .ZN(new_n469));
  INV_X1    g0269(.A(new_n355), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n247), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n455), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g0273(.A(KEYINPUT78), .B(new_n471), .C1(new_n468), .C2(new_n252), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n449), .B(new_n454), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n452), .A2(new_n355), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT79), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n465), .A2(new_n467), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n456), .A2(new_n458), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(KEYINPUT77), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n450), .B1(new_n481), .B2(new_n459), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT78), .B1(new_n482), .B2(new_n471), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n469), .A2(new_n455), .A3(new_n472), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n478), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n447), .A2(G179), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n353), .B2(new_n447), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n475), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n215), .C1(G33), .C2(new_n460), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT20), .ZN(new_n493));
  INV_X1    g0293(.A(G116), .ZN(new_n494));
  AOI22_X1  g0294(.A1(KEYINPUT81), .A2(new_n493), .B1(new_n494), .B2(G20), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n495), .A3(new_n252), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n250), .A2(G116), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n452), .B2(G116), .ZN(new_n500));
  OAI21_X1  g0300(.A(G169), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G41), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n276), .A2(KEYINPUT5), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n254), .A4(G45), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n272), .A3(G270), .A4(new_n275), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n254), .B(G45), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT75), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n503), .A2(KEYINPUT75), .A3(new_n254), .A4(G45), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n510), .A3(new_n504), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n272), .A2(G274), .A3(new_n275), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n281), .A2(new_n283), .A3(G257), .A4(new_n285), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n319), .A2(KEYINPUT80), .A3(G257), .A4(new_n285), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n319), .A2(G264), .A3(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n324), .A2(G303), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n513), .B1(new_n289), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n490), .B1(new_n501), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n500), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n496), .A2(new_n497), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n496), .A2(new_n497), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n521), .A2(new_n526), .A3(G179), .ZN(new_n527));
  INV_X1    g0327(.A(new_n513), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n520), .A2(new_n289), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n530), .A2(new_n526), .A3(KEYINPUT21), .A4(G169), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n522), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n521), .A2(new_n311), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n526), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n530), .A2(new_n368), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n247), .A2(G97), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n453), .B2(G97), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT7), .B1(new_n324), .B2(new_n215), .ZN(new_n541));
  AOI211_X1 g0341(.A(new_n398), .B(G20), .C1(new_n281), .C2(new_n283), .ZN(new_n542));
  OAI21_X1  g0342(.A(G107), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  AND2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n205), .ZN(new_n546));
  INV_X1    g0346(.A(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(KEYINPUT6), .A3(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT74), .B1(new_n551), .B2(new_n252), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT74), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n553), .B(new_n450), .C1(new_n543), .C2(new_n550), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n540), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AND4_X1   g0355(.A1(G257), .A2(new_n505), .A3(new_n272), .A4(new_n275), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n281), .A2(new_n283), .A3(G244), .A4(new_n285), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n319), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n319), .A2(G250), .A3(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n491), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n556), .B1(new_n562), .B2(new_n289), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n511), .A2(new_n512), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n363), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n353), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n555), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n546), .A2(new_n548), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n569), .A2(new_n215), .B1(new_n264), .B2(new_n357), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n547), .B1(new_n399), .B2(new_n395), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n252), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n553), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n252), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n311), .A2(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT76), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n368), .B1(new_n578), .B2(new_n311), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n563), .A2(new_n564), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n575), .A2(new_n577), .A3(new_n540), .A4(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n505), .A2(new_n272), .A3(G264), .A4(new_n275), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n511), .B2(new_n512), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n281), .A2(new_n283), .A3(G250), .A4(new_n285), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n281), .A2(new_n283), .A3(G257), .A4(G1698), .ZN(new_n586));
  INV_X1    g0386(.A(G294), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n586), .C1(new_n261), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n289), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n363), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n589), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n353), .B1(new_n591), .B2(new_n583), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n319), .A2(new_n215), .A3(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n319), .A2(new_n595), .A3(new_n215), .A4(G87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n547), .A2(G20), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT82), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT23), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n215), .A2(G33), .A3(G116), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n598), .B2(KEYINPUT23), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n599), .B1(new_n598), .B2(KEYINPUT23), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT24), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT24), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n597), .A2(new_n608), .A3(new_n605), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n450), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n547), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT25), .B1(new_n250), .B2(new_n547), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(new_n452), .B2(new_n547), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n590), .B(new_n592), .C1(new_n610), .C2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n609), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n608), .B1(new_n597), .B2(new_n605), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n252), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n614), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n584), .A2(new_n589), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(G190), .ZN(new_n621));
  AOI21_X1  g0421(.A(G200), .B1(new_n584), .B2(new_n589), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n618), .B(new_n619), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n568), .A2(new_n581), .A3(new_n615), .A4(new_n623), .ZN(new_n624));
  NOR4_X1   g0424(.A1(new_n438), .A2(new_n489), .A3(new_n538), .A4(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n375), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT17), .B1(new_n409), .B2(new_n418), .ZN(new_n627));
  INV_X1    g0427(.A(new_n435), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n352), .A2(new_n353), .B1(new_n359), .B2(new_n361), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT84), .B1(new_n629), .B2(new_n364), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n365), .A2(KEYINPUT84), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n314), .A2(new_n269), .A3(new_n309), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n627), .B(new_n628), .C1(new_n308), .C2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n424), .A2(new_n434), .A3(KEYINPUT83), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT83), .B1(new_n424), .B2(new_n434), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT85), .ZN(new_n641));
  INV_X1    g0441(.A(new_n344), .ZN(new_n642));
  INV_X1    g0442(.A(new_n346), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n626), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n487), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n592), .A2(new_n590), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n618), .B2(new_n619), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n522), .A2(new_n531), .A3(new_n527), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n475), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n568), .A2(new_n581), .A3(new_n623), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n489), .B2(new_n568), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n483), .A2(new_n484), .B1(G87), .B2(new_n453), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n449), .B1(new_n647), .B2(new_n487), .ZN(new_n658));
  INV_X1    g0458(.A(new_n568), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n654), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n646), .B1(new_n438), .B2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n246), .A2(new_n215), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(G213), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n526), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT87), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n538), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n535), .A2(new_n533), .A3(new_n526), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n651), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n674), .A2(new_n677), .B1(new_n651), .B2(new_n672), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n669), .B1(new_n610), .B2(new_n614), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n615), .A2(new_n623), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n669), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n615), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n663), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n674), .A2(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n672), .A2(new_n651), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND4_X1   g0489(.A1(new_n663), .A2(new_n689), .A3(G330), .A4(new_n684), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n615), .A2(new_n623), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n532), .A2(new_n669), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n650), .A2(new_n683), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n209), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n212), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n660), .A2(new_n656), .ZN(new_n707));
  INV_X1    g0507(.A(new_n654), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n706), .B1(new_n709), .B2(new_n683), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n661), .A2(KEYINPUT29), .A3(new_n669), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AND4_X1   g0513(.A1(new_n615), .A2(new_n568), .A3(new_n581), .A4(new_n623), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n658), .A3(new_n676), .A4(new_n683), .ZN(new_n715));
  NOR2_X1   g0515(.A1(KEYINPUT89), .A2(KEYINPUT30), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n443), .A2(new_n446), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n563), .A2(new_n717), .A3(new_n589), .A4(new_n584), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n528), .A2(new_n529), .A3(G179), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n528), .A2(new_n529), .A3(G179), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n591), .A2(new_n447), .A3(new_n583), .ZN(new_n722));
  INV_X1    g0522(.A(new_n716), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n563), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n717), .A2(G179), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n566), .A3(new_n530), .A4(new_n620), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n720), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n727), .B2(new_n669), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n715), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n711), .A2(new_n713), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n705), .B1(new_n734), .B2(G1), .ZN(G364));
  NAND2_X1  g0535(.A1(new_n678), .A2(new_n679), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT90), .Z(new_n737));
  NAND2_X1  g0537(.A1(new_n689), .A2(G330), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n245), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n254), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n700), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n737), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n214), .B1(G20), .B2(new_n353), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n215), .A2(new_n363), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(new_n311), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n215), .A2(G179), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G190), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n748), .A2(G322), .B1(new_n752), .B2(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(new_n750), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n753), .B(new_n324), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n746), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G190), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n749), .A2(new_n368), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(G283), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n368), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n215), .ZN(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n762), .B1(new_n587), .B2(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n757), .A2(new_n368), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n756), .B(new_n767), .C1(G326), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n760), .A2(new_n547), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n764), .A2(new_n460), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(G68), .C2(new_n758), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n751), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n319), .B1(new_n747), .B2(new_n382), .ZN(new_n778));
  INV_X1    g0578(.A(new_n755), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G77), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n766), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n768), .A2(G50), .B1(new_n781), .B2(G87), .ZN(new_n782));
  AND4_X1   g0582(.A1(new_n774), .A2(new_n777), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n745), .B1(new_n771), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n742), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n243), .A2(G45), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT91), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n699), .A2(new_n319), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(G45), .C2(new_n212), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n319), .A2(new_n209), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(G116), .B2(new_n209), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT92), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n745), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT93), .Z(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n792), .B2(KEYINPUT92), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n785), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n796), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n689), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n744), .A2(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n362), .A2(new_n669), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n629), .A2(KEYINPUT84), .A3(new_n364), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n630), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n371), .B2(new_n805), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n709), .B2(new_n683), .ZN(new_n810));
  INV_X1    g0610(.A(new_n371), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n669), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n709), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n732), .ZN(new_n814));
  OR3_X1    g0614(.A1(new_n813), .A2(KEYINPUT96), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT96), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n742), .B1(new_n813), .B2(new_n814), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n745), .A2(new_n794), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n743), .B1(new_n264), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n745), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n748), .A2(G143), .B1(new_n779), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(new_n768), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  INV_X1    g0625(.A(new_n758), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n760), .A2(new_n219), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n319), .B1(new_n751), .B2(new_n832), .C1(new_n764), .C2(new_n382), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(G50), .C2(new_n781), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n829), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n324), .B1(new_n766), .B2(new_n547), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT95), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n755), .A2(new_n494), .B1(new_n751), .B2(new_n754), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G294), .B2(new_n748), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n773), .B1(G283), .B2(new_n758), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n768), .A2(G303), .B1(new_n761), .B2(G87), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n837), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n820), .B1(new_n821), .B2(new_n843), .C1(new_n809), .C2(new_n795), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n818), .A2(new_n844), .ZN(G384));
  OR2_X1    g0645(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(G116), .A3(new_n216), .A4(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT36), .Z(new_n849));
  OAI211_X1 g0649(.A(new_n213), .B(G77), .C1(new_n382), .C2(new_n219), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n202), .A2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n254), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n739), .A2(new_n254), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n450), .B1(new_n432), .B2(new_n392), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n390), .B1(new_n402), .B2(new_n403), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT16), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n381), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n419), .B1(new_n859), .B2(new_n423), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n667), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n409), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n427), .ZN(new_n864));
  INV_X1    g0664(.A(new_n667), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n419), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n862), .A2(new_n868), .B1(new_n436), .B2(new_n861), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n709), .A2(new_n812), .B1(new_n365), .B2(new_n683), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n270), .A2(new_n669), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n306), .A2(new_n307), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n317), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n633), .A2(new_n872), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n280), .A2(new_n293), .A3(KEYINPUT13), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n297), .B1(new_n296), .B2(new_n300), .ZN(new_n877));
  OAI21_X1  g0677(.A(G169), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT14), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n305), .A3(new_n304), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n875), .B1(new_n880), .B2(new_n270), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT97), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n308), .A2(new_n633), .A3(new_n872), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT97), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n313), .B2(new_n316), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n883), .B(new_n884), .C1(new_n885), .C2(new_n872), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n871), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n870), .A2(new_n888), .B1(new_n638), .B2(new_n667), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT98), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  AOI221_X4 g0691(.A(new_n891), .B1(new_n436), .B2(new_n861), .C1(new_n862), .C2(new_n868), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n862), .A2(new_n868), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n436), .A2(new_n861), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT39), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n894), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n628), .A2(new_n627), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n636), .B2(new_n637), .ZN(new_n900));
  INV_X1    g0700(.A(new_n866), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n864), .A2(new_n866), .A3(new_n419), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n900), .A2(new_n901), .B1(new_n868), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n897), .B(new_n898), .C1(new_n904), .C2(KEYINPUT38), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n308), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n683), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n889), .B(new_n890), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n908), .B1(new_n896), .B2(new_n905), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n638), .A2(new_n667), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n892), .A2(new_n895), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n882), .A2(new_n886), .ZN(new_n913));
  INV_X1    g0713(.A(new_n812), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n629), .A2(new_n364), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n661), .A2(new_n914), .B1(new_n915), .B2(new_n669), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n911), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT98), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n437), .B1(new_n710), .B2(new_n712), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n921), .A2(new_n646), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n920), .B(new_n922), .Z(new_n923));
  OAI21_X1  g0723(.A(new_n898), .B1(new_n904), .B2(KEYINPUT38), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n808), .B1(new_n715), .B2(new_n730), .ZN(new_n925));
  AND4_X1   g0725(.A1(KEYINPUT40), .A2(new_n925), .A3(new_n882), .A4(new_n886), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT99), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(new_n926), .A3(KEYINPUT99), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n913), .B(new_n925), .C1(new_n892), .C2(new_n895), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n437), .A2(new_n731), .ZN(new_n936));
  OAI21_X1  g0736(.A(G330), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n854), .B1(new_n923), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT100), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n939), .A2(new_n940), .B1(new_n938), .B2(new_n923), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n853), .B1(new_n941), .B2(new_n942), .ZN(G367));
  AND2_X1   g0743(.A1(new_n568), .A2(new_n581), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n555), .A2(new_n669), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(new_n650), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n669), .B1(new_n946), .B2(new_n568), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n659), .A2(new_n669), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n693), .A3(new_n694), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n947), .B1(new_n951), .B2(KEYINPUT42), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT42), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n950), .A2(new_n953), .A3(new_n693), .A4(new_n694), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n657), .A2(new_n683), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n647), .A3(new_n487), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n489), .B2(new_n956), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n952), .A2(new_n960), .A3(new_n959), .A4(new_n954), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT101), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n686), .A2(new_n691), .A3(new_n966), .A4(new_n950), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n685), .A2(new_n690), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n969), .B2(new_n950), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n700), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n697), .B2(new_n950), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n695), .A2(new_n696), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n975), .A2(KEYINPUT44), .A3(new_n948), .A4(new_n949), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT102), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT102), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n973), .C1(new_n697), .C2(new_n950), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n697), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT45), .B1(new_n697), .B2(new_n950), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT103), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n692), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n684), .A2(new_n694), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n695), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT104), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n689), .B2(G330), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n678), .A2(KEYINPUT104), .A3(new_n679), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n695), .B(new_n986), .C1(new_n680), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n733), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n977), .B(new_n980), .C1(new_n982), .C2(new_n981), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n969), .A3(KEYINPUT103), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n985), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n972), .B1(new_n997), .B2(new_n734), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n971), .B1(new_n998), .B2(new_n741), .ZN(new_n999));
  INV_X1    g0799(.A(new_n788), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n236), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n798), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n209), .B2(new_n355), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G50), .A2(new_n779), .B1(new_n752), .B2(G137), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1004), .B(new_n319), .C1(new_n825), .C2(new_n747), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n758), .A2(G159), .B1(new_n761), .B2(G77), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n382), .B2(new_n766), .C1(new_n219), .C2(new_n764), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(G143), .C2(new_n770), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G283), .A2(new_n779), .B1(new_n752), .B2(G317), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n319), .B1(new_n748), .B2(G303), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT46), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n766), .B2(new_n494), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n764), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G107), .A2(new_n1015), .B1(new_n758), .B2(G294), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n460), .B2(new_n760), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1014), .B(new_n1017), .C1(G311), .C2(new_n770), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1008), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT47), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n742), .B1(new_n1001), .B2(new_n1003), .C1(new_n1020), .C2(new_n821), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT105), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n801), .B2(new_n958), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n999), .A2(new_n1023), .ZN(G387));
  NOR2_X1   g0824(.A1(new_n994), .A2(new_n701), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT109), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n993), .A2(new_n733), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n993), .A2(new_n733), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(KEYINPUT109), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n702), .A2(new_n791), .B1(G107), .B2(new_n209), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n233), .A2(new_n277), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n702), .ZN(new_n1033));
  AOI211_X1 g0833(.A(G45), .B(new_n1033), .C1(G68), .C2(G77), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n333), .A2(G50), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1000), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1031), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n742), .B1(new_n1038), .B2(new_n798), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n684), .A2(new_n801), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n766), .A2(new_n264), .B1(new_n751), .B2(new_n825), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT107), .Z(new_n1042));
  OAI21_X1  g0842(.A(new_n319), .B1(new_n755), .B2(new_n219), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G50), .B2(new_n748), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n768), .A2(G159), .B1(new_n761), .B2(G97), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n764), .A2(new_n355), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n377), .B2(new_n758), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n748), .A2(G317), .B1(new_n779), .B2(G303), .ZN(new_n1049));
  INV_X1    g0849(.A(G322), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1049), .B1(new_n754), .B2(new_n826), .C1(new_n769), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(G283), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n764), .A2(new_n1054), .B1(new_n766), .B2(new_n587), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n319), .B1(new_n752), .B2(G326), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n494), .C2(new_n760), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1057), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1048), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1039), .B(new_n1040), .C1(new_n745), .C2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT106), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n993), .B2(new_n740), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n991), .A2(new_n992), .A3(KEYINPUT106), .A4(new_n741), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1030), .A2(new_n1067), .ZN(G393));
  XNOR2_X1  g0868(.A(new_n692), .B(new_n995), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n997), .B(new_n700), .C1(new_n1069), .C2(new_n994), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n948), .A2(new_n796), .A3(new_n949), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n324), .B1(new_n752), .B2(G143), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n219), .B2(new_n766), .C1(new_n221), .C2(new_n760), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT110), .Z(new_n1074));
  OAI22_X1  g0874(.A1(new_n823), .A2(new_n825), .B1(new_n775), .B2(new_n747), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n758), .A2(G50), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n764), .A2(new_n264), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n377), .B2(new_n779), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1015), .A2(G116), .B1(new_n779), .B2(G294), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n765), .B2(new_n826), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT111), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G317), .A2(new_n768), .B1(new_n748), .B2(G311), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n324), .B1(new_n751), .B2(new_n1050), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n772), .B(new_n1086), .C1(G283), .C2(new_n781), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n821), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n240), .A2(new_n788), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n798), .B1(G97), .B2(new_n699), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n743), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1069), .A2(new_n741), .B1(new_n1071), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1070), .A2(new_n1093), .ZN(G390));
  NOR4_X1   g0894(.A1(new_n624), .A2(new_n489), .A3(new_n538), .A4(new_n669), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n729), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(G330), .B(new_n809), .C1(new_n1095), .C2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n887), .A2(new_n1099), .A3(KEYINPUT112), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n908), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n913), .B2(new_n916), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1100), .B1(new_n1102), .B2(new_n924), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT112), .B1(new_n887), .B2(new_n1099), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n908), .B1(new_n871), .B2(new_n887), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n896), .A3(new_n905), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n871), .A2(new_n887), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1099), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1110), .A2(new_n917), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n437), .A2(new_n814), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n921), .A2(new_n646), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1111), .B1(new_n1110), .B2(new_n917), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n700), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n741), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n906), .A2(new_n794), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n743), .B1(new_n333), .B2(new_n819), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n826), .A2(new_n547), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1078), .B(new_n1124), .C1(G283), .C2(new_n768), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G97), .A2(new_n779), .B1(new_n752), .B2(G294), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n324), .C1(new_n494), .C2(new_n747), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n831), .B(new_n1127), .C1(G87), .C2(new_n781), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G159), .A2(new_n1015), .B1(new_n768), .B2(G128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n202), .B2(new_n760), .C1(new_n824), .C2(new_n826), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n319), .B1(new_n751), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n747), .A2(new_n832), .B1(new_n755), .B2(new_n1133), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1130), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n766), .A2(new_n825), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1125), .A2(new_n1128), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1122), .B(new_n1123), .C1(new_n821), .C2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1120), .A2(new_n1121), .A3(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(new_n1114), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1119), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n679), .B1(new_n932), .B2(new_n933), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n373), .A2(new_n865), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT55), .Z(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n645), .B2(new_n375), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n626), .B(new_n1147), .C1(new_n640), .C2(new_n644), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n347), .A2(KEYINPUT85), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n642), .A2(new_n643), .A3(new_n641), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n375), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1147), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n645), .A2(new_n375), .A3(new_n1148), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1144), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT99), .B1(new_n924), .B2(new_n926), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n924), .A2(KEYINPUT99), .A3(new_n926), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1143), .B(new_n1158), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1158), .B1(new_n931), .B2(new_n1143), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n920), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1143), .B1(new_n1160), .B2(new_n1159), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1158), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1167), .A2(new_n909), .A3(new_n919), .A4(new_n1161), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1142), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1142), .A2(new_n1164), .A3(KEYINPUT57), .A4(new_n1168), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n700), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1164), .A2(new_n741), .A3(new_n1168), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n743), .B1(new_n202), .B2(new_n819), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1131), .A2(new_n823), .B1(new_n826), .B2(new_n832), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n748), .A2(G128), .B1(new_n779), .B2(G137), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n766), .B2(new_n1133), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(G150), .C2(new_n1015), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G33), .A2(G41), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT113), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n760), .A2(new_n775), .ZN(new_n1185));
  XOR2_X1   g0985(.A(KEYINPUT115), .B(G124), .Z(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1185), .C1(new_n752), .C2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1181), .A2(new_n1182), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n760), .A2(new_n382), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n826), .A2(new_n460), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G116), .C2(new_n768), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G41), .B(new_n319), .C1(new_n752), .C2(G283), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n748), .A2(G107), .B1(new_n779), .B2(new_n470), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1015), .A2(G68), .B1(new_n781), .B2(G77), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT58), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1184), .B(new_n202), .C1(G41), .C2(new_n319), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT114), .Z(new_n1200));
  AND4_X1   g1000(.A1(new_n1188), .A2(new_n1197), .A3(new_n1198), .A4(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1175), .B1(new_n821), .B2(new_n1201), .C1(new_n1158), .C2(new_n795), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1174), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1173), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT117), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(G375));
  NOR2_X1   g1007(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(new_n1141), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n972), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n1117), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n743), .B1(new_n219), .B2(new_n819), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n319), .B1(new_n752), .B2(G303), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n547), .B2(new_n755), .C1(new_n1054), .C2(new_n747), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1046), .B(new_n1215), .C1(G77), .C2(new_n761), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n494), .A2(new_n826), .B1(new_n823), .B2(new_n587), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G97), .B2(new_n781), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n764), .A2(new_n202), .B1(new_n766), .B2(new_n775), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n768), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n324), .B1(new_n752), .B2(G128), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n824), .B2(new_n747), .C1(new_n825), .C2(new_n755), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n826), .A2(new_n1133), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1222), .A2(new_n1189), .A3(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1216), .A2(new_n1218), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1213), .B1(new_n821), .B2(new_n1225), .C1(new_n913), .C2(new_n795), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1208), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n740), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1212), .A2(new_n1229), .ZN(G381));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  OR2_X1    g1031(.A1(G390), .A2(G384), .ZN(new_n1232));
  INV_X1    g1032(.A(G396), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1030), .A2(new_n1233), .A3(new_n1067), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1232), .A2(G387), .A3(G381), .A4(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1206), .A2(new_n1231), .A3(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n1206), .A2(new_n1231), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(new_n1237), .C2(G343), .ZN(G409));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n999), .A2(new_n1023), .A3(G390), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT123), .ZN(new_n1241));
  INV_X1    g1041(.A(G390), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1233), .B1(new_n1030), .B2(new_n1067), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1234), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT123), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n999), .A2(G390), .A3(new_n1247), .A4(new_n1023), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1241), .A2(new_n1243), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT122), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1234), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n1244), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1245), .A2(KEYINPUT122), .A3(new_n1234), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n999), .A2(new_n1023), .A3(G390), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G390), .B1(new_n999), .B2(new_n1023), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1252), .B(new_n1253), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1249), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1239), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n1249), .C2(new_n1256), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n668), .A2(G213), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1174), .A2(KEYINPUT119), .A3(new_n1202), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT119), .B1(new_n1174), .B2(new_n1202), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1142), .A2(new_n1164), .A3(new_n1211), .A4(new_n1168), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT118), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G378), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1173), .A2(G378), .A3(new_n1204), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1262), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1227), .A2(KEYINPUT60), .A3(new_n1114), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n700), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1209), .B1(new_n1117), .B2(KEYINPUT60), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1229), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(G384), .A2(KEYINPUT120), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G384), .A2(KEYINPUT120), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1275), .B(new_n1229), .C1(new_n1273), .C2(new_n1272), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n668), .A2(G213), .A3(G2897), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1280), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1270), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT121), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1261), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT119), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1203), .A2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(KEYINPUT118), .A3(new_n1211), .A4(new_n1142), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1174), .A2(KEYINPUT119), .A3(new_n1202), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT118), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1266), .A2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1231), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1173), .A2(G378), .A3(new_n1204), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1284), .B1(new_n1299), .B2(new_n1262), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1262), .B(new_n1301), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1300), .A2(KEYINPUT121), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1288), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1302), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1299), .A2(new_n1309), .A3(new_n1262), .A4(new_n1301), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1308), .A2(new_n1286), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1257), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1306), .A2(new_n1314), .ZN(G405));
  NAND2_X1  g1115(.A1(new_n1205), .A2(G378), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1237), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1301), .A2(new_n1318), .ZN(new_n1319));
  XOR2_X1   g1119(.A(new_n1257), .B(new_n1319), .Z(new_n1320));
  XNOR2_X1  g1120(.A(new_n1317), .B(new_n1320), .ZN(G402));
endmodule


