//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT69), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n462), .B1(new_n476), .B2(new_n458), .ZN(G160));
  NOR2_X1   g052(.A1(new_n474), .A2(new_n458), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(G162));
  NAND4_X1  g060(.A1(new_n472), .A2(G138), .A3(new_n458), .A4(new_n473), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n459), .A2(new_n490), .A3(G138), .A4(new_n458), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n458), .A2(G102), .A3(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n474), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n494), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT74), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G651), .B1(G50), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT72), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n517), .B(new_n508), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n507), .A2(KEYINPUT73), .A3(new_n508), .A4(new_n517), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n522), .A2(G89), .A3(new_n523), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n513), .A2(KEYINPUT75), .A3(new_n514), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n532));
  AND2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(KEYINPUT6), .A2(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n531), .A2(new_n535), .A3(G51), .A4(G543), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n507), .A2(G63), .A3(G651), .A4(new_n508), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n528), .A2(new_n530), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G168));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n509), .A2(G64), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n522), .A2(G90), .A3(new_n523), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n531), .A2(new_n535), .A3(G543), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT76), .B(G52), .Z(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n545), .A2(KEYINPUT77), .A3(new_n548), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n544), .B1(new_n551), .B2(new_n552), .ZN(G171));
  AND2_X1   g128(.A1(new_n524), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n546), .A2(G43), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n541), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n546), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n524), .A2(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n541), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n551), .A2(new_n552), .ZN(new_n572));
  INV_X1    g147(.A(new_n544), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n545), .A2(KEYINPUT77), .A3(new_n548), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT77), .B1(new_n545), .B2(new_n548), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n571), .B(new_n573), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G301));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n539), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n528), .A2(KEYINPUT79), .A3(new_n538), .A4(new_n530), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G286));
  OAI21_X1  g159(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n546), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(G87), .B2(new_n524), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n524), .A2(G86), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT81), .Z(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n510), .A2(KEYINPUT80), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT80), .B1(new_n510), .B2(new_n592), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G48), .B2(new_n515), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n591), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n510), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G47), .B2(new_n546), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n524), .A2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n522), .A2(new_n523), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n546), .B(KEYINPUT82), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n606), .A2(new_n610), .B1(G54), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n614), .A2(G651), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT84), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n605), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n605), .B1(new_n621), .B2(G868), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  XNOR2_X1  g199(.A(G299), .B(KEYINPUT85), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  INV_X1    g204(.A(new_n558), .ZN(new_n630));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(G559), .B1(new_n618), .B2(new_n620), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g210(.A1(new_n468), .A2(new_n458), .A3(new_n459), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2100), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n478), .A2(G123), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n480), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(new_n458), .B2(G111), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT15), .B(G2435), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n652), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT86), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT17), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT87), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n661), .A3(new_n662), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  INV_X1    g245(.A(new_n663), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n661), .A3(new_n664), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n682), .B1(KEYINPUT20), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(KEYINPUT20), .C2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1991), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n689), .B(new_n694), .ZN(G229));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G27), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G164), .B2(new_n696), .ZN(new_n698));
  MUX2_X1   g273(.A(new_n697), .B(new_n698), .S(KEYINPUT100), .Z(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT101), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G2078), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n480), .A2(G139), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  AOI22_X1  g279(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n702), .B(new_n704), .C1(new_n458), .C2(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G33), .B(new_n706), .S(G29), .Z(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G2072), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(G2072), .ZN(new_n709));
  INV_X1    g284(.A(G28), .ZN(new_n710));
  AOI21_X1  g285(.A(G29), .B1(new_n710), .B2(KEYINPUT30), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(KEYINPUT30), .B2(new_n710), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n644), .B2(new_n696), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n708), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G29), .A2(G32), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n480), .A2(G141), .ZN(new_n716));
  INV_X1    g291(.A(G129), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n472), .A2(new_n473), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G2105), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n468), .A2(G105), .A3(new_n458), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(KEYINPUT98), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT99), .Z(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT26), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT26), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(KEYINPUT98), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n720), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n715), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT31), .B(G11), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n714), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G162), .A2(new_n696), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n696), .B2(G35), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n738), .A2(G2090), .A3(new_n739), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n734), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(new_n696), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G160), .B2(new_n696), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n696), .A2(G26), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT96), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n458), .A2(G116), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G104), .C2(G2105), .ZN(new_n756));
  AND3_X1   g331(.A1(new_n718), .A2(G140), .A3(new_n458), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n478), .A2(KEYINPUT95), .A3(G128), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(KEYINPUT95), .B1(new_n478), .B2(G128), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n756), .B(new_n758), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n754), .B1(new_n762), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G16), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G19), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n558), .B2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1341), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n766), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1966), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n765), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n744), .A2(new_n751), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n621), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT94), .B1(G4), .B2(G16), .ZN(new_n776));
  OR3_X1    g351(.A1(KEYINPUT94), .A2(G4), .A3(G16), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n766), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n766), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n766), .A2(G20), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n787));
  OAI211_X1 g362(.A(KEYINPUT23), .B(new_n786), .C1(new_n787), .C2(new_n766), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT23), .B2(new_n786), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n774), .A2(new_n781), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n766), .A2(G22), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G166), .B2(new_n766), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G1971), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(G1971), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n766), .A2(G6), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G305), .B2(G16), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  AOI211_X1 g373(.A(new_n794), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n766), .A2(G23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n588), .B2(new_n766), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT33), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1976), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n799), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n799), .A2(KEYINPUT93), .A3(new_n800), .A4(new_n804), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n766), .A2(G24), .ZN(new_n811));
  INV_X1    g386(.A(G290), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n766), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT91), .B(G1986), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G25), .A2(G29), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n478), .A2(G119), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n480), .A2(G131), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(G29), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT90), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT35), .B(G1991), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n807), .A2(new_n808), .ZN(new_n828));
  INV_X1    g403(.A(new_n809), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n816), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n816), .A2(new_n833), .A3(new_n827), .A4(new_n830), .ZN(new_n834));
  AOI211_X1 g409(.A(new_n701), .B(new_n791), .C1(new_n832), .C2(new_n834), .ZN(G311));
  AOI21_X1  g410(.A(new_n791), .B1(new_n832), .B2(new_n834), .ZN(new_n836));
  INV_X1    g411(.A(new_n701), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(G150));
  AOI22_X1  g413(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n541), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n522), .A2(G93), .A3(new_n523), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n546), .A2(G55), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n841), .A2(KEYINPUT102), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT102), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n621), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g427(.A(KEYINPUT103), .B(new_n840), .C1(new_n843), .C2(new_n844), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n558), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n630), .A2(new_n851), .A3(new_n845), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n850), .B(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n847), .B1(new_n858), .B2(G860), .ZN(G145));
  NAND2_X1  g434(.A1(new_n478), .A2(G130), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n480), .A2(G142), .ZN(new_n861));
  NOR2_X1   g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(new_n458), .B2(G118), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n860), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G162), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n644), .B(G160), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n865), .B(new_n866), .Z(new_n867));
  INV_X1    g442(.A(new_n756), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n869));
  INV_X1    g444(.A(G128), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n719), .B2(new_n870), .ZN(new_n871));
  AOI211_X1 g446(.A(new_n868), .B(new_n757), .C1(new_n871), .C2(new_n759), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n493), .A2(new_n498), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(G164), .A2(new_n762), .ZN(new_n875));
  INV_X1    g450(.A(new_n729), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n877), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n874), .A2(new_n875), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n729), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n637), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n884), .B(new_n885), .C1(new_n880), .C2(new_n879), .ZN(new_n888));
  INV_X1    g463(.A(new_n637), .ZN(new_n889));
  OAI22_X1  g464(.A1(new_n877), .A2(new_n878), .B1(KEYINPUT104), .B2(new_n706), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n823), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n823), .B1(new_n887), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n867), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n887), .A2(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n822), .ZN(new_n898));
  INV_X1    g473(.A(new_n867), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n892), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  XNOR2_X1  g478(.A(G288), .B(G303), .ZN(new_n904));
  XNOR2_X1  g479(.A(G290), .B(KEYINPUT106), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(G305), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n787), .A2(new_n612), .A3(new_n616), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n787), .B1(new_n616), .B2(new_n612), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n617), .A2(G299), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n909), .A3(KEYINPUT41), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n633), .A2(new_n856), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n633), .A2(new_n856), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n910), .A2(new_n911), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n916), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n922), .A3(KEYINPUT105), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n915), .B(new_n925), .C1(new_n917), .C2(new_n918), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n923), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n907), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  INV_X1    g506(.A(new_n907), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n927), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G868), .ZN(new_n935));
  INV_X1    g510(.A(new_n845), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(G868), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n903), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n631), .B1(new_n930), .B2(new_n933), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n940), .A2(KEYINPUT107), .A3(new_n937), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(G295));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n935), .A2(new_n943), .A3(new_n938), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT108), .B1(new_n940), .B2(new_n937), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(G331));
  AND2_X1   g521(.A1(new_n582), .A2(new_n583), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT109), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  NAND3_X1  g525(.A1(G171), .A2(new_n950), .A3(G286), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(G168), .B1(new_n574), .B2(new_n578), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n952), .A2(KEYINPUT110), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT110), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n857), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  AND3_X1   g533(.A1(G171), .A2(new_n950), .A3(G286), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n950), .B1(G171), .B2(G286), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n948), .A2(KEYINPUT78), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n539), .B1(new_n962), .B2(new_n577), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n958), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(KEYINPUT110), .A3(new_n953), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n856), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n956), .A2(new_n957), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n964), .A2(KEYINPUT111), .A3(new_n856), .A4(new_n965), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n915), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n956), .A2(new_n921), .A3(new_n966), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n907), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n896), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n907), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n921), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n967), .B2(new_n968), .ZN(new_n976));
  INV_X1    g551(.A(new_n915), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n956), .B2(new_n966), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n932), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n896), .A4(new_n971), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n972), .B2(new_n973), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n896), .A3(new_n971), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  MUX2_X1   g560(.A(new_n982), .B(new_n985), .S(KEYINPUT44), .Z(G397));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n873), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  AND2_X1   g564(.A1(G160), .A2(G40), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(G1996), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT114), .B1(new_n994), .B2(G1996), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n876), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n762), .A2(G2067), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n872), .A2(new_n764), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n1000), .B(new_n1001), .C1(G1996), .C2(new_n876), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n822), .A2(new_n826), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n999), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT126), .B1(new_n1006), .B2(new_n1000), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1000), .ZN(new_n1009));
  INV_X1    g584(.A(new_n998), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n994), .A2(KEYINPUT114), .A3(G1996), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n729), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n994), .B2(new_n1002), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1008), .B(new_n1009), .C1(new_n1013), .C2(new_n1005), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n994), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1001), .A2(new_n1000), .A3(new_n876), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n994), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n997), .A2(KEYINPUT46), .A3(new_n998), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT47), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n822), .A2(new_n826), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n994), .B1(new_n1005), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G290), .A2(G1986), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT113), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n992), .A2(new_n1026), .A3(new_n993), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT48), .Z(new_n1028));
  NOR3_X1   g603(.A1(new_n1013), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1015), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n493), .B2(new_n498), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(KEYINPUT117), .A3(new_n750), .A4(new_n990), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n750), .A3(new_n990), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n988), .A2(new_n989), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1032), .A2(KEYINPUT45), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n990), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1034), .A2(new_n1040), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1031), .B1(new_n1046), .B2(new_n539), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1034), .A2(new_n1040), .A3(G168), .A4(new_n1045), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1031), .B1(new_n1048), .B2(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT62), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(KEYINPUT124), .A2(KEYINPUT53), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1054));
  AND3_X1   g629(.A1(new_n1041), .A2(new_n990), .A3(new_n1042), .ZN(new_n1055));
  INV_X1    g630(.A(G2078), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  MUX2_X1   g632(.A(new_n1053), .B(new_n1054), .S(new_n1057), .Z(new_n1058));
  AND3_X1   g633(.A1(new_n1035), .A2(new_n990), .A3(new_n1037), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G1961), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G301), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1049), .A2(KEYINPUT51), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(new_n1064), .C1(new_n1049), .C2(new_n1047), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n597), .A2(new_n590), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G1981), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(G305), .B2(G1981), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1032), .A2(new_n990), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1067), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n588), .A2(G1976), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1071), .A2(new_n1075), .A3(G8), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n588), .A2(G1976), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1071), .A2(G8), .A3(new_n1076), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1075), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1074), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1035), .A2(new_n990), .A3(new_n1037), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1055), .A2(G1971), .B1(G2090), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G303), .A2(G8), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n1090), .B(KEYINPUT55), .Z(new_n1091));
  AND3_X1   g666(.A1(new_n1089), .A2(G8), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1089), .B2(G8), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1087), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1052), .A2(new_n1062), .A3(new_n1065), .A4(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1074), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1046), .A2(G8), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1096), .A2(new_n947), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(KEYINPUT63), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1976), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1074), .A2(new_n1103), .A3(new_n588), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(G1981), .B2(G305), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1099), .A2(new_n1102), .B1(new_n1072), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1097), .A2(new_n1092), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1094), .A2(new_n947), .A3(new_n1101), .A4(new_n1098), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1095), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1060), .A2(KEYINPUT125), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1060), .A2(KEYINPUT125), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1057), .A2(KEYINPUT124), .A3(KEYINPUT53), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1057), .A2(new_n1054), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n1111), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1058), .A2(G301), .A3(new_n1061), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT54), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1094), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1088), .A2(new_n779), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1032), .A2(new_n1120), .A3(new_n990), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1032), .B2(new_n990), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1119), .B1(new_n1123), .B2(G2067), .ZN(new_n1124));
  INV_X1    g699(.A(G1956), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1088), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n787), .A2(KEYINPUT119), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(KEYINPUT119), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1127), .A2(KEYINPUT119), .ZN(new_n1130));
  NAND3_X1  g705(.A1(G299), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1041), .A2(new_n990), .A3(new_n1042), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1126), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n617), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1124), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1956), .B1(new_n1033), .B2(new_n990), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1135), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1132), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(G1341), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1041), .A2(new_n1145), .A3(new_n990), .A4(new_n1042), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n630), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1148), .ZN(new_n1150));
  AOI211_X1 g725(.A(new_n630), .B(new_n1150), .C1(new_n1144), .C2(new_n1146), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1126), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1133), .B1(new_n1126), .B2(new_n1135), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n1157));
  AOI21_X1  g732(.A(G1348), .B1(new_n1033), .B2(new_n990), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1121), .A2(new_n1122), .A3(G2067), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1119), .B(KEYINPUT60), .C1(new_n1123), .C2(G2067), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n1161), .A3(new_n1137), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1152), .A2(new_n1156), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1161), .A2(new_n1137), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1138), .B(new_n1141), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1147), .B(new_n1148), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT61), .B1(new_n1141), .B2(new_n1136), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1165), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(KEYINPUT123), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1118), .B1(new_n1168), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1114), .A2(new_n579), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(new_n1062), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1109), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1013), .A2(new_n1024), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1026), .B1(G1986), .B2(G290), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1183), .B1(new_n994), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1030), .B1(new_n1182), .B2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g761(.A(G319), .ZN(new_n1188));
  NOR4_X1   g762(.A1(G229), .A2(new_n1188), .A3(G401), .A4(G227), .ZN(new_n1189));
  AND2_X1   g763(.A1(new_n901), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n982), .A2(new_n1190), .ZN(G225));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g766(.A1(G225), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n982), .A2(new_n1190), .A3(KEYINPUT127), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1194), .ZN(G308));
endmodule


