//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n453), .A2(G567), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n464), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G137), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT70), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT68), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(G2104), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(new_n468), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n476), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(G113), .A2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n463), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G101), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n475), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(G160));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n470), .A2(G136), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT72), .Z(new_n494));
  AND4_X1   g069(.A1(G2105), .A2(new_n464), .A3(new_n468), .A4(new_n466), .ZN(new_n495));
  AOI211_X1 g070(.A(new_n492), .B(new_n494), .C1(G124), .C2(new_n495), .ZN(G162));
  NAND2_X1  g071(.A1(new_n479), .A2(new_n482), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n464), .A2(new_n466), .A3(new_n500), .A4(new_n468), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n497), .A2(new_n499), .B1(KEYINPUT4), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(G114), .B2(new_n467), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n464), .A2(new_n466), .A3(G2105), .A4(new_n468), .ZN(new_n506));
  INV_X1    g081(.A(G126), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n502), .A2(KEYINPUT73), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n480), .A2(new_n468), .A3(new_n481), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n481), .B1(new_n480), .B2(new_n468), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n499), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G114), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n503), .B1(new_n516), .B2(G2105), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n495), .B2(G126), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n510), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n509), .A2(new_n519), .ZN(G164));
  OR2_X1    g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n526), .A2(new_n535), .ZN(G166));
  NAND3_X1  g111(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT74), .Z(new_n538));
  NAND2_X1  g113(.A1(new_n530), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n539), .B(new_n541), .C1(new_n533), .C2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n525), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n530), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n533), .B2(new_n548), .ZN(new_n549));
  OR3_X1    g124(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT75), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT75), .B1(new_n546), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n525), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n530), .A2(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n533), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n530), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n521), .A2(new_n522), .B1(new_n528), .B2(new_n529), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n565), .B(new_n567), .C1(new_n525), .C2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND2_X1  g147(.A1(new_n530), .A2(G49), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n533), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT76), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n579), .B(G651), .C1(new_n523), .C2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n530), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n533), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n521), .B2(new_n522), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g166(.A(KEYINPUT77), .B(G651), .C1(new_n587), .C2(new_n588), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n585), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n525), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n530), .A2(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n533), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n566), .A2(G92), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT10), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n523), .A2(G66), .ZN(new_n606));
  INV_X1    g181(.A(G79), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n527), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n605), .A2(KEYINPUT78), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT78), .B1(new_n605), .B2(new_n609), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(new_n602), .ZN(G284));
  XOR2_X1   g188(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n602), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(new_n602), .B2(G168), .ZN(G280));
  XOR2_X1   g192(.A(KEYINPUT80), .B(G559), .Z(new_n618));
  OAI21_X1  g193(.A(new_n612), .B1(G860), .B2(new_n618), .ZN(G148));
  NAND2_X1  g194(.A1(new_n612), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n497), .A2(new_n486), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2100), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n495), .A2(G123), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT81), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n470), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n467), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n627), .A2(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT17), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n654), .B2(new_n651), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n656), .B2(new_n658), .ZN(new_n660));
  INV_X1    g235(.A(new_n651), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n657), .A3(new_n653), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n652), .A2(new_n657), .A3(new_n654), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G1981), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT84), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT83), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G6), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n593), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT87), .Z(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(G23), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n575), .B1(new_n578), .B2(new_n580), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n688), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT85), .B(G16), .Z(new_n700));
  MUX2_X1   g275(.A(G303), .B(G22), .S(new_n700), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1971), .ZN(new_n702));
  NOR4_X1   g277(.A1(new_n693), .A2(new_n694), .A3(new_n699), .A4(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n706));
  MUX2_X1   g281(.A(G290), .B(G24), .S(new_n700), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT86), .B(G1986), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n470), .A2(G131), .ZN(new_n712));
  INV_X1    g287(.A(G119), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n467), .A2(G107), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  OAI22_X1  g290(.A1(new_n506), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n717), .B2(new_n710), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n718), .A2(new_n720), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n709), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n705), .A2(new_n706), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  OR3_X1    g300(.A1(new_n724), .A2(KEYINPUT88), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT26), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n731), .A2(new_n732), .B1(G105), .B2(new_n486), .ZN(new_n733));
  INV_X1    g308(.A(G129), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n506), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n470), .A2(G141), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n710), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n710), .B2(G32), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT91), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n688), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n688), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n743), .B1(G1961), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G21), .ZN(new_n747));
  AOI21_X1  g322(.A(KEYINPUT92), .B1(new_n688), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(G168), .A2(G16), .ZN(new_n749));
  MUX2_X1   g324(.A(KEYINPUT92), .B(new_n748), .S(new_n749), .Z(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G1966), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n746), .B(new_n751), .C1(G1961), .C2(new_n745), .ZN(new_n752));
  INV_X1    g327(.A(new_n558), .ZN(new_n753));
  MUX2_X1   g328(.A(new_n753), .B(G19), .S(new_n700), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT89), .B(G1341), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT90), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G28), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT30), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n758), .B2(KEYINPUT30), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n759), .A2(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n764), .B1(new_n710), .B2(new_n633), .C1(new_n754), .C2(new_n756), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n710), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  INV_X1    g342(.A(G128), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n467), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n506), .A2(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n470), .B2(G140), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(new_n710), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2067), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n710), .A2(G33), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT25), .Z(new_n777));
  INV_X1    g352(.A(G139), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n469), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n497), .A2(G127), .ZN(new_n780));
  INV_X1    g355(.A(G115), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n463), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n779), .B1(new_n782), .B2(G2105), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n775), .B1(new_n783), .B2(new_n710), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n739), .A2(new_n742), .B1(new_n784), .B2(G2072), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n765), .A2(new_n774), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(G2072), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n700), .A2(G20), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT23), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G299), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G1966), .B2(new_n750), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n752), .A2(new_n786), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G4), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n612), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1348), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n710), .A2(G35), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G162), .B2(new_n710), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT29), .B(G2090), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G164), .A2(G29), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G27), .B2(G29), .ZN(new_n804));
  INV_X1    g379(.A(G2078), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n798), .A2(new_n802), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(G160), .A2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G34), .ZN(new_n810));
  AOI21_X1  g385(.A(G29), .B1(new_n810), .B2(KEYINPUT24), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(KEYINPUT24), .B2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G2084), .Z(new_n814));
  NOR3_X1   g389(.A1(new_n794), .A2(new_n808), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n726), .A2(new_n728), .A3(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  AOI22_X1  g392(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n525), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n530), .A2(G55), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n533), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(G860), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n612), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n819), .A2(new_n822), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n558), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  AOI21_X1  g405(.A(G860), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(KEYINPUT93), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(KEYINPUT93), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(G145));
  AOI21_X1  g410(.A(new_n508), .B1(new_n514), .B2(new_n513), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n772), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n737), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n839), .B(new_n840), .C1(KEYINPUT94), .C2(new_n783), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n783), .A2(KEYINPUT94), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n841), .B(new_n842), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n495), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n467), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G142), .B2(new_n470), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n625), .B(new_n848), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n717), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n843), .A2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(G160), .B(new_n633), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G162), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n859));
  INV_X1    g434(.A(new_n853), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n851), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n859), .B1(new_n861), .B2(new_n856), .ZN(new_n862));
  NOR4_X1   g437(.A1(new_n860), .A2(new_n851), .A3(KEYINPUT95), .A4(new_n857), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g440(.A1(new_n605), .A2(new_n609), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(G299), .Z(new_n867));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n828), .B(KEYINPUT96), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n620), .B(new_n870), .ZN(new_n871));
  MUX2_X1   g446(.A(new_n869), .B(new_n867), .S(new_n871), .Z(new_n872));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  XOR2_X1   g450(.A(G166), .B(new_n600), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n696), .B(new_n593), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n880));
  OAI21_X1  g455(.A(G868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g457(.A(new_n881), .B1(G868), .B2(new_n827), .ZN(G331));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n884));
  AOI21_X1  g459(.A(G168), .B1(G301), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n828), .ZN(new_n887));
  NAND2_X1  g462(.A1(G171), .A2(KEYINPUT97), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n885), .A3(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n869), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n894), .A3(new_n867), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n878), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n878), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n901), .A3(new_n897), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT43), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n905), .B2(KEYINPUT101), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT98), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n901), .B1(new_n898), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n896), .A2(KEYINPUT98), .A3(new_n897), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n912), .A2(KEYINPUT100), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT100), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n906), .B(new_n908), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n904), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n913), .A4(new_n899), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n899), .A2(new_n913), .A3(new_n903), .A4(new_n902), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT99), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n919), .B(new_n921), .C1(new_n913), .C2(new_n912), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n907), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n916), .A2(new_n923), .ZN(G397));
  NAND2_X1  g499(.A1(new_n515), .A2(new_n518), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT45), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n928), .B2(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n475), .A2(new_n485), .A3(G40), .A4(new_n487), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n737), .B(G1996), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n772), .B(G2067), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n717), .A2(new_n719), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n720), .B1(new_n712), .B2(new_n716), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n600), .B(G1986), .Z(new_n942));
  OAI21_X1  g517(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(new_n926), .C1(new_n509), .C2(new_n519), .ZN(new_n945));
  INV_X1    g520(.A(new_n932), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT105), .B1(new_n836), .B2(G1384), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n925), .A2(new_n949), .A3(new_n926), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n944), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n791), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT116), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n925), .B2(new_n926), .ZN(new_n954));
  AOI211_X1 g529(.A(KEYINPUT105), .B(G1384), .C1(new_n515), .C2(new_n518), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT50), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n946), .A3(new_n945), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT116), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n791), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(G299), .B(KEYINPUT57), .Z(new_n961));
  OAI21_X1  g536(.A(new_n926), .B1(new_n509), .B2(new_n519), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n836), .A2(new_n963), .A3(G1384), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n932), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT56), .B(G2072), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n960), .A2(new_n961), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n961), .B1(new_n960), .B2(new_n968), .ZN(new_n970));
  INV_X1    g545(.A(new_n612), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT118), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n948), .A2(new_n950), .A3(new_n944), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n946), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT73), .B1(new_n502), .B2(new_n508), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n515), .A2(new_n510), .A3(new_n518), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(new_n944), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n972), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(KEYINPUT118), .A3(new_n973), .A4(new_n946), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n797), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n946), .A2(new_n983), .A3(new_n948), .A4(new_n950), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT117), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n971), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n969), .B1(new_n970), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n932), .B1(new_n977), .B2(new_n944), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT116), .B(G1956), .C1(new_n988), .C2(new_n956), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n958), .B1(new_n957), .B2(new_n791), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n968), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n961), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT61), .A3(new_n969), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT121), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n993), .A2(new_n969), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n982), .A2(new_n985), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT60), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n971), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n982), .A2(KEYINPUT60), .A3(new_n985), .A4(new_n612), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT61), .ZN(new_n1005));
  INV_X1    g580(.A(new_n968), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n1006), .B(new_n992), .C1(new_n953), .C2(new_n959), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n970), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n964), .A2(new_n966), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT119), .B(G1996), .Z(new_n1010));
  NAND3_X1  g585(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(G1341), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1009), .A2(new_n1010), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n558), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT59), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1004), .A2(new_n1008), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n987), .B1(new_n998), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT123), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n948), .A2(new_n950), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n963), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n946), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1966), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT115), .B(G2084), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n980), .A2(new_n973), .A3(new_n946), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1021), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G168), .A2(new_n1021), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1020), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1029), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n932), .B1(new_n1022), .B2(new_n963), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1966), .B1(new_n1037), .B2(new_n1024), .ZN(new_n1038));
  OAI21_X1  g613(.A(G8), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(KEYINPUT123), .A3(new_n1033), .A4(new_n1032), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1032), .B1(new_n1030), .B2(KEYINPUT122), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT51), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1041), .A2(new_n1045), .B1(new_n1031), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1961), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n979), .A2(new_n1048), .A3(new_n981), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n966), .B(new_n805), .C1(KEYINPUT45), .C2(new_n977), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT124), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1054), .A3(new_n1051), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n930), .A2(KEYINPUT53), .A3(new_n805), .A4(new_n966), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1049), .A2(new_n1053), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G171), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1050), .A2(new_n1054), .A3(new_n1051), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1054), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1037), .A2(KEYINPUT53), .A3(new_n805), .A4(new_n1024), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(G301), .A3(new_n1062), .A4(new_n1049), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1063), .A3(KEYINPUT54), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1971), .B1(new_n964), .B2(new_n966), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT104), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT104), .ZN(new_n1068));
  INV_X1    g643(.A(G1971), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n965), .A2(new_n932), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1068), .B(new_n1069), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G2090), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n980), .A2(new_n1073), .A3(new_n973), .A4(new_n946), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1067), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G166), .A2(new_n1021), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT106), .B(KEYINPUT55), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n1079));
  OAI22_X1  g654(.A1(G166), .A2(new_n1021), .B1(KEYINPUT106), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1075), .A2(KEYINPUT107), .A3(G8), .A4(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1074), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1072), .ZN(new_n1084));
  OAI211_X1 g659(.A(G8), .B(new_n1081), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT107), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1066), .B1(G2090), .B2(new_n957), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1081), .B1(new_n1089), .B2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT111), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n566), .A2(G86), .B1(new_n530), .B2(G48), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n679), .B1(new_n1092), .B2(new_n589), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n593), .B2(new_n679), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1094), .B2(KEYINPUT49), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n591), .A2(new_n592), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n679), .A3(new_n1092), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1093), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1091), .A2(new_n1097), .A3(KEYINPUT49), .A4(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(new_n1011), .C1(new_n1095), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT49), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1094), .A2(KEYINPUT109), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT110), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT110), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1100), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1976), .ZN(new_n1110));
  NOR3_X1   g685(.A1(G288), .A2(KEYINPUT108), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT108), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n696), .B2(G1976), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n1011), .A3(G8), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT52), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(G288), .B2(new_n1110), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1114), .A2(new_n1011), .A3(G8), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT114), .B1(new_n1109), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1103), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1107), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1121), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1118), .A4(new_n1116), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1090), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1064), .A2(new_n1088), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1047), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1049), .A2(new_n1053), .A3(new_n1062), .A4(new_n1055), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(G171), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1132), .B2(G171), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1057), .A2(G171), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1131), .B1(new_n1137), .B2(KEYINPUT54), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1132), .A2(G171), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1132), .A2(new_n1133), .A3(G171), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT126), .B(new_n1139), .C1(new_n1143), .C2(new_n1136), .ZN(new_n1144));
  AND4_X1   g719(.A1(new_n1019), .A2(new_n1130), .A3(new_n1138), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1030), .A2(G168), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT112), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1125), .A2(new_n1148), .A3(new_n1118), .A4(new_n1116), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT112), .B1(new_n1109), .B2(new_n1119), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1075), .A2(G8), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1146), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1155), .A2(new_n1087), .A3(new_n1082), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1125), .A2(new_n1110), .A3(new_n696), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1097), .B(KEYINPUT113), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1021), .B(new_n1012), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1154), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1088), .A2(new_n1128), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1161), .A2(new_n1146), .A3(G168), .A4(new_n1030), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1046), .A2(new_n1031), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1031), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1030), .A2(KEYINPUT122), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1033), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1163), .B(new_n1164), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1161), .A2(new_n1169), .A3(new_n1143), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1163), .B1(new_n1171), .B2(new_n1164), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1160), .B(new_n1162), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n943), .B1(new_n1145), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT47), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n935), .A2(G1996), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT46), .Z(new_n1177));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n737), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(KEYINPUT127), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT127), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1186), .A2(KEYINPUT47), .A3(new_n1180), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n935), .A2(G1986), .A3(G290), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1188), .A2(KEYINPUT48), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1188), .A2(KEYINPUT48), .B1(new_n936), .B2(new_n941), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n772), .A2(new_n983), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n937), .A2(new_n938), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1191), .B1(new_n1192), .B2(new_n939), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1189), .A2(new_n1190), .B1(new_n936), .B2(new_n1193), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1183), .A2(new_n1187), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1174), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g771(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n1198), .A2(new_n864), .A3(new_n922), .ZN(G225));
  INV_X1    g773(.A(G225), .ZN(G308));
endmodule


