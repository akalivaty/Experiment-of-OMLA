//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(new_n464), .A3(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT69), .B1(new_n472), .B2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NOR4_X1   g049(.A1(new_n470), .A2(new_n471), .A3(new_n474), .A4(new_n464), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n463), .B(new_n469), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT71), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G125), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G160));
  INV_X1    g067(.A(G136), .ZN(new_n493));
  NOR2_X1   g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n476), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n466), .A2(new_n468), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  INV_X1    g073(.A(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(KEYINPUT3), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(new_n474), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n500), .A2(KEYINPUT69), .A3(KEYINPUT3), .A4(new_n501), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n497), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  XOR2_X1   g081(.A(new_n506), .B(KEYINPUT72), .Z(new_n507));
  AOI21_X1  g082(.A(new_n496), .B1(new_n507), .B2(G124), .ZN(G162));
  INV_X1    g083(.A(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT4), .B1(new_n476), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n509), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n484), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(G126), .A2(G2105), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n469), .B(new_n517), .C1(new_n473), .C2(new_n475), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n505), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n463), .A2(G114), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n523), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT74), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  INV_X1    g101(.A(new_n524), .ZN(new_n527));
  AOI211_X1 g102(.A(new_n526), .B(new_n527), .C1(new_n519), .C2(new_n521), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n516), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G164));
  XNOR2_X1  g105(.A(KEYINPUT5), .B(G543), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n531), .A2(new_n532), .A3(G88), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n532), .A2(G543), .ZN(new_n537));
  AOI211_X1 g112(.A(new_n533), .B(new_n536), .C1(G50), .C2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n532), .A2(new_n531), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n532), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G51), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT5), .B(G543), .Z(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n535), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(new_n553), .B2(new_n552), .ZN(new_n555));
  INV_X1    g130(.A(G90), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n541), .A2(new_n556), .B1(new_n545), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n555), .A2(new_n559), .ZN(G171));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n541), .A2(new_n561), .B1(new_n545), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n531), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n535), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n537), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(new_n541), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G91), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n531), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n535), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(G299));
  NAND2_X1  g154(.A1(new_n555), .A2(new_n559), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  XNOR2_X1  g157(.A(G166), .B(new_n582), .ZN(G303));
  NAND2_X1  g158(.A1(new_n575), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n537), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n575), .A2(G86), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT79), .Z(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n550), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n537), .B2(G48), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n541), .A2(new_n595), .B1(new_n545), .B2(new_n596), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT80), .Z(new_n598));
  AOI22_X1  g173(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n535), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(G290));
  AND3_X1   g176(.A1(new_n531), .A2(new_n532), .A3(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT81), .B(G66), .Z(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n550), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(new_n537), .B2(G54), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G321));
  XOR2_X1   g186(.A(G321), .B(KEYINPUT82), .Z(G284));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(new_n608), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(new_n566), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n609), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n608), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g199(.A(new_n479), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n625), .A2(new_n485), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  NAND2_X1  g204(.A1(KEYINPUT84), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(KEYINPUT84), .A2(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n507), .A2(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n635));
  INV_X1    g210(.A(G99), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n463), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n477), .B2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n633), .A2(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n648), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(new_n657), .A3(G14), .ZN(G401));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n661), .A2(new_n659), .A3(new_n662), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n659), .A3(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n640), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(G227));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(new_n677), .A3(new_n675), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n682), .C1(new_n677), .C2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  INV_X1    g263(.A(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(G229));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT86), .B(G16), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(G22), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n694), .A2(new_n700), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT34), .Z(new_n708));
  NOR2_X1   g283(.A1(G25), .A2(G29), .ZN(new_n709));
  OR2_X1    g284(.A1(G95), .A2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n711));
  INV_X1    g286(.A(G131), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n476), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n507), .B2(G119), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n709), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n696), .A2(G24), .ZN(new_n718));
  INV_X1    g293(.A(G290), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n696), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(new_n684), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n708), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT36), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n507), .A2(G128), .ZN(new_n727));
  OR2_X1    g302(.A1(G104), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n477), .B2(G140), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n726), .B1(new_n733), .B2(new_n724), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT88), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2067), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G33), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT89), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT25), .Z(new_n740));
  INV_X1    g315(.A(G139), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n476), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(KEYINPUT90), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(KEYINPUT90), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n743), .A2(new_n744), .B1(new_n463), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT91), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n738), .B1(new_n747), .B2(new_n724), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2072), .Z(new_n749));
  NOR2_X1   g324(.A1(new_n736), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n724), .B1(KEYINPUT24), .B2(G34), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(KEYINPUT24), .B2(G34), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n491), .B2(G29), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT93), .Z(new_n756));
  NOR2_X1   g331(.A1(G171), .A2(new_n701), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G5), .B2(new_n701), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n507), .A2(G129), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  INV_X1    g338(.A(G105), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n625), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n477), .B2(G141), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(new_n724), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n724), .B2(G32), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n756), .B(new_n760), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT94), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n696), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n566), .B2(new_n696), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT87), .B(G1341), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n617), .A2(new_n701), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G4), .B2(new_n701), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n695), .A2(G20), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT23), .Z(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G299), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1956), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT31), .B(G11), .Z(new_n787));
  INV_X1    g362(.A(G28), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(KEYINPUT30), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT92), .Z(new_n790));
  AOI21_X1  g365(.A(G29), .B1(new_n788), .B2(KEYINPUT30), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G168), .A2(new_n701), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n701), .B2(G21), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n786), .B(new_n797), .C1(new_n759), .C2(new_n758), .ZN(new_n798));
  INV_X1    g373(.A(new_n639), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n782), .B(new_n798), .C1(G29), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n770), .A2(new_n771), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n800), .B(new_n801), .C1(new_n754), .C2(new_n753), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n724), .A2(G35), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n724), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT29), .B(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n724), .A2(G27), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G164), .B2(new_n724), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2078), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n802), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n723), .A2(new_n750), .A3(new_n773), .A4(new_n810), .ZN(G150));
  INV_X1    g386(.A(G150), .ZN(G311));
  NAND2_X1  g387(.A1(G80), .A2(G543), .ZN(new_n813));
  INV_X1    g388(.A(G67), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n550), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n535), .B1(new_n815), .B2(KEYINPUT95), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(KEYINPUT95), .B2(new_n815), .ZN(new_n817));
  INV_X1    g392(.A(G93), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n541), .A2(new_n818), .B1(new_n545), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n620), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n817), .A2(new_n566), .A3(new_n821), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n617), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT96), .Z(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n830), .B2(new_n831), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n824), .B1(new_n833), .B2(new_n835), .ZN(G145));
  INV_X1    g411(.A(new_n628), .ZN(new_n837));
  INV_X1    g412(.A(new_n714), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n477), .A2(G142), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT99), .Z(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n841));
  INV_X1    g416(.A(G106), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n463), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n507), .B2(G130), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n838), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n840), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n714), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n845), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n837), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n845), .A2(new_n847), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT100), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n628), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n747), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n768), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n747), .A2(new_n859), .A3(new_n767), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n520), .B1(new_n505), .B2(new_n517), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n524), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n505), .A2(G138), .A3(new_n463), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n514), .B1(new_n868), .B2(KEYINPUT4), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n864), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n527), .B1(new_n519), .B2(new_n521), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n516), .A2(new_n871), .A3(KEYINPUT97), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n732), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n862), .A3(new_n861), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n851), .A2(new_n855), .A3(KEYINPUT101), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n858), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n856), .A2(new_n857), .A3(new_n875), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G162), .B(new_n491), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n799), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n884), .A3(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g465(.A1(new_n822), .A2(new_n609), .ZN(new_n891));
  XNOR2_X1  g466(.A(G290), .B(G305), .ZN(new_n892));
  XNOR2_X1  g467(.A(G166), .B(new_n703), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT42), .Z(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(G299), .A2(KEYINPUT102), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n617), .B1(G299), .B2(KEYINPUT102), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n614), .A2(new_n617), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n897), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n614), .A2(new_n902), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n617), .A3(new_n898), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n900), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n827), .B(new_n622), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n901), .B2(new_n903), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n910), .B1(new_n914), .B2(new_n909), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n895), .B1(new_n896), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n896), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n895), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n891), .B1(new_n918), .B2(new_n609), .ZN(G295));
  XNOR2_X1  g494(.A(G295), .B(KEYINPUT105), .ZN(G331));
  NAND2_X1  g495(.A1(G171), .A2(G168), .ZN(new_n921));
  NAND2_X1  g496(.A1(G301), .A2(G286), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n827), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(new_n825), .A3(new_n826), .A4(new_n922), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(KEYINPUT108), .A3(new_n827), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n907), .A3(new_n906), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(KEYINPUT107), .A3(new_n926), .ZN(new_n931));
  OR3_X1    g506(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n827), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n904), .A2(new_n908), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n933), .A3(new_n894), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n934), .B2(KEYINPUT109), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n930), .A2(new_n933), .A3(new_n936), .A4(new_n894), .ZN(new_n937));
  INV_X1    g512(.A(new_n894), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n914), .B1(new_n932), .B2(new_n931), .ZN(new_n939));
  AND4_X1   g514(.A1(new_n908), .A2(new_n904), .A3(new_n927), .A4(new_n928), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n930), .A2(new_n933), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n938), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n935), .A2(new_n944), .A3(new_n937), .A4(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n944), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n937), .A4(new_n946), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(KEYINPUT119), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n490), .A2(G40), .A3(new_n478), .A4(new_n481), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n529), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n872), .A4(new_n958), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n957), .B(new_n961), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n699), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n529), .A2(new_n968), .A3(new_n958), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n958), .B1(new_n867), .B2(new_n869), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n956), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT118), .ZN(new_n973));
  AOI21_X1  g548(.A(G2090), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(KEYINPUT118), .A3(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n955), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(G303), .A2(G8), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT55), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n954), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n516), .B2(new_n871), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n955), .B1(new_n957), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n703), .A2(G1976), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT114), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n986), .B(new_n987), .C1(G1976), .C2(new_n703), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n589), .A2(new_n990), .A3(new_n689), .A4(new_n593), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n593), .A2(new_n588), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G1981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n992), .B(new_n994), .C1(KEYINPUT116), .C2(KEYINPUT49), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n983), .A3(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n988), .B(new_n999), .C1(new_n987), .C2(new_n986), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n970), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n867), .A2(new_n526), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n871), .A2(KEYINPUT74), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1005), .B2(new_n516), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n957), .B(new_n1002), .C1(new_n1006), .C2(new_n968), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(G2090), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n955), .B1(new_n967), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n979), .B(KEYINPUT113), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n699), .A2(new_n966), .B1(new_n974), .B2(new_n975), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT119), .B(new_n979), .C1(new_n1012), .C2(new_n955), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n968), .B1(new_n529), .B2(new_n958), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n956), .A2(G2084), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1014), .A2(new_n1001), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n960), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n529), .A2(new_n958), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n956), .B1(new_n970), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1966), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G286), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n981), .A2(new_n1011), .A3(new_n1013), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT63), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1007), .A2(G2090), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n699), .B2(new_n966), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n979), .B1(new_n1029), .B2(new_n955), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1023), .A2(new_n1026), .A3(G286), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1011), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1011), .A2(KEYINPUT120), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1027), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(G299), .B(KEYINPUT57), .Z(new_n1037));
  INV_X1    g612(.A(G1956), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n972), .A2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT56), .B(G2072), .Z(new_n1040));
  OAI211_X1 g615(.A(new_n1037), .B(new_n1039), .C1(new_n966), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n957), .A2(new_n982), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G2067), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n1007), .B2(new_n780), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(new_n608), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1039), .B1(new_n966), .B2(new_n1040), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1041), .ZN(new_n1051));
  NOR2_X1   g626(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1051), .A2(KEYINPUT61), .B1(new_n1041), .B2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n962), .A2(new_n963), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n962), .A2(new_n963), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1055), .A2(new_n1056), .B1(new_n960), .B2(new_n959), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n956), .A2(G1996), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT58), .B(G1341), .Z(new_n1060));
  AND2_X1   g635(.A1(new_n1042), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n566), .B(new_n1054), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1054), .A2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1057), .A2(new_n1058), .B1(new_n1042), .B2(new_n1060), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n620), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n617), .B(new_n1043), .C1(new_n1007), .C2(new_n780), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT60), .B1(new_n1045), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1044), .A2(new_n1069), .A3(new_n617), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1062), .A2(new_n1066), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1050), .B1(new_n1053), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n981), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n966), .B2(G2078), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(G2078), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1019), .A2(new_n1021), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1007), .A2(new_n759), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(G301), .B(KEYINPUT54), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n795), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1002), .B(new_n1015), .C1(new_n1006), .C2(new_n968), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1082), .B(G8), .C1(new_n1086), .C2(G286), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G168), .A2(new_n955), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1023), .A2(KEYINPUT51), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1092));
  AOI211_X1 g667(.A(KEYINPUT123), .B(new_n1089), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1087), .B(new_n1090), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n488), .A2(G40), .A3(new_n1076), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n482), .B(KEYINPUT124), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n873), .A2(new_n958), .ZN(new_n1097));
  AOI211_X1 g672(.A(new_n1095), .B(new_n1096), .C1(new_n1097), .C2(new_n960), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1080), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1081), .A2(new_n1094), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1073), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1072), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G288), .A2(G1976), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n999), .A2(new_n1105), .B1(new_n989), .B2(new_n991), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(KEYINPUT117), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n983), .B1(new_n1106), .B2(KEYINPUT117), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1107), .A2(new_n1108), .B1(new_n1109), .B2(new_n1000), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1079), .A2(G171), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1094), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1088), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT123), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1086), .A2(new_n1091), .A3(new_n1088), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1117), .A2(KEYINPUT62), .A3(new_n1090), .A4(new_n1087), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1111), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n981), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1110), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1036), .A2(new_n1104), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1097), .A2(new_n960), .A3(new_n957), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1123), .A2(G1986), .A3(G290), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1018), .B(new_n956), .C1(new_n873), .C2(new_n958), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n719), .A2(new_n684), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n1127), .B(KEYINPUT111), .Z(new_n1128));
  INV_X1    g703(.A(G2067), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n732), .B(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1996), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n767), .B(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n714), .B(new_n716), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n1123), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1128), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1122), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n714), .A2(new_n716), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1133), .A2(new_n1140), .B1(G2067), .B2(new_n732), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1125), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1123), .B1(new_n1130), .B2(new_n768), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT46), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1123), .A2(new_n1146), .A3(G1996), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT46), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT47), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1135), .A2(new_n1123), .B1(KEYINPUT48), .B2(new_n1124), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(KEYINPUT48), .B2(new_n1124), .ZN(new_n1152));
  OR4_X1    g727(.A1(new_n1139), .A2(new_n1144), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1144), .A2(new_n1152), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1139), .B1(new_n1154), .B2(new_n1150), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1138), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g732(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1159));
  NOR2_X1   g733(.A1(G229), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g734(.A1(new_n1160), .A2(new_n949), .A3(new_n950), .ZN(new_n1161));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n884), .B1(new_n880), .B2(new_n881), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n888), .A2(new_n887), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n1161), .B(new_n1162), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g739(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n889), .B2(new_n1161), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1167), .ZN(G308));
  NAND2_X1  g742(.A1(new_n889), .A2(new_n1161), .ZN(G225));
endmodule


