

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596;

  INV_X1 U328 ( .A(KEYINPUT55), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n408), .B(n318), .ZN(n540) );
  XOR2_X1 U330 ( .A(KEYINPUT37), .B(n498), .Z(n296) );
  XNOR2_X1 U331 ( .A(n320), .B(KEYINPUT31), .ZN(n321) );
  XNOR2_X1 U332 ( .A(n426), .B(n321), .ZN(n322) );
  XNOR2_X1 U333 ( .A(G99GAT), .B(G71GAT), .ZN(n303) );
  XNOR2_X1 U334 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U335 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n403) );
  XNOR2_X1 U336 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U337 ( .A(n404), .B(n403), .ZN(n557) );
  XNOR2_X1 U338 ( .A(n500), .B(KEYINPUT38), .ZN(n508) );
  XNOR2_X1 U339 ( .A(n461), .B(G190GAT), .ZN(n462) );
  XNOR2_X1 U340 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(G176GAT), .B(G183GAT), .Z(n298) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U344 ( .A(KEYINPUT86), .B(KEYINPUT18), .Z(n300) );
  XNOR2_X1 U345 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U347 ( .A(n302), .B(n301), .Z(n408) );
  XNOR2_X1 U348 ( .A(n303), .B(G120GAT), .ZN(n333) );
  XOR2_X1 U349 ( .A(G43GAT), .B(G134GAT), .Z(n367) );
  XNOR2_X1 U350 ( .A(n333), .B(n367), .ZN(n304) );
  AND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  NAND2_X1 U352 ( .A1(n304), .A2(n305), .ZN(n309) );
  INV_X1 U353 ( .A(n304), .ZN(n307) );
  INV_X1 U354 ( .A(n305), .ZN(n306) );
  NAND2_X1 U355 ( .A1(n307), .A2(n306), .ZN(n308) );
  NAND2_X1 U356 ( .A1(n309), .A2(n308), .ZN(n310) );
  XOR2_X1 U357 ( .A(n310), .B(KEYINPUT20), .Z(n313) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n311), .B(KEYINPUT83), .ZN(n446) );
  XNOR2_X1 U360 ( .A(n446), .B(KEYINPUT87), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n315) );
  INV_X1 U362 ( .A(KEYINPUT85), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n317) );
  XOR2_X1 U364 ( .A(G15GAT), .B(G127GAT), .Z(n342) );
  XNOR2_X1 U365 ( .A(n342), .B(KEYINPUT84), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  INV_X1 U367 ( .A(n540), .ZN(n530) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(G78GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n319), .B(G148GAT), .ZN(n426) );
  AND2_X1 U370 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n322), .B(G176GAT), .ZN(n327) );
  XOR2_X1 U372 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n324) );
  XOR2_X1 U373 ( .A(G85GAT), .B(G92GAT), .Z(n359) );
  XOR2_X1 U374 ( .A(G204GAT), .B(G64GAT), .Z(n412) );
  XNOR2_X1 U375 ( .A(n359), .B(n412), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U377 ( .A(n325), .B(KEYINPUT33), .Z(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n329) );
  XNOR2_X1 U380 ( .A(KEYINPUT71), .B(KEYINPUT32), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U383 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n332), .B(KEYINPUT13), .ZN(n338) );
  XNOR2_X1 U385 ( .A(n333), .B(n338), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n588) );
  XOR2_X1 U387 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n341) );
  XOR2_X1 U388 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n337) );
  XNOR2_X1 U389 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n346) );
  XOR2_X1 U393 ( .A(G22GAT), .B(G155GAT), .Z(n421) );
  XOR2_X1 U394 ( .A(n421), .B(n342), .Z(n344) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U397 ( .A(n346), .B(n345), .Z(n351) );
  XOR2_X1 U398 ( .A(G8GAT), .B(G1GAT), .Z(n387) );
  XOR2_X1 U399 ( .A(G78GAT), .B(G211GAT), .Z(n348) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G71GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n387), .B(n349), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n591) );
  XOR2_X1 U404 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n353) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n352) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n372) );
  XOR2_X1 U407 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n355) );
  XNOR2_X1 U408 ( .A(G99GAT), .B(KEYINPUT77), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U410 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XOR2_X1 U411 ( .A(n356), .B(n422), .Z(n358) );
  XNOR2_X1 U412 ( .A(G190GAT), .B(G218GAT), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U414 ( .A(n359), .B(KEYINPUT10), .Z(n361) );
  NAND2_X1 U415 ( .A1(G232GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n370) );
  XOR2_X1 U418 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n365) );
  XNOR2_X1 U419 ( .A(G36GAT), .B(G29GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U421 ( .A(KEYINPUT7), .B(n366), .ZN(n393) );
  INV_X1 U422 ( .A(n393), .ZN(n368) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n568) );
  XNOR2_X1 U426 ( .A(KEYINPUT36), .B(n568), .ZN(n593) );
  NAND2_X1 U427 ( .A1(n591), .A2(n593), .ZN(n375) );
  XOR2_X1 U428 ( .A(KEYINPUT114), .B(KEYINPUT45), .Z(n373) );
  XNOR2_X1 U429 ( .A(KEYINPUT64), .B(n373), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n394) );
  XOR2_X1 U431 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n377) );
  XNOR2_X1 U432 ( .A(KEYINPUT69), .B(KEYINPUT67), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n391) );
  XOR2_X1 U434 ( .A(G22GAT), .B(G141GAT), .Z(n379) );
  XNOR2_X1 U435 ( .A(G43GAT), .B(G50GAT), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U437 ( .A(G113GAT), .B(G15GAT), .Z(n381) );
  XNOR2_X1 U438 ( .A(G169GAT), .B(G197GAT), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U440 ( .A(n383), .B(n382), .Z(n389) );
  XOR2_X1 U441 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n385) );
  NAND2_X1 U442 ( .A1(G229GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U446 ( .A(n391), .B(n390), .Z(n392) );
  XOR2_X1 U447 ( .A(n393), .B(n392), .Z(n558) );
  NAND2_X1 U448 ( .A1(n394), .A2(n558), .ZN(n395) );
  NOR2_X1 U449 ( .A1(n588), .A2(n395), .ZN(n396) );
  XOR2_X1 U450 ( .A(KEYINPUT115), .B(n396), .Z(n402) );
  XNOR2_X1 U451 ( .A(KEYINPUT41), .B(n588), .ZN(n510) );
  OR2_X1 U452 ( .A1(n510), .A2(n558), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n397), .B(KEYINPUT46), .ZN(n399) );
  INV_X1 U454 ( .A(n568), .ZN(n550) );
  INV_X1 U455 ( .A(n591), .ZN(n546) );
  AND2_X1 U456 ( .A1(n550), .A2(n546), .ZN(n398) );
  AND2_X1 U457 ( .A1(n399), .A2(n398), .ZN(n400) );
  XOR2_X1 U458 ( .A(n400), .B(KEYINPUT47), .Z(n401) );
  NOR2_X1 U459 ( .A1(n402), .A2(n401), .ZN(n404) );
  XOR2_X1 U460 ( .A(KEYINPUT21), .B(G218GAT), .Z(n406) );
  XNOR2_X1 U461 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U463 ( .A(G197GAT), .B(n407), .Z(n433) );
  XNOR2_X1 U464 ( .A(n408), .B(n433), .ZN(n416) );
  XOR2_X1 U465 ( .A(KEYINPUT94), .B(G92GAT), .Z(n410) );
  XNOR2_X1 U466 ( .A(G36GAT), .B(G8GAT), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U468 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n527) );
  NOR2_X1 U472 ( .A1(n557), .A2(n527), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n417), .B(KEYINPUT54), .ZN(n581) );
  XOR2_X1 U474 ( .A(KEYINPUT91), .B(KEYINPUT2), .Z(n419) );
  XNOR2_X1 U475 ( .A(KEYINPUT3), .B(KEYINPUT90), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U477 ( .A(G141GAT), .B(n420), .Z(n445) );
  XOR2_X1 U478 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n424) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U481 ( .A(n425), .B(KEYINPUT92), .Z(n431) );
  XOR2_X1 U482 ( .A(n426), .B(KEYINPUT24), .Z(n428) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n429), .B(G204GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n445), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n473) );
  XOR2_X1 U489 ( .A(KEYINPUT79), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U490 ( .A(G29GAT), .B(G148GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U492 ( .A(G134GAT), .B(G85GAT), .Z(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n452) );
  XOR2_X1 U494 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n440) );
  XNOR2_X1 U495 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U497 ( .A(G57GAT), .B(G155GAT), .Z(n442) );
  XNOR2_X1 U498 ( .A(G127GAT), .B(G120GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n450) );
  XOR2_X1 U501 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n448) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n454) );
  NAND2_X1 U506 ( .A1(G225GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n580) );
  INV_X1 U508 ( .A(n580), .ZN(n554) );
  NOR2_X1 U509 ( .A1(n473), .A2(n554), .ZN(n455) );
  AND2_X1 U510 ( .A1(n581), .A2(n455), .ZN(n459) );
  XNOR2_X1 U511 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n457) );
  NOR2_X1 U512 ( .A1(n530), .A2(n460), .ZN(n577) );
  NAND2_X1 U513 ( .A1(n577), .A2(n568), .ZN(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT127), .B(KEYINPUT58), .Z(n461) );
  NAND2_X1 U515 ( .A1(n473), .A2(n530), .ZN(n464) );
  XNOR2_X1 U516 ( .A(n464), .B(KEYINPUT26), .ZN(n583) );
  XNOR2_X1 U517 ( .A(n527), .B(KEYINPUT95), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n465), .B(KEYINPUT27), .ZN(n475) );
  INV_X1 U519 ( .A(n475), .ZN(n466) );
  NOR2_X1 U520 ( .A1(n583), .A2(n466), .ZN(n555) );
  INV_X1 U521 ( .A(n527), .ZN(n486) );
  AND2_X1 U522 ( .A1(n540), .A2(n486), .ZN(n467) );
  NOR2_X1 U523 ( .A1(n473), .A2(n467), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT25), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT97), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n555), .A2(n470), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n471), .A2(n554), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT98), .ZN(n479) );
  XOR2_X1 U529 ( .A(n530), .B(KEYINPUT88), .Z(n477) );
  XNOR2_X1 U530 ( .A(KEYINPUT28), .B(n473), .ZN(n507) );
  NOR2_X1 U531 ( .A1(n580), .A2(n507), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n539) );
  XNOR2_X1 U533 ( .A(n539), .B(KEYINPUT96), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n495) );
  NAND2_X1 U536 ( .A1(n591), .A2(n550), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n480), .B(KEYINPUT82), .ZN(n481) );
  XNOR2_X1 U538 ( .A(n481), .B(KEYINPUT16), .ZN(n482) );
  NOR2_X1 U539 ( .A1(n495), .A2(n482), .ZN(n512) );
  NOR2_X1 U540 ( .A1(n588), .A2(n558), .ZN(n499) );
  NAND2_X1 U541 ( .A1(n512), .A2(n499), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(KEYINPUT99), .ZN(n491) );
  NAND2_X1 U543 ( .A1(n554), .A2(n491), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(KEYINPUT100), .ZN(n488) );
  NAND2_X1 U547 ( .A1(n491), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U550 ( .A1(n491), .A2(n540), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n493) );
  NAND2_X1 U553 ( .A1(n491), .A2(n507), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(n494), .ZN(G1327GAT) );
  NOR2_X1 U556 ( .A1(n591), .A2(n495), .ZN(n496) );
  NAND2_X1 U557 ( .A1(n593), .A2(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT103), .B(n497), .ZN(n498) );
  NAND2_X1 U559 ( .A1(n499), .A2(n296), .ZN(n500) );
  NOR2_X1 U560 ( .A1(n508), .A2(n580), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n527), .A2(n508), .ZN(n503) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  INV_X1 U565 ( .A(KEYINPUT40), .ZN(n505) );
  NOR2_X1 U566 ( .A1(n530), .A2(n508), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(G43GAT), .ZN(G1330GAT) );
  INV_X1 U569 ( .A(n507), .ZN(n535) );
  NOR2_X1 U570 ( .A1(n508), .A2(n535), .ZN(n509) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  INV_X1 U572 ( .A(n510), .ZN(n574) );
  NAND2_X1 U573 ( .A1(n558), .A2(n574), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT105), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n512), .A2(n525), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n520), .A2(n580), .ZN(n516) );
  XOR2_X1 U577 ( .A(KEYINPUT104), .B(KEYINPUT106), .Z(n514) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n527), .A2(n520), .ZN(n517) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n530), .A2(n520), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n535), .ZN(n524) );
  XOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n522) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT108), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NAND2_X1 U591 ( .A1(n296), .A2(n525), .ZN(n534) );
  NOR2_X1 U592 ( .A1(n580), .A2(n534), .ZN(n526) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n526), .Z(G1336GAT) );
  NOR2_X1 U594 ( .A1(n527), .A2(n534), .ZN(n528) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(n528), .Z(n529) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U597 ( .A1(n530), .A2(n534), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G99GAT), .B(n533), .ZN(G1338GAT) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NOR2_X1 U605 ( .A1(n557), .A2(n539), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n558), .A2(n549), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  NOR2_X1 U610 ( .A1(n510), .A2(n549), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n549), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(n547), .Z(n548) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n567) );
  INV_X1 U622 ( .A(n558), .ZN(n584) );
  NAND2_X1 U623 ( .A1(n567), .A2(n584), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n561) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT52), .B(n562), .Z(n564) );
  NAND2_X1 U629 ( .A1(n567), .A2(n574), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  XOR2_X1 U631 ( .A(G155GAT), .B(KEYINPUT121), .Z(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n591), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n577), .A2(n584), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT56), .B(n573), .Z(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U644 ( .A1(n577), .A2(n591), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n586) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n594) );
  NAND2_X1 U650 ( .A1(n594), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(n587), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .Z(n590) );
  NAND2_X1 U654 ( .A1(n594), .A2(n588), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  NAND2_X1 U656 ( .A1(n594), .A2(n591), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n595), .B(KEYINPUT62), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

