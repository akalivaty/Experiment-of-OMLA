//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OR3_X1    g0007(.A1(new_n207), .A2(KEYINPUT64), .A3(G13), .ZN(new_n208));
  OAI21_X1  g0008(.A(KEYINPUT64), .B1(new_n207), .B2(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n206), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n214), .A2(KEYINPUT0), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(KEYINPUT0), .B2(new_n214), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n201), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G97), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n227), .B1(new_n202), .B2(new_n228), .C1(new_n229), .C2(new_n212), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n207), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n221), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G222), .A2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G223), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n257), .B(new_n258), .C1(G77), .C2(new_n253), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n215), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(new_n251), .B2(new_n260), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT65), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n264), .A2(new_n266), .A3(new_n269), .A4(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n258), .A2(new_n262), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G226), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n259), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n273), .A2(G179), .ZN(new_n274));
  OAI21_X1  g0074(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n216), .A2(G33), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n275), .B1(new_n276), .B2(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n215), .B1(new_n207), .B2(new_n251), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n267), .A2(KEYINPUT66), .A3(G13), .A4(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n281), .A2(new_n282), .B1(new_n201), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n282), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n216), .A2(G1), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(G50), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n274), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n273), .A2(G200), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n301), .B1(new_n302), .B2(new_n273), .C1(new_n303), .C2(new_n296), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT9), .B1(new_n289), .B2(new_n295), .ZN(new_n305));
  OR3_X1    g0105(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT10), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n288), .A2(new_n224), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n278), .A2(new_n201), .B1(new_n216), .B2(G68), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n280), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n282), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT11), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT67), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n291), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n287), .A2(new_n290), .A3(KEYINPUT67), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n294), .A2(G68), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n311), .B(new_n316), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n228), .A2(G1698), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n253), .B(new_n323), .C1(G226), .C2(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n266), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n271), .A2(G238), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n270), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT13), .B1(new_n326), .B2(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(G169), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n333), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n333), .B2(G169), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n322), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n333), .A2(new_n302), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n331), .B2(new_n332), .ZN(new_n342));
  OR3_X1    g0142(.A1(new_n340), .A2(new_n322), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n250), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT68), .B(G33), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(KEYINPUT3), .ZN(new_n347));
  NOR2_X1   g0147(.A1(G223), .A2(G1698), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n223), .B2(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G87), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n266), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT69), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n347), .A2(new_n349), .B1(G33), .B2(G87), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT69), .B1(new_n355), .B2(new_n266), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n271), .A2(G232), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n270), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(G190), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n341), .B1(new_n352), .B2(new_n358), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n252), .B1(new_n346), .B2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(G20), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n250), .A2(new_n252), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n216), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n365), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n224), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(G58), .B(G68), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n363), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT68), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G33), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n250), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n380), .B2(new_n365), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n347), .A2(KEYINPUT7), .A3(G20), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT16), .B(new_n373), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n375), .A2(new_n282), .A3(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n291), .A2(new_n279), .A3(new_n293), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n288), .B2(new_n279), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n362), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n362), .A2(KEYINPUT17), .A3(new_n384), .A4(new_n386), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n384), .A2(new_n386), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n350), .A2(new_n351), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n258), .ZN(new_n394));
  INV_X1    g0194(.A(new_n358), .ZN(new_n395));
  AOI21_X1  g0195(.A(G169), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n353), .B1(new_n393), .B2(new_n258), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n355), .A2(KEYINPUT69), .A3(new_n266), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n358), .A2(G179), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n392), .A2(new_n401), .A3(KEYINPUT18), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n391), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(G232), .A2(G1698), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n255), .A2(G238), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n253), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n258), .C1(G107), .C2(new_n253), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n271), .A2(G244), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n270), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n297), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G179), .B2(new_n413), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n320), .A2(new_n313), .A3(new_n293), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n417), .A2(new_n280), .B1(new_n216), .B2(new_n313), .ZN(new_n418));
  INV_X1    g0218(.A(new_n279), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n277), .B2(new_n419), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n290), .B1(G77), .B2(new_n287), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n415), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n413), .A2(G200), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n422), .B(new_n425), .C1(new_n302), .C2(new_n413), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n309), .A2(new_n344), .A3(new_n407), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT19), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n216), .B1(new_n325), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G87), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n229), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n216), .A2(G33), .A3(G97), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n430), .A2(new_n433), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n379), .A2(new_n250), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n216), .A2(G68), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n282), .B1(new_n288), .B2(new_n417), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n267), .A2(G33), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n292), .A2(G87), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n225), .A2(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n376), .A2(new_n378), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n347), .A2(new_n443), .B1(G116), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n347), .A2(KEYINPUT73), .A3(G244), .A4(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n379), .A2(G244), .A3(G1698), .A4(new_n250), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT73), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n258), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n261), .A2(G1), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n453), .A2(G274), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n206), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n266), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n442), .B1(new_n457), .B2(G200), .ZN(new_n458));
  INV_X1    g0258(.A(new_n456), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n450), .B2(new_n258), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(G190), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n451), .A2(G190), .A3(new_n456), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT75), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT76), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n457), .A2(new_n297), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n460), .A2(new_n336), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n438), .A2(new_n282), .ZN(new_n469));
  INV_X1    g0269(.A(new_n417), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n287), .A2(new_n290), .A3(new_n470), .A4(new_n440), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n288), .A2(new_n417), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT74), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n439), .A2(KEYINPUT74), .A3(new_n471), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n467), .A2(new_n468), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n465), .A2(new_n466), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n466), .B1(new_n465), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n212), .A2(G1698), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G303), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n436), .A2(new_n483), .B1(new_n484), .B2(new_n253), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT78), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n213), .A2(new_n255), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n347), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n379), .A2(new_n250), .A3(new_n487), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT78), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n485), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT5), .B(G41), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n452), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G270), .A3(new_n266), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n266), .A2(G274), .A3(new_n492), .A4(new_n452), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT77), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n494), .A2(KEYINPUT77), .A3(new_n495), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n491), .A2(new_n266), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n267), .B2(G33), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n318), .A2(new_n319), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT79), .B1(new_n287), .B2(G116), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT79), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n285), .A2(new_n503), .A3(new_n499), .A4(new_n286), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n505), .B(new_n216), .C1(G33), .C2(new_n229), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n499), .A2(G20), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n282), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n506), .A2(new_n282), .A3(KEYINPUT20), .A4(new_n507), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n502), .A2(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n297), .B1(new_n501), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n498), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT21), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  AOI211_X1 g0317(.A(KEYINPUT80), .B(new_n517), .C1(new_n498), .C2(new_n513), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n488), .A2(new_n490), .ZN(new_n520));
  INV_X1    g0320(.A(new_n485), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n496), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n494), .A2(KEYINPUT77), .A3(new_n495), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n522), .A2(new_n258), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n501), .A2(new_n512), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(G179), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n498), .B2(G200), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n302), .B2(new_n498), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n519), .A2(KEYINPUT81), .A3(new_n527), .A4(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n529), .B(new_n527), .C1(new_n516), .C2(new_n518), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n379), .A2(G244), .A3(new_n255), .A4(new_n250), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n255), .A2(KEYINPUT4), .A3(G244), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n206), .B2(new_n255), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n253), .A2(new_n539), .B1(G33), .B2(G283), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n266), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n493), .A2(G257), .A3(new_n266), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n495), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT71), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT71), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n546), .A3(new_n495), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n542), .A2(new_n302), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n547), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n541), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n550), .B2(G200), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n287), .A2(G97), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n291), .B1(new_n267), .B2(G33), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G97), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n432), .B1(new_n367), .B2(new_n370), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n557), .A2(new_n229), .A3(G107), .ZN(new_n558));
  XNOR2_X1  g0358(.A(G97), .B(G107), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n560), .A2(new_n216), .B1(new_n313), .B2(new_n278), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n282), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT70), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n559), .A2(new_n557), .ZN(new_n564));
  INV_X1    g0364(.A(new_n558), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n364), .A2(new_n366), .B1(new_n369), .B2(new_n365), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(new_n432), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT70), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n282), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n555), .B1(new_n563), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n551), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n297), .B1(new_n549), .B2(new_n541), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n542), .A2(new_n336), .A3(new_n545), .A4(new_n547), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT72), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n572), .A2(new_n576), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT72), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n551), .A2(new_n572), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(G250), .A2(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n212), .B2(G1698), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(new_n379), .A3(new_n250), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n444), .A2(G294), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n258), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n493), .A2(G264), .A3(new_n266), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n495), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G169), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n588), .A2(G179), .A3(new_n495), .A4(new_n589), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n595), .A2(new_n431), .A3(G20), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n379), .A2(new_n596), .A3(new_n250), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n250), .A2(new_n252), .A3(new_n216), .A4(G87), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n595), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT23), .B1(new_n216), .B2(G107), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT23), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n432), .A3(G20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n444), .A2(new_n216), .A3(G116), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n597), .A2(new_n599), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT24), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n598), .B2(new_n595), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT24), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n597), .A4(new_n605), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n290), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n285), .A2(new_n432), .A3(new_n286), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT25), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n287), .A2(new_n290), .A3(G107), .A4(new_n440), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n593), .B(new_n594), .C1(new_n611), .C2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n266), .B1(new_n585), .B2(new_n586), .ZN(new_n618));
  INV_X1    g0418(.A(new_n589), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n619), .A3(new_n336), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n495), .A2(new_n620), .B1(new_n590), .B2(G169), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n607), .A2(new_n610), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n616), .B1(new_n622), .B2(new_n282), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT82), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n590), .A2(G200), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n623), .B(new_n625), .C1(new_n302), .C2(new_n590), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n617), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n578), .A2(new_n582), .A3(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n428), .A2(new_n481), .A3(new_n534), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n481), .B2(new_n577), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n457), .A2(new_n297), .B1(new_n475), .B2(new_n476), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(new_n468), .B1(new_n458), .B2(new_n463), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n631), .A3(new_n577), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n527), .B1(new_n516), .B2(new_n518), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT83), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n593), .B(new_n637), .C1(new_n611), .C2(new_n616), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT83), .B1(new_n621), .B2(new_n623), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(new_n579), .A3(new_n581), .A4(new_n626), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n478), .B(new_n635), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n428), .B1(new_n632), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g0445(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n392), .A2(new_n401), .A3(KEYINPUT18), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT18), .B1(new_n392), .B2(new_n401), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n404), .A2(new_n405), .A3(new_n646), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n343), .A2(new_n423), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(new_n339), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n389), .A2(new_n390), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n306), .A2(new_n307), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n300), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n645), .A2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n267), .A2(new_n216), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n526), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n534), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n636), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n593), .B(new_n665), .C1(new_n611), .C2(new_n616), .ZN(new_n674));
  INV_X1    g0474(.A(new_n665), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n623), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n627), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n636), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n628), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n665), .B(KEYINPUT87), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n640), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(G399));
  NOR2_X1   g0485(.A1(new_n211), .A2(G41), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n433), .A2(G116), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n267), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n219), .B2(new_n686), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  NAND4_X1  g0491(.A1(new_n534), .A2(new_n629), .A3(new_n481), .A4(new_n681), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n590), .A2(new_n336), .ZN(new_n693));
  OR4_X1    g0493(.A1(new_n460), .A2(new_n525), .A3(new_n550), .A4(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n525), .A2(new_n550), .A3(new_n460), .A4(new_n620), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(KEYINPUT30), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(KEYINPUT30), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT31), .B1(new_n698), .B2(new_n665), .ZN(new_n699));
  INV_X1    g0499(.A(new_n681), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(KEYINPUT31), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n672), .B1(new_n692), .B2(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n460), .A2(new_n461), .A3(G190), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n439), .A2(new_n441), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n460), .B2(new_n341), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n461), .B1(new_n460), .B2(G190), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n467), .A2(new_n468), .A3(new_n477), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT76), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n465), .A2(new_n466), .A3(new_n478), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n631), .A3(new_n711), .A4(new_n577), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n634), .A2(new_n577), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n709), .B1(new_n713), .B2(KEYINPUT26), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT88), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n714), .A3(KEYINPUT88), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n617), .A2(new_n624), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n636), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n642), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n718), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n632), .A2(new_n643), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n700), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n703), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n691), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(new_n673), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n671), .A2(new_n672), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n216), .A2(G13), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n267), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n686), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT89), .Z(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(new_n731), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n210), .A2(new_n253), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT90), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(G355), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n211), .A2(new_n347), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G45), .B2(new_n218), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n247), .A2(new_n261), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(G116), .B2(new_n210), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n265), .B1(new_n216), .B2(G169), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT91), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT92), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n746), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n737), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n341), .A2(G190), .ZN(new_n757));
  OAI21_X1  g0557(.A(G20), .B1(new_n757), .B2(G179), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT93), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n229), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n216), .A2(new_n336), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n302), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n216), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n767), .A2(G50), .B1(new_n770), .B2(G87), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n302), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G107), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n766), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n771), .B(new_n774), .C1(new_n224), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G190), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G159), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n765), .A2(new_n778), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n757), .A2(new_n216), .A3(new_n336), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n253), .B1(new_n313), .B2(new_n783), .C1(new_n785), .C2(new_n202), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n777), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n759), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G294), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n780), .A2(G329), .B1(new_n784), .B2(G322), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n368), .C1(new_n791), .C2(new_n783), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT33), .B(G317), .Z(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n776), .A2(new_n793), .B1(new_n772), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n767), .A2(G326), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n484), .B2(new_n769), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n792), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n764), .A2(new_n787), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n756), .B1(new_n748), .B2(new_n799), .C1(new_n670), .C2(new_n752), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n738), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n424), .A2(KEYINPUT97), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n665), .B1(new_n416), .B2(new_n421), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT97), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n423), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n803), .A2(new_n426), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n423), .A2(new_n665), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n726), .B2(new_n700), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n681), .B(new_n809), .C1(new_n632), .C2(new_n643), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n703), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n736), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n811), .A2(new_n703), .A3(new_n812), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n748), .A2(new_n750), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT95), .Z(new_n818));
  OAI21_X1  g0618(.A(new_n736), .B1(new_n818), .B2(G77), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n785), .A2(new_n820), .B1(new_n779), .B2(new_n791), .ZN(new_n821));
  INV_X1    g0621(.A(new_n783), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n253), .B(new_n821), .C1(G116), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n772), .A2(new_n431), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G303), .B2(new_n767), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n775), .A2(G283), .B1(new_n770), .B2(G107), .ZN(new_n826));
  AND4_X1   g0626(.A1(new_n764), .A2(new_n823), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(KEYINPUT96), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n822), .A2(G159), .B1(new_n784), .B2(G143), .ZN(new_n830));
  INV_X1    g0630(.A(new_n767), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n276), .C2(new_n776), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n788), .A2(G58), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n201), .A2(new_n769), .B1(new_n772), .B2(new_n224), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n436), .B(new_n838), .C1(G132), .C2(new_n780), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n828), .A2(new_n829), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n748), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n819), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n809), .B2(new_n750), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n816), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  OAI211_X1 g0646(.A(G116), .B(new_n217), .C1(new_n566), .C2(KEYINPUT35), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(KEYINPUT98), .B1(KEYINPUT35), .B2(new_n566), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(KEYINPUT98), .B2(new_n847), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT36), .Z(new_n850));
  OAI211_X1 g0650(.A(new_n219), .B(G77), .C1(new_n202), .C2(new_n224), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n201), .A2(G68), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n267), .B(G13), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n663), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n652), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n322), .A2(new_n665), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n344), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n857), .B1(new_n339), .B2(new_n343), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n803), .A2(new_n806), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n675), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT99), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n812), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n373), .B1(new_n381), .B2(new_n382), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n363), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n383), .A2(new_n282), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n386), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n855), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n391), .B2(new_n406), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n392), .A2(new_n855), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n402), .A2(new_n873), .A3(new_n387), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n387), .A2(KEYINPUT37), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n870), .B1(new_n401), .B2(new_n855), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n866), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n648), .A2(new_n649), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n855), .B(new_n870), .C1(new_n882), .C2(new_n655), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n875), .A2(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n856), .B1(new_n865), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT39), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n872), .A2(new_n880), .A3(new_n866), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n873), .A2(new_n387), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n890), .B2(KEYINPUT85), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n874), .ZN(new_n892));
  INV_X1    g0692(.A(new_n890), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(KEYINPUT85), .A3(KEYINPUT37), .A4(new_n402), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n655), .B1(new_n650), .B2(new_n651), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n892), .B(new_n894), .C1(new_n895), .C2(new_n873), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n889), .B1(new_n896), .B2(new_n866), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n888), .B1(new_n897), .B2(KEYINPUT39), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n339), .A2(new_n665), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(KEYINPUT100), .A2(new_n887), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n887), .A2(KEYINPUT100), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n724), .A2(new_n428), .A3(new_n727), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n658), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT101), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(new_n699), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n692), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n809), .B1(new_n859), .B2(new_n860), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT40), .B1(new_n914), .B2(new_n897), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n881), .A2(new_n885), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(KEYINPUT101), .A2(KEYINPUT40), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n912), .B1(new_n692), .B2(new_n910), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n911), .A2(new_n428), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(G330), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n907), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n267), .B2(new_n732), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n907), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n854), .B1(new_n928), .B2(new_n929), .ZN(G367));
  NOR2_X1   g0730(.A1(new_n705), .A2(new_n675), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n634), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n709), .A2(KEYINPUT102), .A3(new_n931), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT102), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n478), .B2(new_n932), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n579), .B(new_n581), .C1(new_n572), .C2(new_n681), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n577), .A2(new_n700), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n939), .A2(KEYINPUT103), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT103), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n719), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n700), .B1(new_n945), .B2(new_n579), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n943), .A2(KEYINPUT42), .A3(new_n680), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT42), .B1(new_n943), .B2(new_n680), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n938), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n678), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n944), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT104), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n952), .A2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(KEYINPUT104), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n680), .B1(new_n679), .B2(new_n677), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n728), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n943), .A2(new_n683), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT45), .ZN(new_n966));
  NOR2_X1   g0766(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n944), .B2(new_n684), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n943), .B(new_n683), .C1(KEYINPUT105), .C2(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g0769(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n953), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n953), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n728), .B1(new_n964), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n686), .B(KEYINPUT41), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(KEYINPUT107), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT107), .ZN(new_n981));
  INV_X1    g0781(.A(new_n728), .ZN(new_n982));
  INV_X1    g0782(.A(new_n975), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n973), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n982), .B1(new_n984), .B2(new_n963), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n981), .B1(new_n985), .B2(new_n978), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n986), .A3(new_n733), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n960), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n937), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n751), .ZN(new_n990));
  INV_X1    g0790(.A(new_n742), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n991), .A2(new_n240), .B1(new_n210), .B2(new_n417), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n736), .B1(new_n754), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n762), .A2(new_n224), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n772), .A2(new_n313), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G159), .B2(new_n775), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n767), .A2(G143), .B1(new_n770), .B2(G58), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n368), .B1(new_n784), .B2(G150), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G50), .A2(new_n822), .B1(new_n780), .B2(G137), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n772), .A2(new_n229), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G311), .B2(new_n767), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n347), .B1(new_n775), .B2(G294), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n432), .C2(new_n759), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n780), .A2(G317), .B1(new_n784), .B2(G303), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT46), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n769), .B2(new_n499), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n822), .A2(G283), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n994), .A2(new_n1000), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT47), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n748), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n993), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n990), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n988), .A2(new_n1016), .ZN(G387));
  OR2_X1    g0817(.A1(new_n677), .A2(new_n752), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n822), .A2(G303), .B1(new_n784), .B2(G317), .ZN(new_n1019));
  INV_X1    g0819(.A(G322), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(new_n831), .B2(new_n1020), .C1(new_n791), .C2(new_n776), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n788), .A2(G283), .B1(G294), .B2(new_n770), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n772), .A2(new_n499), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n347), .B(new_n1030), .C1(G326), .C2(new_n780), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n775), .A2(new_n419), .B1(new_n770), .B2(G77), .ZN(new_n1033));
  INV_X1    g0833(.A(G159), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n831), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G68), .A2(new_n822), .B1(new_n780), .B2(G150), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n201), .B2(new_n785), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1035), .A2(new_n1037), .A3(new_n436), .A4(new_n1001), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n417), .B2(new_n762), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n748), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n754), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n740), .A2(new_n688), .B1(new_n432), .B2(new_n211), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n688), .C1(G68), .C2(G77), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1043), .A2(KEYINPUT108), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(KEYINPUT108), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT50), .B1(new_n279), .B2(G50), .ZN(new_n1046));
  OR3_X1    g0846(.A1(new_n279), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(KEYINPUT109), .A3(new_n742), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n261), .B2(new_n237), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT109), .B1(new_n1048), .B2(new_n742), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1042), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n737), .B(new_n1040), .C1(new_n1041), .C2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n963), .A2(new_n734), .B1(new_n1018), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n964), .A2(new_n686), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n963), .A2(new_n728), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(G393));
  NAND2_X1  g0857(.A1(new_n984), .A2(new_n734), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n742), .A2(new_n244), .B1(G97), .B2(new_n211), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1041), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n737), .B1(new_n1060), .B2(KEYINPUT110), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT110), .B2(new_n1060), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n368), .B1(new_n779), .B2(new_n1020), .C1(new_n820), .C2(new_n783), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n774), .B1(new_n794), .B2(new_n769), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(G303), .C2(new_n775), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n767), .A2(G317), .B1(G311), .B2(new_n784), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT52), .Z(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(new_n499), .C2(new_n759), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n767), .A2(G150), .B1(G159), .B2(new_n784), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT51), .Z(new_n1070));
  AOI21_X1  g0870(.A(new_n824), .B1(G68), .B2(new_n770), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n419), .A2(new_n822), .B1(new_n780), .B2(G143), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n775), .A2(G50), .ZN(new_n1073));
  AND4_X1   g0873(.A1(new_n347), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1070), .B(new_n1074), .C1(new_n762), .C2(new_n313), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n748), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1062), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n944), .B2(new_n752), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n984), .B1(new_n728), .B2(new_n963), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n686), .B1(new_n964), .B2(new_n976), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1058), .B(new_n1078), .C1(new_n1079), .C2(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(new_n861), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n862), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n426), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n721), .B1(new_n715), .B2(new_n716), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n665), .B(new_n1084), .C1(new_n1085), .C2(new_n718), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n863), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n896), .A2(new_n866), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n885), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n900), .B(KEYINPUT111), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n812), .A2(new_n864), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n1082), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n900), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1088), .A2(new_n1092), .B1(new_n1095), .B2(new_n898), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n809), .A2(G330), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n692), .B2(new_n910), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT112), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n1082), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1098), .B2(new_n1082), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT113), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n898), .B1(new_n865), .B2(new_n901), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1084), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n723), .A2(new_n675), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n861), .B1(new_n1106), .B2(new_n863), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT113), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1102), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n665), .B1(new_n1085), .B2(new_n718), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1087), .B1(new_n1113), .B2(new_n1105), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1092), .B1(new_n1114), .B2(new_n861), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n692), .A2(new_n702), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1097), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1082), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n1104), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1103), .A2(new_n734), .A3(new_n1112), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT115), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1122), .A2(KEYINPUT113), .B1(new_n1096), .B2(new_n1118), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT115), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n734), .A4(new_n1112), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n818), .A2(new_n419), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n737), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n776), .A2(new_n832), .B1(new_n783), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n762), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(G159), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT116), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n770), .A2(G150), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n368), .B1(new_n780), .B2(G125), .ZN(new_n1136));
  INV_X1    g0936(.A(G132), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n785), .ZN(new_n1138));
  INV_X1    g0938(.A(G128), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n831), .A2(new_n1139), .B1(new_n772), .B2(new_n201), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n253), .B1(G116), .B2(new_n784), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n229), .B2(new_n783), .C1(new_n820), .C2(new_n779), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n770), .A2(G87), .B1(new_n773), .B2(G68), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n432), .B2(new_n776), .C1(new_n794), .C2(new_n831), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(new_n1131), .C2(G77), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1128), .B1(new_n748), .B2(new_n1147), .C1(new_n899), .C2(new_n750), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT117), .Z(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n911), .A2(G330), .A3(new_n428), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT114), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n911), .A2(KEYINPUT114), .A3(G330), .A4(new_n428), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n658), .A3(new_n905), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1098), .A2(new_n1082), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT112), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n861), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1098), .A2(new_n1099), .A3(new_n1082), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1093), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1114), .B(new_n1118), .C1(new_n1082), .C2(new_n1098), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1156), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1102), .B1(new_n1115), .B2(new_n1104), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1119), .B1(new_n1167), .B2(new_n1110), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1112), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1166), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1103), .A2(new_n1165), .A3(new_n1112), .A4(new_n1119), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n686), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1126), .A2(new_n1150), .A3(new_n1172), .ZN(G378));
  INV_X1    g0973(.A(new_n1156), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n296), .A2(new_n855), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n308), .B(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n922), .B2(G330), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n672), .B(new_n1185), .C1(new_n915), .C2(new_n921), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n904), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1090), .B1(new_n920), .B2(new_n908), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1188), .A2(KEYINPUT40), .B1(new_n920), .B2(new_n919), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1185), .B1(new_n1189), .B2(new_n672), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n922), .A2(G330), .A3(new_n1183), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(new_n903), .A4(new_n902), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1176), .B1(new_n1187), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1175), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n686), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1175), .B2(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1185), .A2(new_n749), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n736), .B1(G50), .B2(new_n817), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n436), .A2(new_n260), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n994), .B1(G116), .B2(new_n767), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT119), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n769), .A2(new_n313), .B1(new_n779), .B2(new_n794), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1205), .B(new_n1201), .C1(G58), .C2(new_n773), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT118), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n822), .A2(new_n470), .B1(new_n784), .B2(G107), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n229), .B2(new_n776), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1204), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1202), .B1(new_n1210), .B2(KEYINPUT58), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT120), .Z(new_n1212));
  OAI22_X1  g1012(.A1(new_n785), .A2(new_n1139), .B1(new_n783), .B2(new_n832), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1129), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n770), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G125), .A2(new_n767), .B1(new_n775), .B2(G132), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n762), .C2(new_n276), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1034), .B2(new_n772), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1217), .B2(KEYINPUT59), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1210), .A2(KEYINPUT58), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1212), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1200), .B1(new_n1223), .B2(new_n842), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1196), .A2(new_n734), .B1(new_n1199), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1198), .A2(new_n1225), .ZN(G375));
  AND2_X1   g1026(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT121), .B1(new_n1227), .B2(new_n733), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT121), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n734), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n736), .B1(new_n818), .B2(G68), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n762), .A2(new_n417), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n995), .B1(G294), .B2(new_n767), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n775), .A2(G116), .B1(new_n770), .B2(G97), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n253), .B1(new_n822), .B2(G107), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n780), .A2(G303), .B1(new_n784), .B2(G283), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n762), .A2(new_n201), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n767), .A2(G132), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT122), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n785), .A2(new_n832), .B1(new_n783), .B2(new_n276), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G128), .B2(new_n780), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n436), .B1(G58), .B2(new_n773), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n775), .A2(new_n1214), .B1(new_n770), .B2(G159), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1241), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1233), .A2(new_n1238), .B1(new_n1239), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1232), .B1(new_n1247), .B2(new_n842), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1082), .B2(new_n750), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1228), .A2(new_n1231), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1227), .A2(new_n1156), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n979), .A3(new_n1166), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(G381));
  INV_X1    g1053(.A(G390), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n988), .A2(new_n1016), .A3(new_n1254), .ZN(new_n1255));
  OR3_X1    g1055(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1255), .A2(new_n1256), .A3(G381), .ZN(new_n1257));
  INV_X1    g1057(.A(G378), .ZN(new_n1258));
  INV_X1    g1058(.A(G375), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(G407));
  INV_X1    g1060(.A(KEYINPUT123), .ZN(new_n1261));
  INV_X1    g1061(.A(G213), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(G343), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n664), .A2(KEYINPUT123), .A3(G213), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT124), .Z(new_n1266));
  NAND3_X1  g1066(.A1(new_n1259), .A2(new_n1258), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(new_n1267), .A3(G213), .ZN(G409));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G378), .B(new_n1225), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n686), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1103), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(new_n1166), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1149), .B1(new_n1273), .B2(new_n1171), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1175), .A2(new_n979), .A3(new_n1196), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1225), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1126), .B(new_n1274), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1227), .B2(new_n1156), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1165), .A2(new_n1271), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1250), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n845), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1250), .B(G384), .C1(new_n1282), .C2(new_n1284), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AND4_X1   g1088(.A1(KEYINPUT126), .A2(new_n1278), .A3(new_n1265), .A4(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1265), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT126), .B1(new_n1291), .B2(new_n1288), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1269), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1266), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1288), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1286), .A2(new_n1287), .B1(G2897), .B2(new_n1266), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1290), .A2(G2897), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1288), .B2(new_n1297), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1298), .A2(new_n1291), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(new_n801), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1254), .B1(new_n988), .B2(new_n1016), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1016), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n1302), .B(G390), .C1(new_n960), .C2(new_n987), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n977), .A2(new_n979), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n734), .B1(new_n1306), .B2(new_n981), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n959), .B1(new_n1307), .B2(new_n980), .ZN(new_n1308));
  OAI21_X1  g1108(.A(G390), .B1(new_n1308), .B2(new_n1302), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1300), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1255), .A3(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1304), .A2(new_n1305), .A3(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1293), .A2(new_n1295), .A3(new_n1299), .A4(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1298), .B2(new_n1294), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1294), .A2(KEYINPUT62), .A3(new_n1288), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1315), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1304), .A2(new_n1311), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1313), .B1(new_n1319), .B2(new_n1321), .ZN(G405));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1258), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1270), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1288), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1288), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1323), .A2(new_n1326), .A3(new_n1270), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1320), .ZN(G402));
endmodule


