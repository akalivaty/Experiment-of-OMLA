//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n203), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G107), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n207), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(new_n203), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n207), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n229), .B(new_n232), .C1(new_n220), .C2(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n222), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n203), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(new_n214), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n226), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(KEYINPUT11), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n252), .A2(new_n262), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n227), .A2(G1), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G68), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n254), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT11), .B1(new_n260), .B2(new_n262), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n257), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G232), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G1698), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n274), .B(new_n276), .C1(G226), .C2(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G97), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  AND2_X1   g0083(.A1(G1), .A2(G13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n284), .A2(new_n285), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n287), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n291), .B2(new_n209), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n281), .A2(new_n282), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n282), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n290), .B1(new_n277), .B2(new_n278), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n292), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT69), .B1(new_n298), .B2(G200), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT69), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  AOI211_X1 g0101(.A(new_n300), .B(new_n301), .C1(new_n294), .C2(new_n297), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n270), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n296), .A2(new_n295), .A3(new_n292), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT13), .B1(new_n296), .B2(new_n292), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT70), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(KEYINPUT13), .C1(new_n296), .C2(new_n292), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT71), .B1(new_n309), .B2(G190), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(KEYINPUT71), .A3(G190), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n303), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n294), .B2(new_n297), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT14), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT72), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n315), .ZN(new_n322));
  AOI22_X1  g0122(.A1(KEYINPUT14), .A2(new_n322), .B1(new_n309), .B2(G179), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n270), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT73), .B1(new_n313), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n274), .A2(G222), .A3(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G77), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n274), .A2(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G223), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n327), .B(new_n331), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n280), .ZN(new_n335));
  INV_X1    g0135(.A(G226), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n289), .B1(new_n291), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n301), .B1(new_n335), .B2(new_n338), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT67), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n261), .A2(new_n226), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n258), .B1(G150), .B2(new_n255), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT66), .ZN(new_n349));
  NOR3_X1   g0149(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n227), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n204), .A2(KEYINPUT66), .A3(G20), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n345), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n265), .A2(new_n201), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n264), .A2(new_n355), .B1(new_n201), .B2(new_n252), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n344), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  INV_X1    g0159(.A(new_n255), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n346), .A2(new_n259), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n351), .B2(new_n352), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT67), .B(new_n356), .C1(new_n362), .C2(new_n345), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT9), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n358), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n358), .B2(new_n363), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n343), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n348), .A2(new_n353), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n262), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT67), .B1(new_n370), .B2(new_n356), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n354), .A2(new_n357), .A3(new_n344), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT9), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n358), .A2(new_n363), .A3(new_n364), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n343), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n368), .A2(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n347), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n259), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n381), .A2(new_n262), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n264), .A2(G77), .A3(new_n266), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G77), .B2(new_n251), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n330), .A2(new_n326), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G238), .B1(G107), .B2(new_n330), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n274), .A2(new_n326), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n275), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n280), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n280), .A2(new_n288), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(G244), .B1(new_n288), .B2(new_n286), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n385), .B1(new_n393), .B2(new_n314), .ZN(new_n394));
  INV_X1    g0194(.A(new_n393), .ZN(new_n395));
  INV_X1    g0195(.A(G179), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n339), .A2(new_n314), .B1(new_n370), .B2(new_n356), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(G179), .B2(new_n339), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n385), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n395), .B2(G190), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n393), .A2(G200), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n378), .A2(new_n398), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n391), .A2(G232), .B1(new_n288), .B2(new_n286), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n333), .A2(new_n326), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n336), .A2(G1698), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(new_n328), .C2(new_n329), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n290), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n301), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n289), .B1(new_n275), .B2(new_n291), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT77), .B(G190), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n416), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n345), .A2(new_n251), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n346), .A2(new_n265), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(KEYINPUT76), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(KEYINPUT76), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n422), .A2(new_n423), .B1(new_n252), .B2(new_n346), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G58), .A2(G68), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT75), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT75), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(G58), .A3(G68), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n428), .A3(new_n223), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G20), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n255), .A2(G159), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT7), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n328), .A2(new_n329), .A3(new_n433), .A4(G20), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT74), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n328), .B2(new_n329), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n272), .A2(KEYINPUT74), .A3(new_n273), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n227), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n438), .B2(new_n433), .ZN(new_n439));
  OAI211_X1 g0239(.A(KEYINPUT16), .B(new_n432), .C1(new_n439), .C2(new_n203), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT16), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n433), .B1(new_n274), .B2(G20), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n330), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n203), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n430), .A2(new_n431), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n262), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n419), .B(new_n424), .C1(new_n441), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n407), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n422), .A2(new_n423), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n251), .B2(new_n347), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT7), .B1(new_n330), .B2(new_n227), .ZN(new_n454));
  OAI21_X1  g0254(.A(G68), .B1(new_n454), .B2(new_n434), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n432), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n345), .B1(new_n456), .B2(new_n442), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n453), .B1(new_n457), .B2(new_n440), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(KEYINPUT78), .A3(KEYINPUT17), .A4(new_n419), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n416), .A2(new_n413), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G179), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n314), .B2(new_n460), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT18), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n424), .B1(new_n441), .B2(new_n448), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n451), .A2(new_n459), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n270), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n316), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT72), .B1(new_n315), .B2(new_n316), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n309), .A2(G179), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n470), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n298), .A2(G200), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n300), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n298), .A2(KEYINPUT69), .A3(G200), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n470), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n312), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n310), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT73), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n477), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n325), .A2(new_n406), .A3(new_n469), .A4(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n227), .B2(G107), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n216), .A2(KEYINPUT23), .A3(G20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(G20), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n227), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT22), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT22), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n274), .A2(new_n497), .A3(new_n227), .A4(G87), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT24), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n345), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n498), .ZN(new_n504));
  INV_X1    g0304(.A(new_n494), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT85), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n499), .A2(new_n500), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT24), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT25), .B1(new_n252), .B2(new_n216), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n216), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n250), .A2(G33), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n345), .A2(new_n251), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n216), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G294), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n388), .C2(new_n211), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n250), .A2(G45), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT5), .B(G41), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n280), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n522), .A2(new_n280), .B1(G264), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n286), .A2(new_n524), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g0328(.A(G169), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n531), .B2(new_n396), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n519), .A2(new_n532), .A3(KEYINPUT86), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT86), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n527), .A2(new_n396), .A3(new_n528), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n531), .B2(G169), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n517), .B1(new_n503), .B2(new_n509), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n531), .A2(G190), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n530), .A2(G200), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n533), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT6), .ZN(new_n543));
  INV_X1    g0343(.A(G97), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n543), .A2(new_n544), .A3(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(G97), .B(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n227), .B1(new_n214), .B2(new_n360), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n216), .B1(new_n443), .B2(new_n444), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n262), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  MUX2_X1   g0350(.A(new_n251), .B(new_n516), .S(G97), .Z(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n274), .A2(G244), .A3(new_n326), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n326), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n290), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n526), .A2(G257), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n528), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n562), .A2(new_n396), .A3(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n553), .A2(new_n554), .B1(G33), .B2(G283), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT81), .B1(new_n386), .B2(G250), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n559), .A2(new_n560), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n566), .B(new_n557), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n280), .ZN(new_n570));
  INV_X1    g0370(.A(new_n564), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n314), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n552), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(G200), .B1(new_n562), .B2(new_n564), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(G190), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT80), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n550), .A2(new_n577), .A3(new_n551), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G116), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n252), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n264), .A2(G116), .A3(new_n515), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n556), .B(new_n227), .C1(G33), .C2(new_n544), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(new_n262), .C1(new_n227), .C2(G116), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n582), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n525), .A2(new_n524), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(G270), .A3(new_n290), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n528), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n274), .A2(G257), .A3(new_n326), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n330), .A2(G303), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(new_n332), .C2(new_n217), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n280), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n417), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n589), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n301), .B2(new_n596), .ZN(new_n599));
  INV_X1    g0399(.A(new_n592), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n280), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n589), .A3(G169), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n600), .A2(new_n601), .A3(G179), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n589), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n602), .A2(new_n589), .A3(KEYINPUT21), .A4(G169), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n599), .A2(new_n605), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT19), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n259), .B2(new_n544), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n274), .A2(new_n227), .A3(G68), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n210), .A2(new_n544), .A3(new_n216), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n210), .A2(new_n544), .A3(new_n216), .A4(KEYINPUT82), .ZN(new_n618));
  NAND3_X1  g0418(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n617), .A2(new_n618), .B1(new_n227), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n262), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n380), .A2(new_n252), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n380), .C2(new_n516), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n215), .A2(G1698), .ZN(new_n624));
  OAI221_X1 g0424(.A(new_n624), .B1(G238), .B2(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n290), .B1(new_n625), .B2(new_n493), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n290), .A2(G250), .A3(new_n523), .ZN(new_n627));
  INV_X1    g0427(.A(new_n286), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n628), .B2(new_n523), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n314), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n626), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n396), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n623), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(G200), .B1(new_n626), .B2(new_n629), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT83), .B1(new_n516), .B2(new_n210), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT83), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n264), .A2(new_n636), .A3(G87), .A4(new_n515), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n634), .A2(new_n638), .A3(new_n621), .A4(new_n622), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n631), .A2(G190), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n633), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n580), .A2(new_n610), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n488), .A2(new_n542), .A3(new_n645), .ZN(G372));
  OR2_X1    g0446(.A1(new_n634), .A2(KEYINPUT87), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n634), .A2(KEYINPUT87), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n638), .A2(new_n621), .A3(new_n622), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n633), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n519), .A2(new_n532), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n608), .A2(new_n609), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(new_n605), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n654), .A2(new_n657), .A3(new_n573), .A4(new_n579), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n564), .B1(new_n569), .B2(new_n280), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G179), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n314), .B2(new_n659), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT88), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n661), .A2(KEYINPUT88), .B1(new_n576), .B2(new_n578), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  INV_X1    g0464(.A(new_n633), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n649), .B2(new_n650), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n644), .A2(new_n573), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n665), .B1(new_n668), .B2(KEYINPUT26), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n658), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n488), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n464), .A2(new_n467), .ZN(new_n672));
  INV_X1    g0472(.A(new_n398), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n324), .B1(new_n483), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n451), .A2(new_n459), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n367), .A2(KEYINPUT10), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n376), .B1(new_n375), .B2(new_n343), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n368), .A2(new_n377), .A3(KEYINPUT89), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n401), .B1(new_n676), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n671), .A2(new_n683), .ZN(G369));
  NAND2_X1  g0484(.A1(new_n656), .A2(new_n605), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n250), .A2(new_n227), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n589), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT90), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n610), .B2(new_n693), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n519), .A2(new_n691), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n542), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n655), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n691), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n691), .B1(new_n656), .B2(new_n605), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n542), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n691), .B(KEYINPUT91), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(G399));
  NAND3_X1  g0512(.A1(new_n617), .A2(new_n581), .A3(new_n618), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n230), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(G1), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n224), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT92), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n570), .A2(new_n571), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n596), .A2(G179), .A3(new_n527), .A4(new_n631), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT30), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n527), .A2(new_n631), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n606), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n659), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT93), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n396), .B1(new_n626), .B2(new_n629), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n596), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n731), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n602), .A2(new_n733), .A3(KEYINPUT93), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n531), .A2(new_n659), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n725), .A2(new_n729), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n691), .B1(new_n737), .B2(KEYINPUT94), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n735), .A2(new_n736), .ZN(new_n739));
  INV_X1    g0539(.A(new_n729), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n728), .B1(new_n727), .B2(new_n659), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT94), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n722), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n645), .A2(new_n542), .A3(new_n708), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n697), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n662), .A2(new_n663), .A3(KEYINPUT26), .A4(new_n666), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT96), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n652), .A2(new_n580), .A3(new_n653), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n533), .A2(new_n538), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(new_n755), .B2(new_n685), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n668), .A2(new_n664), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n751), .A3(new_n752), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n753), .A2(new_n756), .A3(new_n758), .A4(new_n633), .ZN(new_n759));
  INV_X1    g0559(.A(new_n691), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(KEYINPUT29), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n670), .A2(new_n708), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT95), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT29), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n750), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n721), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n695), .A2(G330), .ZN(new_n771));
  INV_X1    g0571(.A(G13), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n250), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n716), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n698), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT97), .Z(new_n778));
  AOI21_X1  g0578(.A(new_n226), .B1(G20), .B2(new_n314), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n227), .B1(new_n781), .B2(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n544), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n227), .A2(G179), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n340), .A3(G200), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n274), .B1(new_n785), .B2(new_n216), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n227), .A2(new_n396), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n417), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n783), .B(new_n786), .C1(G50), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n301), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G190), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G68), .A2(new_n791), .B1(new_n793), .B2(G77), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n210), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n792), .A2(new_n417), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(new_n797), .B2(G58), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n781), .A2(G20), .A3(new_n340), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n790), .A2(new_n794), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n782), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n799), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n274), .B(new_n805), .C1(G329), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  INV_X1    g0608(.A(new_n785), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n791), .A2(new_n808), .B1(new_n809), .B2(G283), .ZN(new_n810));
  INV_X1    g0610(.A(new_n795), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n797), .A2(G322), .B1(new_n811), .B2(G303), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n789), .A2(G326), .B1(new_n793), .B2(G311), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n807), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n780), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n274), .A2(new_n230), .ZN(new_n816));
  INV_X1    g0616(.A(G355), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(G116), .B2(new_n230), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n436), .A2(new_n437), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n715), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G45), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n225), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n245), .A2(new_n822), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G13), .A2(G33), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n227), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT98), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n779), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n776), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n815), .B(new_n832), .C1(new_n696), .C2(new_n829), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT99), .Z(new_n834));
  NAND2_X1  g0634(.A1(new_n778), .A2(new_n834), .ZN(G396));
  NAND2_X1  g0635(.A1(new_n673), .A2(new_n760), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n403), .A2(new_n404), .B1(new_n402), .B2(new_n691), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n673), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n762), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n838), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n670), .A2(new_n708), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n776), .B1(new_n750), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n750), .B2(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(new_n776), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n779), .A2(new_n826), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n214), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n819), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n811), .A2(G50), .B1(new_n809), .B2(G68), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n202), .B2(new_n782), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n848), .B(new_n850), .C1(G132), .C2(new_n806), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT101), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n797), .A2(G143), .B1(new_n791), .B2(G150), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n789), .A2(G137), .B1(new_n793), .B2(G159), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT34), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n851), .A2(new_n852), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G116), .A2(new_n793), .B1(new_n791), .B2(G283), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT100), .Z(new_n861));
  AOI211_X1 g0661(.A(new_n274), .B(new_n783), .C1(G311), .C2(new_n806), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n797), .A2(G294), .B1(new_n811), .B2(G107), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n789), .A2(G303), .B1(new_n809), .B2(G87), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n826), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n847), .B1(new_n780), .B2(new_n866), .C1(new_n840), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n844), .A2(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n773), .A2(new_n250), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n438), .A2(new_n433), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n444), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n446), .B1(new_n872), .B2(G68), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n262), .B1(new_n873), .B2(KEYINPUT16), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT103), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n432), .B1(new_n439), .B2(new_n203), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n345), .B1(new_n877), .B2(new_n442), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n441), .B1(new_n878), .B2(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n689), .B1(new_n880), .B2(new_n424), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n468), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  OAI211_X1 g0683(.A(KEYINPUT103), .B(new_n262), .C1(new_n873), .C2(KEYINPUT16), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n440), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n878), .A2(KEYINPUT103), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n424), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n689), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n462), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n883), .B1(new_n891), .B2(new_n449), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n449), .B1(new_n458), .B2(new_n463), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n458), .A2(new_n689), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT37), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT38), .B(new_n882), .C1(new_n892), .C2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n468), .A2(new_n894), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n465), .A2(new_n462), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n465), .A2(new_n888), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n883), .A4(new_n449), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n896), .A2(new_n897), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n453), .B1(new_n876), .B2(new_n879), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n449), .B1(new_n908), .B2(new_n889), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n895), .B1(new_n909), .B2(KEYINPUT37), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n468), .A2(new_n881), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n897), .B1(new_n912), .B2(new_n896), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT104), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT105), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n477), .A2(new_n691), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n910), .A2(new_n911), .A3(new_n905), .ZN(new_n920));
  INV_X1    g0720(.A(new_n449), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n887), .B2(new_n890), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n902), .B1(new_n922), .B2(new_n883), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n923), .B2(new_n882), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT39), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n896), .A2(new_n906), .A3(new_n897), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(KEYINPUT104), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT105), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(new_n916), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n918), .A2(new_n919), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n672), .A2(new_n888), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n270), .A2(new_n760), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n324), .B2(new_n313), .ZN(new_n933));
  INV_X1    g0733(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n477), .A2(new_n483), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n836), .B(KEYINPUT102), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n841), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n912), .A2(new_n896), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n931), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n930), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n762), .A2(new_n764), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT95), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n488), .A2(new_n944), .A3(new_n765), .A4(new_n761), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n683), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n942), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT94), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n745), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n949), .A2(KEYINPUT31), .A3(new_n691), .A4(new_n742), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n744), .A2(new_n748), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n488), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n896), .A2(new_n906), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n838), .B1(new_n933), .B2(new_n935), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n951), .A2(new_n954), .A3(KEYINPUT40), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n940), .A2(new_n951), .A3(new_n954), .ZN(new_n956));
  XNOR2_X1  g0756(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n953), .A2(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n697), .B1(new_n952), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n952), .B2(new_n958), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n870), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n947), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(new_n547), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT35), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT35), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n964), .A2(G116), .A3(new_n228), .A4(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n225), .A2(G77), .A3(new_n428), .A4(new_n426), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(G50), .B2(new_n203), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n772), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n967), .A3(new_n970), .ZN(G367));
  OAI21_X1  g0771(.A(new_n830), .B1(new_n230), .B2(new_n380), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n821), .A2(new_n241), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n776), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n785), .A2(new_n214), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n330), .B(new_n975), .C1(G137), .C2(new_n806), .ZN(new_n976));
  INV_X1    g0776(.A(new_n782), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n811), .A2(G58), .B1(new_n977), .B2(G68), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n797), .A2(G150), .B1(new_n793), .B2(G50), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n789), .A2(G143), .B1(new_n791), .B2(G159), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n976), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n789), .A2(G311), .ZN(new_n982));
  INV_X1    g0782(.A(new_n793), .ZN(new_n983));
  INV_X1    g0783(.A(G283), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n797), .ZN(new_n986));
  INV_X1    g0786(.A(G303), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n986), .A2(new_n987), .B1(new_n216), .B2(new_n782), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n985), .B(new_n988), .C1(G294), .C2(new_n791), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT110), .B1(new_n811), .B2(G116), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n848), .B1(new_n544), .B2(new_n785), .C1(new_n993), .C2(new_n799), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT111), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n981), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n974), .B1(new_n998), .B2(new_n779), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n650), .A2(new_n760), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n666), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT107), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1000), .A2(new_n633), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(KEYINPUT107), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n999), .B1(new_n1006), .B2(new_n828), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n716), .B(KEYINPUT41), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n705), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n700), .A2(new_n702), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n706), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n698), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n750), .C1(new_n766), .C2(new_n767), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n708), .B1(new_n576), .B2(new_n578), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n580), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n662), .A2(new_n663), .A3(new_n707), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT108), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT108), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n1023), .A2(KEYINPUT45), .A3(new_n711), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT45), .B1(new_n1023), .B2(new_n711), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1020), .A2(new_n710), .A3(new_n1022), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT44), .Z(new_n1028));
  INV_X1    g0828(.A(KEYINPUT109), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n704), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n698), .A2(KEYINPUT109), .A3(new_n703), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1026), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1027), .B(KEYINPUT44), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1029), .B(new_n704), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1015), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1010), .B1(new_n1036), .B2(new_n768), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n774), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1006), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT43), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1021), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n542), .B(new_n705), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT42), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1023), .A2(new_n755), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n707), .B1(new_n1047), .B2(new_n573), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1041), .B(new_n1042), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1048), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT42), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1045), .B(new_n1051), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1050), .A2(new_n1052), .A3(new_n1040), .A4(new_n1039), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1023), .A2(new_n698), .A3(new_n703), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1055), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1049), .A2(new_n1053), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1008), .B1(new_n1038), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(G387));
  NAND3_X1  g0862(.A1(new_n700), .A2(new_n702), .A3(new_n829), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n820), .B1(new_n238), .B2(new_n822), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n714), .B2(new_n816), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n346), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1066));
  OAI21_X1  g0866(.A(KEYINPUT50), .B1(new_n346), .B2(G50), .ZN(new_n1067));
  AOI21_X1  g0867(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n714), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1065), .A2(new_n1069), .B1(new_n216), .B2(new_n715), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n776), .B1(new_n1070), .B2(new_n831), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n986), .A2(new_n201), .B1(new_n983), .B2(new_n203), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n347), .B2(new_n791), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n848), .B1(G150), .B2(new_n806), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n380), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n809), .A2(G97), .B1(new_n977), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n789), .A2(G159), .B1(new_n811), .B2(G77), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n819), .B1(G326), .B2(new_n806), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n795), .A2(new_n804), .B1(new_n782), .B2(new_n984), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G303), .A2(new_n793), .B1(new_n791), .B2(G311), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n789), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT113), .B(G322), .Z(new_n1083));
  OAI221_X1 g0883(.A(new_n1081), .B1(new_n993), .B2(new_n986), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT48), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1080), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT49), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1079), .B1(new_n581), .B2(new_n785), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1078), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1071), .B1(new_n1091), .B2(new_n779), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1014), .A2(new_n775), .B1(new_n1063), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1015), .A2(KEYINPUT114), .A3(new_n716), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n769), .B2(new_n1014), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT114), .B1(new_n1015), .B2(new_n716), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(G393));
  INV_X1    g0897(.A(KEYINPUT117), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1036), .A2(new_n717), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1032), .A2(new_n1035), .A3(new_n1015), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT116), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1098), .B(new_n1099), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1023), .A2(new_n828), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n248), .A2(new_n820), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n830), .B1(new_n544), .B2(new_n230), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n795), .A2(new_n203), .B1(new_n782), .B2(new_n214), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n848), .B1(G143), .B2(new_n806), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(new_n210), .B2(new_n785), .C1(new_n346), .C2(new_n983), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1108), .B(new_n1110), .C1(G50), .C2(new_n791), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G150), .A2(new_n789), .B1(new_n797), .B2(G159), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT51), .Z(new_n1113));
  AOI22_X1  g0913(.A1(G311), .A2(new_n797), .B1(new_n789), .B2(G317), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT52), .Z(new_n1115));
  OAI22_X1  g0915(.A1(new_n983), .A2(new_n804), .B1(new_n581), .B2(new_n782), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n791), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1117), .A2(new_n987), .B1(new_n984), .B2(new_n795), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n330), .B1(new_n785), .B2(new_n216), .C1(new_n799), .C2(new_n1083), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1111), .A2(new_n1113), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n776), .B1(new_n1106), .B2(new_n1107), .C1(new_n1121), .C2(new_n780), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1105), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT115), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n774), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1032), .A2(new_n1035), .A3(KEYINPUT115), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1104), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1100), .B(new_n1101), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1098), .B1(new_n1129), .B2(new_n1099), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT118), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT118), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n1104), .A4(new_n1127), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1131), .A2(new_n1135), .ZN(G390));
  AND2_X1   g0936(.A1(new_n951), .A2(G330), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1137), .A2(new_n954), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n939), .A2(new_n919), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n918), .B2(new_n929), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n919), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n953), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n759), .B(new_n760), .C1(new_n673), .C2(new_n837), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n836), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n1144), .B2(new_n936), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1138), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n927), .A2(new_n928), .A3(new_n916), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n928), .B1(new_n927), .B2(new_n916), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1147), .A2(new_n1148), .B1(new_n919), .B2(new_n939), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1145), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n749), .A2(new_n840), .A3(new_n936), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1146), .A2(new_n775), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n826), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n274), .B(new_n796), .C1(G294), .C2(new_n806), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n797), .A2(G116), .B1(new_n791), .B2(G107), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n789), .A2(G283), .B1(new_n793), .B2(G97), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n809), .A2(G68), .B1(new_n977), .B2(G77), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n791), .A2(G137), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n800), .B2(new_n782), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G50), .B2(new_n809), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n330), .B1(new_n806), .B2(G125), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n983), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n811), .A2(G150), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(KEYINPUT53), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1162), .B(new_n1167), .C1(KEYINPUT53), .C2(new_n1166), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G128), .A2(new_n789), .B1(new_n797), .B2(G132), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT119), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1159), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n779), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n845), .B1(new_n346), .B2(new_n846), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1154), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1153), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n488), .A2(new_n1137), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n945), .A2(new_n683), .A3(new_n1177), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1143), .A2(new_n836), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1137), .A2(new_n840), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1151), .C1(new_n936), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n841), .A2(new_n938), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n936), .B1(new_n749), .B2(new_n840), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n1138), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1178), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n717), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1146), .A2(new_n1152), .A3(new_n1185), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1175), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G378));
  INV_X1    g0990(.A(KEYINPUT122), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n368), .A2(KEYINPUT89), .A3(new_n377), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT89), .B1(new_n368), .B2(new_n377), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n400), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n689), .B1(new_n358), .B2(new_n363), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n682), .A2(new_n400), .A3(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1191), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1199), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(KEYINPUT122), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(G330), .A3(new_n958), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n955), .A2(new_n953), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n956), .A2(new_n957), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(G330), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1209), .A2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1147), .A2(new_n1148), .A3(new_n1141), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n941), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n930), .A2(new_n941), .A3(new_n1209), .A4(new_n1214), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n775), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n845), .B1(new_n201), .B2(new_n846), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n819), .A2(G41), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n986), .A2(new_n216), .B1(new_n983), .B2(new_n380), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1117), .A2(new_n544), .B1(new_n202), .B2(new_n785), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n977), .A2(G68), .B1(new_n806), .B2(G283), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n789), .A2(G116), .B1(new_n811), .B2(G77), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1228), .A2(new_n1223), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT58), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1225), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G33), .A2(G41), .ZN(new_n1235));
  INV_X1    g1035(.A(G124), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n799), .B2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G125), .A2(new_n789), .B1(new_n797), .B2(G128), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n793), .A2(G137), .B1(G150), .B2(new_n977), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1164), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n791), .A2(G132), .B1(new_n811), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1243));
  XNOR2_X1  g1043(.A(new_n1242), .B(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT121), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1237), .B(new_n1246), .C1(G159), .C2(new_n809), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1234), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1222), .B1(new_n780), .B2(new_n1249), .C1(new_n1208), .C2(new_n867), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1221), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1178), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1188), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1215), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1255), .A2(KEYINPUT123), .A3(new_n930), .A4(new_n941), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT123), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1218), .A2(new_n1257), .A3(new_n1219), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(KEYINPUT57), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1188), .A2(new_n1253), .B1(new_n1219), .B2(new_n1218), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n716), .B1(new_n1261), .B2(KEYINPUT57), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1252), .B1(new_n1260), .B2(new_n1262), .ZN(G375));
  NAND3_X1  g1063(.A1(new_n1181), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1186), .A2(new_n1010), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n937), .A2(new_n826), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n983), .A2(new_n359), .B1(new_n201), .B2(new_n782), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G159), .B2(new_n811), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n848), .B1(G128), .B2(new_n806), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n797), .A2(G137), .B1(new_n809), .B2(G58), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n789), .A2(G132), .B1(new_n791), .B2(new_n1240), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n274), .B(new_n975), .C1(G303), .C2(new_n806), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n797), .A2(G283), .B1(new_n791), .B2(G116), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n789), .A2(G294), .B1(new_n793), .B2(G107), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n811), .A2(G97), .B1(new_n977), .B2(new_n1075), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n780), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n845), .B(new_n1279), .C1(new_n203), .C2(new_n846), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1266), .A2(new_n775), .B1(new_n1267), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1265), .A2(new_n1281), .ZN(G381));
  NOR2_X1   g1082(.A1(G375), .A2(G378), .ZN(new_n1283));
  INV_X1    g1083(.A(G396), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1093), .B(new_n1284), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(G387), .A2(G384), .A3(G381), .A4(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1135), .A3(new_n1131), .A4(new_n1286), .ZN(G407));
  INV_X1    g1087(.A(new_n1283), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G343), .C2(new_n1288), .ZN(G409));
  NAND2_X1  g1089(.A1(new_n690), .A2(G213), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1281), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1266), .A2(new_n1253), .A3(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1293), .A2(new_n717), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1264), .B1(new_n1185), .B2(new_n1292), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1291), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  OR2_X1    g1096(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1254), .A2(new_n1220), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT57), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n717), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n1189), .B(new_n1251), .C1(new_n1306), .C2(new_n1259), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1258), .A2(new_n775), .A3(new_n1256), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1250), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1309), .A2(KEYINPUT124), .B1(new_n1010), .B2(new_n1261), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT124), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1308), .A2(new_n1311), .A3(new_n1250), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G378), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1290), .B(new_n1303), .C1(new_n1307), .C2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT62), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1290), .B1(new_n1307), .B2(new_n1313), .ZN(new_n1316));
  INV_X1    g1116(.A(G2897), .ZN(new_n1317));
  OAI22_X1  g1117(.A1(new_n1299), .A2(new_n1302), .B1(new_n1317), .B2(new_n1290), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1290), .A2(new_n1317), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1298), .B(new_n1319), .C1(new_n1296), .C2(new_n1301), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1316), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1309), .A2(KEYINPUT124), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1261), .A2(new_n1010), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1312), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1189), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G378), .B(new_n1252), .C1(new_n1260), .C2(new_n1262), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1290), .A4(new_n1303), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1315), .A2(new_n1322), .A3(new_n1323), .A4(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G393), .A2(G396), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1285), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1061), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1059), .B1(new_n1037), .B2(new_n774), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1285), .B(new_n1333), .C1(new_n1336), .C2(new_n1008), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1338), .A2(new_n1135), .A3(new_n1131), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1135), .B2(new_n1131), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1332), .A2(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1323), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1343));
  XOR2_X1   g1143(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1344));
  AOI21_X1  g1144(.A(new_n1343), .B1(new_n1314), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT127), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1316), .A2(new_n1346), .A3(new_n1321), .ZN(new_n1347));
  AOI22_X1  g1147(.A1(new_n1327), .A2(new_n1328), .B1(G213), .B2(new_n690), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1321), .ZN(new_n1349));
  OAI21_X1  g1149(.A(KEYINPUT127), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1348), .A2(KEYINPUT63), .A3(new_n1303), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1345), .A2(new_n1347), .A3(new_n1350), .A4(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1342), .A2(new_n1352), .ZN(G405));
  AND2_X1   g1153(.A1(G375), .A2(new_n1189), .ZN(new_n1354));
  OR3_X1    g1154(.A1(new_n1354), .A2(new_n1307), .A3(new_n1303), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1303), .B1(new_n1354), .B2(new_n1307), .ZN(new_n1356));
  AND3_X1   g1156(.A1(new_n1355), .A2(new_n1341), .A3(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1341), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1357), .A2(new_n1358), .ZN(G402));
endmodule


