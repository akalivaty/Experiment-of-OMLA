

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U320 ( .A(n323), .B(KEYINPUT13), .ZN(n373) );
  XOR2_X1 U321 ( .A(n402), .B(n401), .Z(n505) );
  XOR2_X1 U322 ( .A(n329), .B(n328), .Z(n288) );
  AND2_X1 U323 ( .A1(n561), .A2(n444), .ZN(n445) );
  XNOR2_X1 U324 ( .A(n330), .B(n288), .ZN(n331) );
  INV_X1 U325 ( .A(n373), .ZN(n374) );
  XNOR2_X1 U326 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U327 ( .A(KEYINPUT41), .B(n338), .Z(n524) );
  XOR2_X1 U328 ( .A(n305), .B(n389), .Z(n516) );
  XNOR2_X1 U329 ( .A(n448), .B(G190GAT), .ZN(n449) );
  XNOR2_X1 U330 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(G71GAT), .B(G176GAT), .Z(n290) );
  XNOR2_X1 U332 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n301) );
  XOR2_X1 U334 ( .A(G99GAT), .B(KEYINPUT20), .Z(n292) );
  XNOR2_X1 U335 ( .A(G43GAT), .B(KEYINPUT84), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n294) );
  XNOR2_X1 U337 ( .A(G134GAT), .B(G127GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n293), .B(KEYINPUT0), .ZN(n435) );
  XOR2_X1 U339 ( .A(n294), .B(n435), .Z(n299) );
  XOR2_X1 U340 ( .A(G120GAT), .B(G15GAT), .Z(n296) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(n297), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U346 ( .A(KEYINPUT17), .B(G190GAT), .Z(n303) );
  XNOR2_X1 U347 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U349 ( .A(KEYINPUT19), .B(n304), .Z(n389) );
  XOR2_X1 U350 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n388) );
  XOR2_X1 U351 ( .A(G43GAT), .B(G29GAT), .Z(n307) );
  XNOR2_X1 U352 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U354 ( .A(n308), .B(KEYINPUT69), .Z(n310) );
  XNOR2_X1 U355 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n345) );
  XOR2_X1 U357 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n312) );
  NAND2_X1 U358 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U360 ( .A(n313), .B(KEYINPUT30), .Z(n317) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(G113GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n314), .B(G1GAT), .ZN(n441) );
  XNOR2_X1 U363 ( .A(G22GAT), .B(G15GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n315), .B(KEYINPUT70), .ZN(n372) );
  XNOR2_X1 U365 ( .A(n441), .B(n372), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U367 ( .A(G169GAT), .B(G8GAT), .Z(n396) );
  XOR2_X1 U368 ( .A(n318), .B(n396), .Z(n320) );
  XNOR2_X1 U369 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U371 ( .A(n345), .B(n321), .Z(n564) );
  XNOR2_X1 U372 ( .A(G120GAT), .B(G148GAT), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n322), .B(G57GAT), .ZN(n440) );
  XOR2_X1 U374 ( .A(G71GAT), .B(KEYINPUT72), .Z(n323) );
  XNOR2_X1 U375 ( .A(n440), .B(n373), .ZN(n332) );
  XOR2_X1 U376 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n325) );
  NAND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n327) );
  XNOR2_X1 U379 ( .A(G176GAT), .B(G92GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n326), .B(G64GAT), .ZN(n392) );
  XNOR2_X1 U381 ( .A(n327), .B(n392), .ZN(n330) );
  XOR2_X1 U382 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n329) );
  XNOR2_X1 U383 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n328) );
  XNOR2_X1 U384 ( .A(G106GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n333), .B(G204GAT), .ZN(n413) );
  XNOR2_X1 U386 ( .A(G99GAT), .B(G85GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n334), .B(KEYINPUT75), .ZN(n348) );
  XNOR2_X1 U388 ( .A(n413), .B(n348), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n570) );
  INV_X1 U390 ( .A(KEYINPUT64), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n570), .B(n337), .ZN(n338) );
  INV_X1 U392 ( .A(n524), .ZN(n555) );
  NAND2_X1 U393 ( .A1(n564), .A2(n555), .ZN(n339) );
  OR2_X1 U394 ( .A1(KEYINPUT46), .A2(n339), .ZN(n341) );
  NAND2_X1 U395 ( .A1(KEYINPUT46), .A2(n339), .ZN(n340) );
  NAND2_X1 U396 ( .A1(n341), .A2(n340), .ZN(n379) );
  XOR2_X1 U397 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n343) );
  XNOR2_X1 U398 ( .A(KEYINPUT78), .B(KEYINPUT9), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n358) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(KEYINPUT79), .Z(n347) );
  XNOR2_X1 U402 ( .A(G190GAT), .B(G218GAT), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n356) );
  XOR2_X1 U404 ( .A(KEYINPUT80), .B(n348), .Z(n350) );
  NAND2_X1 U405 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U407 ( .A(G92GAT), .B(G106GAT), .Z(n352) );
  XNOR2_X1 U408 ( .A(G134GAT), .B(G162GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(n354), .B(n353), .Z(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(n358), .B(n357), .Z(n531) );
  XOR2_X1 U413 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n360) );
  XNOR2_X1 U414 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n368) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XOR2_X1 U417 ( .A(G57GAT), .B(G78GAT), .Z(n362) );
  XNOR2_X1 U418 ( .A(G183GAT), .B(G127GAT), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U420 ( .A(G155GAT), .B(G211GAT), .Z(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n377) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U425 ( .A(G1GAT), .B(G8GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n375) );
  XOR2_X1 U428 ( .A(n375), .B(n374), .Z(n376) );
  XOR2_X1 U429 ( .A(n377), .B(n376), .Z(n573) );
  INV_X1 U430 ( .A(n573), .ZN(n527) );
  AND2_X1 U431 ( .A1(n531), .A2(n527), .ZN(n378) );
  AND2_X1 U432 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n380), .B(KEYINPUT47), .ZN(n386) );
  XOR2_X1 U434 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n382) );
  XOR2_X1 U435 ( .A(KEYINPUT36), .B(n531), .Z(n576) );
  NAND2_X1 U436 ( .A1(n576), .A2(n573), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  NOR2_X1 U438 ( .A1(n570), .A2(n383), .ZN(n384) );
  XOR2_X1 U439 ( .A(n564), .B(KEYINPUT71), .Z(n550) );
  INV_X1 U440 ( .A(n550), .ZN(n520) );
  NAND2_X1 U441 ( .A1(n384), .A2(n520), .ZN(n385) );
  AND2_X1 U442 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n534) );
  INV_X1 U444 ( .A(n389), .ZN(n402) );
  XOR2_X1 U445 ( .A(G211GAT), .B(KEYINPUT21), .Z(n391) );
  XNOR2_X1 U446 ( .A(G197GAT), .B(G218GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n415) );
  XNOR2_X1 U448 ( .A(n415), .B(n392), .ZN(n400) );
  XOR2_X1 U449 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n394) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(G204GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U452 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  NOR2_X1 U456 ( .A1(n534), .A2(n505), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n403), .B(KEYINPUT54), .ZN(n561) );
  XNOR2_X1 U458 ( .A(KEYINPUT87), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(KEYINPUT88), .ZN(n405) );
  XOR2_X1 U460 ( .A(n405), .B(KEYINPUT2), .Z(n407) );
  XNOR2_X1 U461 ( .A(G155GAT), .B(G162GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n432) );
  XOR2_X1 U463 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n409) );
  XNOR2_X1 U464 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U466 ( .A(G50GAT), .B(KEYINPUT23), .Z(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n419) );
  XNOR2_X1 U468 ( .A(G22GAT), .B(KEYINPUT89), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n412), .B(G148GAT), .ZN(n414) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n417) );
  XNOR2_X1 U471 ( .A(G141GAT), .B(n415), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n421) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n432), .B(n422), .ZN(n461) );
  XOR2_X1 U477 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n426) );
  XNOR2_X1 U481 ( .A(G29GAT), .B(G85GAT), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U483 ( .A(n428), .B(n427), .Z(n434) );
  XOR2_X1 U484 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n430) );
  XNOR2_X1 U485 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n439) );
  XOR2_X1 U489 ( .A(KEYINPUT96), .B(n435), .Z(n437) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n460) );
  XNOR2_X1 U495 ( .A(KEYINPUT97), .B(n460), .ZN(n463) );
  NOR2_X1 U496 ( .A1(n461), .A2(n463), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NOR2_X1 U498 ( .A1(n516), .A2(n446), .ZN(n447) );
  XNOR2_X1 U499 ( .A(KEYINPUT120), .B(n447), .ZN(n558) );
  INV_X1 U500 ( .A(n531), .ZN(n546) );
  NAND2_X1 U501 ( .A1(n558), .A2(n546), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n448) );
  INV_X1 U503 ( .A(n463), .ZN(n560) );
  NOR2_X1 U504 ( .A1(n570), .A2(n520), .ZN(n451) );
  XOR2_X1 U505 ( .A(KEYINPUT77), .B(n451), .Z(n483) );
  NOR2_X1 U506 ( .A1(n516), .A2(n505), .ZN(n452) );
  NOR2_X1 U507 ( .A1(n461), .A2(n452), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT25), .ZN(n458) );
  XOR2_X1 U509 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n455) );
  NAND2_X1 U510 ( .A1(n461), .A2(n516), .ZN(n454) );
  XOR2_X1 U511 ( .A(n455), .B(n454), .Z(n562) );
  INV_X1 U512 ( .A(n562), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(n505), .Z(n462) );
  NAND2_X1 U514 ( .A1(n456), .A2(n462), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n458), .A2(n457), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n460), .A2(n459), .ZN(n466) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(n461), .Z(n513) );
  INV_X1 U518 ( .A(n513), .ZN(n464) );
  NAND2_X1 U519 ( .A1(n463), .A2(n462), .ZN(n536) );
  NOR2_X1 U520 ( .A1(n464), .A2(n536), .ZN(n518) );
  NAND2_X1 U521 ( .A1(n518), .A2(n516), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n479) );
  NAND2_X1 U523 ( .A1(n531), .A2(n573), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(n467), .Z(n468) );
  AND2_X1 U525 ( .A1(n479), .A2(n468), .ZN(n493) );
  NAND2_X1 U526 ( .A1(n483), .A2(n493), .ZN(n475) );
  NOR2_X1 U527 ( .A1(n560), .A2(n475), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT34), .B(n469), .Z(n470) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n470), .ZN(G1324GAT) );
  NOR2_X1 U530 ( .A1(n505), .A2(n475), .ZN(n472) );
  XNOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(G1325GAT) );
  NOR2_X1 U533 ( .A1(n516), .A2(n475), .ZN(n474) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NOR2_X1 U536 ( .A1(n513), .A2(n475), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT102), .B(n476), .Z(n477) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(n477), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT104), .Z(n478) );
  XNOR2_X1 U540 ( .A(KEYINPUT39), .B(n478), .ZN(n486) );
  NAND2_X1 U541 ( .A1(n527), .A2(n479), .ZN(n480) );
  XNOR2_X1 U542 ( .A(KEYINPUT103), .B(n480), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n481), .A2(n576), .ZN(n482) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n482), .ZN(n503) );
  NAND2_X1 U545 ( .A1(n483), .A2(n503), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(KEYINPUT38), .ZN(n491) );
  NOR2_X1 U547 ( .A1(n560), .A2(n491), .ZN(n485) );
  XOR2_X1 U548 ( .A(n486), .B(n485), .Z(G1328GAT) );
  NOR2_X1 U549 ( .A1(n491), .A2(n505), .ZN(n487) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n487), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n491), .A2(n516), .ZN(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n491), .A2(n513), .ZN(n492) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n492), .Z(G1331GAT) );
  NOR2_X1 U557 ( .A1(n564), .A2(n524), .ZN(n502) );
  NAND2_X1 U558 ( .A1(n502), .A2(n493), .ZN(n499) );
  NOR2_X1 U559 ( .A1(n560), .A2(n499), .ZN(n495) );
  XNOR2_X1 U560 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n494) );
  XNOR2_X1 U561 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n496), .Z(G1332GAT) );
  NOR2_X1 U563 ( .A1(n505), .A2(n499), .ZN(n497) );
  XOR2_X1 U564 ( .A(G64GAT), .B(n497), .Z(G1333GAT) );
  NOR2_X1 U565 ( .A1(n516), .A2(n499), .ZN(n498) );
  XOR2_X1 U566 ( .A(G71GAT), .B(n498), .Z(G1334GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n499), .ZN(n501) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(G1335GAT) );
  NAND2_X1 U570 ( .A1(n503), .A2(n502), .ZN(n512) );
  NOR2_X1 U571 ( .A1(n560), .A2(n512), .ZN(n504) );
  XOR2_X1 U572 ( .A(G85GAT), .B(n504), .Z(G1336GAT) );
  NOR2_X1 U573 ( .A1(n505), .A2(n512), .ZN(n507) );
  XNOR2_X1 U574 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(G1337GAT) );
  NOR2_X1 U576 ( .A1(n516), .A2(n512), .ZN(n508) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(n508), .Z(n509) );
  XNOR2_X1 U578 ( .A(G99GAT), .B(n509), .ZN(G1338GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n511) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n510) );
  XNOR2_X1 U581 ( .A(n511), .B(n510), .ZN(n515) );
  NOR2_X1 U582 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U583 ( .A(n515), .B(n514), .Z(G1339GAT) );
  NOR2_X1 U584 ( .A1(n516), .A2(n534), .ZN(n517) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(KEYINPUT112), .B(n519), .ZN(n530) );
  NOR2_X1 U587 ( .A1(n530), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n523), .ZN(G1340GAT) );
  XNOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n524), .A2(n530), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1341GAT) );
  NOR2_X1 U594 ( .A1(n527), .A2(n530), .ZN(n528) );
  XOR2_X1 U595 ( .A(KEYINPUT50), .B(n528), .Z(n529) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  XNOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n533) );
  NOR2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1343GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n538) );
  OR2_X1 U601 ( .A1(n534), .A2(n562), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n547), .A2(n564), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n541) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(KEYINPUT117), .B(n542), .Z(n544) );
  NAND2_X1 U610 ( .A1(n547), .A2(n555), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n573), .A2(n547), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U614 ( .A(G162GAT), .B(KEYINPUT119), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n558), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(n554), .Z(n557) );
  NAND2_X1 U623 ( .A1(n558), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n573), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n566) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n577) );
  NAND2_X1 U630 ( .A1(n577), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(n567), .B(KEYINPUT124), .Z(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n577), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

