//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  AOI211_X1 g0013(.A(new_n211), .B(new_n213), .C1(G77), .C2(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n220), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NOR3_X1   g0027(.A1(new_n219), .A2(new_n222), .A3(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  XNOR2_X1  g0045(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT15), .B(G87), .Z(new_n249));
  NAND2_X1  g0049(.A1(new_n216), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n247), .A2(new_n248), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(new_n216), .B2(new_n204), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n221), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n253), .A2(new_n255), .B1(new_n204), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n255), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(new_n216), .B2(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n215), .A2(KEYINPUT69), .A3(G20), .ZN(new_n262));
  AND4_X1   g0062(.A1(new_n256), .A2(new_n259), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G77), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G238), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G232), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n266), .B(new_n267), .C1(new_n268), .C2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(new_n221), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n269), .B(new_n273), .C1(G107), .C2(new_n266), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n215), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n277), .A2(new_n272), .A3(G274), .A4(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G244), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n272), .A2(new_n275), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n274), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n265), .B(new_n284), .C1(G179), .C2(new_n282), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(G200), .ZN(new_n286));
  INV_X1    g0086(.A(G190), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n282), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n265), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G58), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n209), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G58), .A2(G68), .ZN(new_n292));
  OAI21_X1  g0092(.A(G20), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n248), .A2(G159), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT7), .ZN(new_n297));
  INV_X1    g0097(.A(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT3), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G33), .ZN(new_n301));
  AOI211_X1 g0101(.A(new_n297), .B(G20), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n299), .B2(new_n301), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n216), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n306), .B2(new_n297), .ZN(new_n307));
  OAI211_X1 g0107(.A(KEYINPUT16), .B(new_n296), .C1(new_n307), .C2(new_n209), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n297), .B1(new_n266), .B2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n299), .A2(new_n301), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n209), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n313), .B2(new_n295), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT74), .B(new_n309), .C1(new_n313), .C2(new_n295), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n308), .A2(new_n316), .A3(new_n255), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G226), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G1698), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n266), .B(new_n320), .C1(G223), .C2(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G87), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n272), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n272), .A2(G232), .A3(new_n275), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n279), .A2(KEYINPUT75), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT75), .B1(new_n279), .B2(new_n325), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n324), .B(new_n287), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n328), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n323), .B1(new_n330), .B2(new_n326), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n331), .B2(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n246), .A2(new_n256), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n263), .B2(new_n246), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n318), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n318), .A2(new_n334), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n324), .B(G179), .C1(new_n327), .C2(new_n328), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n331), .B2(new_n283), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT76), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G169), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT76), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n338), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n337), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n337), .A2(new_n340), .A3(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT18), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n336), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT77), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n289), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n268), .A2(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G226), .B2(G1698), .ZN(new_n357));
  INV_X1    g0157(.A(G97), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n357), .A2(new_n311), .B1(new_n298), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n273), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n360), .A2(new_n279), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n272), .A2(G238), .A3(new_n275), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n355), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n355), .A3(new_n362), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n248), .ZN(new_n369));
  INV_X1    g0169(.A(G50), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n369), .A2(new_n370), .B1(new_n250), .B2(new_n204), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n216), .A2(G68), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n255), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT11), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n263), .A2(G68), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n374), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(new_n215), .A3(G13), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT12), .ZN(new_n379));
  AND4_X1   g0179(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n364), .A2(new_n365), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n287), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n368), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(KEYINPUT72), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n366), .B2(new_n283), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n366), .A2(G179), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n381), .B(G169), .C1(KEYINPUT72), .C2(new_n384), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n380), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n248), .A2(G150), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n392), .B1(new_n250), .B2(new_n246), .C1(new_n203), .C2(new_n216), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n255), .B1(new_n370), .B2(new_n257), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n263), .A2(G50), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT70), .B1(new_n397), .B2(KEYINPUT9), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G223), .A2(G1698), .ZN(new_n399));
  INV_X1    g0199(.A(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G222), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n266), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n273), .C1(G77), .C2(new_n266), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n279), .C1(new_n319), .C2(new_n281), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n287), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n397), .B2(KEYINPUT9), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(G200), .ZN(new_n407));
  XOR2_X1   g0207(.A(new_n407), .B(KEYINPUT71), .Z(new_n408));
  INV_X1    g0208(.A(KEYINPUT70), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT9), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n396), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n398), .A2(new_n406), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT10), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n404), .A2(new_n283), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n404), .A2(G179), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n396), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n354), .A2(new_n391), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G179), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n210), .A2(new_n400), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n280), .A2(G1698), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n299), .A2(new_n422), .A3(new_n301), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G116), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n273), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n215), .A2(G45), .ZN(new_n428));
  INV_X1    g0228(.A(new_n271), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(G250), .C1(new_n429), .C2(new_n221), .ZN(new_n430));
  INV_X1    g0230(.A(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G274), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT79), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n272), .B1(new_n424), .B2(new_n425), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT79), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n436), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n421), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n249), .A2(new_n256), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT19), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n250), .B2(new_n358), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT80), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n266), .A2(new_n216), .A3(G68), .ZN(new_n445));
  NAND3_X1  g0245(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n216), .ZN(new_n447));
  INV_X1    g0247(.A(G87), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n358), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT80), .B(new_n441), .C1(new_n250), .C2(new_n358), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n444), .A2(new_n445), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n440), .B1(new_n453), .B2(new_n255), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n215), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n256), .A2(new_n455), .A3(new_n221), .A4(new_n254), .ZN(new_n456));
  INV_X1    g0256(.A(new_n249), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n435), .A2(new_n438), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n439), .B(new_n458), .C1(new_n459), .C2(G169), .ZN(new_n460));
  OAI21_X1  g0260(.A(G190), .B1(new_n435), .B2(new_n438), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n456), .A2(new_n448), .ZN(new_n462));
  AOI211_X1 g0262(.A(new_n440), .B(new_n462), .C1(new_n453), .C2(new_n255), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n461), .B(new_n463), .C1(new_n459), .C2(new_n367), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n256), .A2(G107), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n467), .A2(KEYINPUT25), .B1(new_n456), .B2(new_n449), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT23), .ZN(new_n469));
  OAI211_X1 g0269(.A(G20), .B(new_n449), .C1(new_n469), .C2(KEYINPUT83), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n299), .A2(new_n301), .A3(new_n216), .A4(G87), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT22), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n473), .A2(new_n474), .B1(G116), .B2(new_n251), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n266), .A2(KEYINPUT22), .A3(new_n216), .A4(G87), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT24), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n472), .A2(new_n475), .A3(new_n479), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n468), .B1(new_n481), .B2(new_n255), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n467), .A2(KEYINPUT25), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT78), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(G41), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n428), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(G41), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(G274), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n266), .B1(G250), .B2(G1698), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n400), .A2(G257), .ZN(new_n494));
  INV_X1    g0294(.A(G294), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n493), .A2(new_n494), .B1(new_n298), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n273), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n487), .A2(new_n489), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n491), .A3(new_n431), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G264), .A3(new_n272), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n273), .B1(new_n490), .B2(new_n491), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT84), .B1(new_n503), .B2(G264), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n492), .B(new_n497), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n283), .ZN(new_n506));
  INV_X1    g0306(.A(new_n505), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n421), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n484), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n465), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(G200), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n500), .A2(new_n501), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n503), .A2(KEYINPUT84), .A3(G264), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(G190), .A3(new_n492), .A4(new_n497), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n482), .A2(new_n511), .A3(new_n515), .A4(new_n483), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n299), .A2(new_n301), .A3(G244), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n517), .A2(new_n518), .B1(G33), .B2(G283), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n400), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n266), .B2(G250), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n400), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n273), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n503), .A2(G257), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n492), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n283), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n256), .A2(G97), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n456), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G97), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n449), .B1(new_n310), .B2(new_n312), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n369), .A2(new_n204), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n358), .A2(new_n449), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n216), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n532), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n529), .B(new_n531), .C1(new_n540), .C2(new_n259), .ZN(new_n541));
  INV_X1    g0341(.A(new_n492), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n519), .B(new_n520), .C1(new_n400), .C2(new_n522), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n273), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(new_n421), .A3(new_n525), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n527), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n540), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n528), .B1(new_n547), .B2(new_n255), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n526), .A2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n544), .A2(G190), .A3(new_n525), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n531), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n516), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n510), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n499), .A2(G270), .A3(new_n272), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n492), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT81), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G303), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n311), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n400), .A2(G257), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G264), .A2(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n299), .A2(new_n301), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n273), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT82), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n559), .A2(new_n273), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n554), .A2(KEYINPUT81), .A3(new_n492), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n557), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n530), .A2(G116), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(G33), .B2(G283), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G33), .B2(new_n358), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n255), .C1(new_n216), .C2(G116), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  OAI221_X1 g0376(.A(new_n570), .B1(G116), .B2(new_n256), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n569), .A2(new_n577), .A3(G169), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n569), .A2(G200), .ZN(new_n581));
  INV_X1    g0381(.A(new_n577), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n557), .A2(G190), .A3(new_n567), .A4(new_n568), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n557), .A2(G179), .A3(new_n567), .A4(new_n568), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n569), .A2(new_n577), .A3(KEYINPUT21), .A4(G169), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n580), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n420), .A2(new_n553), .A3(new_n588), .ZN(G372));
  XOR2_X1   g0389(.A(new_n285), .B(KEYINPUT88), .Z(new_n590));
  OR2_X1    g0390(.A1(new_n368), .A2(new_n382), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n389), .A2(new_n390), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n336), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n318), .A2(new_n334), .B1(new_n342), .B2(new_n338), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(new_n346), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n414), .B1(new_n598), .B2(KEYINPUT89), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n594), .A2(new_n597), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT89), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n418), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n354), .A2(new_n391), .A3(new_n413), .A4(new_n417), .ZN(new_n604));
  INV_X1    g0404(.A(new_n509), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n580), .A2(new_n586), .A3(new_n587), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n516), .A2(new_n546), .A3(new_n551), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n436), .A2(new_n433), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(KEYINPUT85), .A3(G200), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT85), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n609), .B2(new_n367), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n461), .A2(new_n611), .A3(new_n463), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n283), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n439), .A2(new_n458), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n608), .A2(KEYINPUT86), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT86), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n552), .B2(new_n617), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n607), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n527), .A2(new_n545), .A3(new_n541), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n465), .A2(KEYINPUT26), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n617), .B2(new_n546), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(KEYINPUT87), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n616), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n624), .A2(KEYINPUT87), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n603), .B1(new_n604), .B2(new_n630), .ZN(G369));
  NAND2_X1  g0431(.A1(new_n509), .A2(new_n516), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n223), .A2(G20), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n215), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n484), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n605), .A2(new_n640), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n577), .A2(new_n640), .ZN(new_n645));
  MUX2_X1   g0445(.A(new_n606), .B(new_n588), .S(new_n645), .Z(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n646), .A3(G330), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n482), .A2(new_n483), .B1(new_n507), .B2(new_n421), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n640), .B(KEYINPUT90), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n506), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n640), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n606), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n633), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n647), .A2(new_n651), .A3(new_n655), .ZN(G399));
  NOR2_X1   g0456(.A1(new_n224), .A2(G41), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n450), .A2(G116), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n657), .A2(new_n659), .A3(new_n215), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT91), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  INV_X1    g0463(.A(new_n657), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n662), .B(new_n663), .C1(new_n220), .C2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n630), .A2(KEYINPUT29), .A3(new_n649), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n623), .A2(new_n625), .A3(new_n460), .A4(new_n464), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n617), .B2(new_n546), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n616), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT95), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n608), .B(new_n618), .C1(new_n605), .C2(new_n606), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT95), .A4(new_n616), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n675), .A2(KEYINPUT96), .A3(new_n652), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT96), .B1(new_n675), .B2(new_n652), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n667), .B1(new_n678), .B2(KEYINPUT29), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n544), .A2(new_n514), .A3(new_n497), .A4(new_n525), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n435), .A2(new_n438), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n681), .A2(new_n585), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n680), .B1(new_n683), .B2(KEYINPUT30), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n585), .A2(new_n682), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT92), .B(new_n685), .C1(new_n686), .C2(new_n681), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(KEYINPUT30), .ZN(new_n688));
  AOI21_X1  g0488(.A(G179), .B1(new_n544), .B2(new_n525), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n505), .A3(new_n610), .A4(new_n569), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n684), .A2(new_n687), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n640), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n460), .A2(new_n464), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n648), .B2(new_n506), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n588), .A2(new_n696), .A3(new_n608), .A4(new_n650), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT93), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n553), .A2(KEYINPUT93), .A3(new_n588), .A4(new_n650), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n688), .A2(new_n690), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n683), .A2(KEYINPUT30), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT31), .B(new_n649), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n704), .A2(KEYINPUT94), .A3(G330), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT94), .B1(new_n704), .B2(G330), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n679), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n666), .B1(new_n708), .B2(G1), .ZN(G364));
  NOR2_X1   g0509(.A1(new_n287), .A2(new_n367), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n216), .A2(G179), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G87), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n266), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT98), .Z(new_n716));
  NOR2_X1   g0516(.A1(new_n367), .A2(G190), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT99), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n716), .B1(new_n449), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT100), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n287), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n216), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n358), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n216), .A2(new_n421), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(new_n287), .A3(G200), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n717), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n727), .A2(G58), .B1(G68), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n725), .A2(new_n710), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n370), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n724), .B(new_n732), .C1(G77), .C2(new_n733), .ZN(new_n734));
  XOR2_X1   g0534(.A(KEYINPUT97), .B(G159), .Z(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n711), .A2(new_n287), .A3(new_n367), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT32), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n721), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n733), .ZN(new_n741));
  INV_X1    g0541(.A(G311), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G326), .ZN(new_n744));
  INV_X1    g0544(.A(G329), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n744), .A2(new_n731), .B1(new_n737), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(KEYINPUT33), .B(G317), .Z(new_n747));
  OAI22_X1  g0547(.A1(new_n723), .A2(new_n495), .B1(new_n747), .B2(new_n728), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n746), .B(new_n748), .C1(G322), .C2(new_n727), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n311), .B1(new_n712), .B2(new_n558), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT101), .Z(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n749), .B(new_n751), .C1(new_n752), .C2(new_n719), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n740), .B1(new_n743), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n221), .B1(G20), .B2(new_n283), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n755), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n304), .A2(new_n305), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n224), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n220), .A2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(G45), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n761), .B(new_n762), .C1(new_n244), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G355), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n225), .A2(new_n266), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n764), .B1(G116), .B2(new_n225), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n754), .A2(new_n755), .B1(new_n759), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n758), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n646), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n215), .B1(new_n634), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n657), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n646), .A2(G330), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n646), .A2(G330), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n774), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n770), .A2(new_n774), .B1(new_n775), .B2(new_n777), .ZN(G396));
  AND2_X1   g0578(.A1(new_n627), .A2(new_n616), .ZN(new_n779));
  INV_X1    g0579(.A(new_n629), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n619), .A2(new_n621), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n607), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n265), .A2(new_n640), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n289), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n590), .B2(new_n783), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n782), .A2(new_n650), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n782), .B2(new_n650), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(new_n707), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n774), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n727), .A2(G143), .B1(G150), .B2(new_n729), .ZN(new_n793));
  INV_X1    g0593(.A(G137), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n794), .B2(new_n731), .C1(new_n741), .C2(new_n736), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n713), .A2(G50), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n760), .B1(new_n798), .B2(new_n737), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT102), .ZN(new_n800));
  INV_X1    g0600(.A(new_n719), .ZN(new_n801));
  INV_X1    g0601(.A(new_n723), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n801), .A2(G68), .B1(G58), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G116), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n741), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n727), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n807), .A2(new_n495), .B1(new_n742), .B2(new_n737), .ZN(new_n808));
  INV_X1    g0608(.A(new_n731), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n266), .B(new_n808), .C1(G303), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n801), .A2(G87), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n712), .A2(new_n449), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n812), .B(new_n724), .C1(G283), .C2(new_n729), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n804), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n755), .A2(new_n756), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n815), .A2(new_n755), .B1(new_n204), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n773), .B(new_n817), .C1(new_n786), .C2(new_n757), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n792), .A2(new_n818), .ZN(G384));
  NAND2_X1  g0619(.A1(new_n596), .A2(new_n638), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n391), .B1(new_n380), .B2(new_n652), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n390), .B(new_n640), .C1(new_n389), .C2(new_n383), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n300), .A2(G33), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT73), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n827));
  AOI21_X1  g0627(.A(G20), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n312), .B1(new_n828), .B2(KEYINPUT7), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n295), .B1(new_n829), .B2(G68), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n259), .B1(new_n830), .B2(KEYINPUT16), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT16), .B2(new_n830), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n638), .B1(new_n832), .B2(new_n334), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n350), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n339), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n832), .A2(new_n334), .B1(new_n835), .B2(new_n638), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n318), .A2(new_n332), .A3(new_n334), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT37), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n638), .B1(new_n318), .B2(new_n334), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n348), .A2(new_n840), .A3(new_n841), .A4(new_n335), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n834), .A2(KEYINPUT38), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT38), .B1(new_n834), .B2(new_n843), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n285), .A2(new_n640), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n823), .B1(new_n845), .B2(new_n846), .C1(new_n788), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT39), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT103), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n837), .A2(new_n839), .ZN(new_n853));
  INV_X1    g0653(.A(new_n595), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n841), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n334), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT7), .B1(new_n311), .B2(new_n216), .ZN(new_n857));
  OAI21_X1  g0657(.A(G68), .B1(new_n857), .B2(new_n302), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n296), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT74), .B1(new_n859), .B2(new_n309), .ZN(new_n860));
  INV_X1    g0660(.A(new_n317), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n856), .B1(new_n862), .B2(new_n831), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n841), .B(new_n335), .C1(new_n863), .C2(new_n638), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n345), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n852), .B1(new_n855), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT17), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n335), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n839), .B1(new_n596), .B2(new_n868), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n837), .A2(new_n595), .A3(new_n839), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n842), .B(KEYINPUT103), .C1(new_n870), .C2(new_n841), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n866), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n872), .A2(KEYINPUT104), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT104), .B1(new_n872), .B2(new_n873), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n874), .A2(new_n875), .A3(new_n845), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n851), .B1(new_n876), .B2(KEYINPUT39), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n593), .A2(new_n652), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n820), .B(new_n848), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n599), .A2(new_n602), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n417), .ZN(new_n881));
  INV_X1    g0681(.A(new_n667), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n675), .A2(new_n652), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT96), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n675), .A2(KEYINPUT96), .A3(new_n652), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(KEYINPUT29), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n604), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n879), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n872), .A2(new_n873), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT104), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n872), .A2(KEYINPUT104), .A3(new_n873), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n844), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n785), .B1(new_n821), .B2(new_n822), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(KEYINPUT40), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n898), .B(new_n896), .C1(new_n845), .C2(new_n846), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n895), .A2(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n420), .A2(new_n898), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(G330), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n890), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n215), .B2(new_n634), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n537), .A2(new_n538), .ZN(new_n909));
  OAI211_X1 g0709(.A(G20), .B(new_n270), .C1(new_n909), .C2(KEYINPUT35), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n805), .B(new_n910), .C1(KEYINPUT35), .C2(new_n909), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT36), .Z(new_n912));
  OAI21_X1  g0712(.A(G77), .B1(new_n290), .B2(new_n209), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n913), .A2(new_n220), .B1(G50), .B2(new_n209), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n223), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n912), .A3(new_n915), .ZN(G367));
  INV_X1    g0716(.A(G150), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n266), .B1(new_n807), .B2(new_n917), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n741), .A2(new_n370), .B1(new_n728), .B2(new_n736), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n918), .B(new_n919), .C1(G143), .C2(new_n809), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n712), .A2(new_n290), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n723), .A2(new_n209), .ZN(new_n922));
  INV_X1    g0722(.A(new_n718), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n921), .B(new_n922), .C1(G77), .C2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n920), .B(new_n924), .C1(new_n794), .C2(new_n737), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n731), .A2(new_n742), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n741), .A2(new_n752), .B1(new_n449), .B2(new_n723), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(G97), .B2(new_n923), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n713), .A2(G116), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT46), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n760), .B1(G294), .B2(new_n729), .ZN(new_n931));
  INV_X1    g0731(.A(new_n737), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n727), .A2(G303), .B1(G317), .B2(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n928), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n925), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT47), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n774), .B1(new_n936), .B2(new_n755), .ZN(new_n937));
  INV_X1    g0737(.A(new_n761), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n759), .B1(new_n225), .B2(new_n457), .C1(new_n236), .C2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n463), .A2(new_n652), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n940), .A2(new_n439), .A3(new_n458), .A4(new_n615), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n617), .B2(new_n940), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(new_n769), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n937), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n647), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n644), .B1(G330), .B2(new_n646), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n654), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n644), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n776), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n647), .A3(new_n653), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n649), .A2(new_n541), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n551), .A2(new_n546), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n623), .A2(new_n649), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n651), .B(new_n956), .C1(new_n653), .C2(new_n632), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT45), .Z(new_n958));
  OAI21_X1  g0758(.A(new_n651), .B1(new_n653), .B2(new_n632), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT44), .B1(new_n960), .B2(new_n956), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  INV_X1    g0762(.A(new_n956), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n647), .A3(new_n961), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n964), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n957), .B(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n945), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n679), .B(new_n707), .C1(new_n952), .C2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n657), .B(KEYINPUT41), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n970), .A2(KEYINPUT106), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT106), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n972), .A2(new_n973), .A3(new_n772), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT107), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n655), .A2(new_n963), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT42), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n546), .B1(new_n954), .B2(new_n509), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n650), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n942), .B(KEYINPUT43), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT105), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n977), .A2(new_n984), .A3(new_n979), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT105), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n986), .A3(new_n981), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n945), .A2(new_n956), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n974), .A2(new_n975), .A3(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n988), .B(new_n989), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n970), .A2(new_n971), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT106), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n970), .A2(KEYINPUT106), .A3(new_n971), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n771), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT107), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n944), .B1(new_n991), .B2(new_n998), .ZN(G387));
  INV_X1    g0799(.A(new_n760), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n805), .B2(new_n718), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n727), .A2(G317), .B1(G311), .B2(new_n729), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n558), .B2(new_n741), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G322), .B2(new_n809), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT48), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n752), .B2(new_n723), .C1(new_n495), .C2(new_n712), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT49), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .C1(new_n744), .C2(new_n737), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n712), .A2(new_n204), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n457), .A2(new_n723), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G68), .C2(new_n733), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1000), .B1(new_n247), .B2(new_n729), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G159), .A2(new_n809), .B1(new_n932), .B2(G150), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n370), .B2(new_n807), .C1(new_n358), .C2(new_n719), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n761), .B1(new_n232), .B2(new_n763), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n658), .B2(new_n766), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n209), .A2(new_n204), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n247), .A2(new_n1021), .A3(new_n370), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT50), .B1(new_n246), .B2(G50), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1022), .A2(new_n763), .A3(new_n658), .A4(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1019), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(G107), .B2(new_n225), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1017), .A2(new_n755), .B1(new_n759), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n773), .C1(new_n644), .C2(new_n769), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n708), .A2(new_n951), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n657), .B1(new_n708), .B2(new_n951), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1028), .B1(new_n771), .B2(new_n952), .C1(new_n1029), .C2(new_n1030), .ZN(G393));
  INV_X1    g0831(.A(new_n969), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n708), .A2(new_n951), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT108), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT108), .B2(new_n968), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n657), .B(new_n1033), .C1(new_n1029), .C2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n963), .A2(new_n758), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n759), .B1(new_n358), .B2(new_n225), .C1(new_n241), .C2(new_n938), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n727), .A2(G159), .B1(new_n809), .B2(G150), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT109), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n733), .A2(new_n247), .B1(G50), .B2(new_n729), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n802), .A2(G77), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n713), .A2(G68), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1000), .B1(G143), .B2(new_n932), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n811), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n712), .A2(new_n752), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n311), .B1(new_n741), .B2(new_n495), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n727), .A2(G311), .B1(new_n809), .B2(G317), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(KEYINPUT52), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n932), .A2(G322), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n723), .A2(new_n805), .B1(new_n728), .B2(new_n558), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n801), .B2(G107), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1041), .A2(new_n1047), .B1(new_n1048), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n774), .B1(new_n1057), .B2(new_n755), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n1037), .A2(new_n1038), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1035), .B2(new_n772), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1036), .A2(new_n1060), .ZN(G390));
  NAND3_X1  g0861(.A1(new_n898), .A2(G330), .A3(new_n786), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n823), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n895), .A2(new_n878), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n786), .B1(new_n676), .B2(new_n677), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n847), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT110), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n785), .B1(new_n885), .B2(new_n886), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n823), .B1(new_n1071), .B2(new_n847), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT110), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1072), .A2(new_n1073), .A3(new_n878), .A4(new_n895), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n788), .A2(new_n847), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n878), .B1(new_n1076), .B2(new_n1063), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n877), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1065), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n786), .B(new_n823), .C1(new_n705), .C2(new_n706), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1071), .A2(new_n847), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n786), .B1(new_n705), .B2(new_n706), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1064), .B1(new_n1085), .B2(new_n1063), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1084), .B1(new_n1086), .B2(new_n1076), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n420), .A2(G330), .A3(new_n898), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n881), .A2(new_n1088), .A3(new_n888), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT111), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1075), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1080), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT111), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1075), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n1079), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(new_n1097), .A3(new_n657), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n733), .A2(G97), .B1(G107), .B2(new_n729), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n752), .B2(new_n731), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT113), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n266), .B1(new_n727), .B2(G116), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n714), .A3(new_n1043), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G68), .B2(new_n801), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(new_n495), .C2(new_n737), .ZN(new_n1105));
  INV_X1    g0905(.A(G128), .ZN(new_n1106));
  INV_X1    g0906(.A(G125), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1106), .A2(new_n731), .B1(new_n737), .B2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G159), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n741), .A2(new_n1110), .B1(new_n1111), .B2(new_n723), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1108), .B(new_n1112), .C1(G132), .C2(new_n727), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n712), .A2(new_n917), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1113), .B(new_n1115), .C1(new_n794), .C2(new_n728), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n266), .B1(new_n718), .B2(new_n370), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT112), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1105), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1119), .A2(new_n755), .B1(new_n246), .B2(new_n816), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n850), .B1(new_n895), .B2(new_n849), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n773), .B(new_n1120), .C1(new_n1121), .C2(new_n757), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1096), .A2(new_n1079), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n772), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1098), .A2(new_n1125), .ZN(G378));
  NAND2_X1  g0926(.A1(new_n413), .A2(new_n417), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n397), .A2(new_n638), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1130), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n413), .A2(new_n417), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1132), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n756), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n816), .A2(new_n370), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1010), .B1(G58), .B2(new_n923), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n752), .B2(new_n737), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1141), .A2(G41), .A3(new_n760), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT114), .Z(new_n1143));
  OAI22_X1  g0943(.A1(new_n741), .A2(new_n457), .B1(new_n358), .B2(new_n728), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n922), .B(new_n1144), .C1(G107), .C2(new_n727), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(new_n805), .C2(new_n731), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT58), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n733), .A2(G137), .B1(G132), .B2(new_n729), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT115), .Z(new_n1149));
  OAI22_X1  g0949(.A1(new_n807), .A2(new_n1106), .B1(new_n917), .B2(new_n723), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n713), .B2(new_n1109), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(new_n1107), .C2(new_n731), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT59), .Z(new_n1153));
  AOI21_X1  g0953(.A(G41), .B1(new_n923), .B2(new_n735), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G33), .B1(new_n932), .B2(G124), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G41), .B1(new_n760), .B2(G33), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1147), .B(new_n1156), .C1(G50), .C2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n774), .B1(new_n1158), .B2(new_n755), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1138), .A2(new_n1139), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n902), .A2(new_n901), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(G330), .C1(new_n876), .C2(new_n899), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT118), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n903), .B2(G330), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n879), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n846), .ZN(new_n1170));
  AOI221_X4 g0970(.A(new_n1063), .B1(new_n1170), .B2(new_n844), .C1(new_n787), .C2(new_n1068), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n878), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1121), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n895), .A2(new_n900), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1164), .A2(new_n1174), .A3(G330), .A4(new_n1161), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1169), .A2(new_n1173), .A3(new_n820), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1168), .A2(new_n1176), .A3(KEYINPUT119), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT119), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n879), .B(new_n1178), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1160), .B1(new_n1180), .B2(new_n771), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1070), .A2(new_n1074), .B1(new_n1077), .B2(new_n877), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1093), .B(new_n1087), .C1(new_n1183), .C2(new_n1065), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1089), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1168), .B2(new_n1176), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n657), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT57), .B1(new_n1190), .B2(new_n1185), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1182), .B1(new_n1189), .B2(new_n1191), .ZN(G375));
  NAND3_X1  g0992(.A1(new_n420), .A2(G330), .A3(new_n898), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n603), .B(new_n1193), .C1(new_n604), .C2(new_n679), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1194), .B(new_n1084), .C1(new_n1076), .C2(new_n1086), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n971), .B(KEYINPUT120), .Z(new_n1196));
  NAND3_X1  g0996(.A1(new_n1090), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n774), .B1(new_n209), .B2(new_n816), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT121), .Z(new_n1199));
  NOR2_X1   g0999(.A1(new_n823), .A2(new_n757), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n807), .A2(new_n794), .B1(new_n1106), .B2(new_n737), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1000), .B(new_n1201), .C1(G58), .C2(new_n923), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n723), .A2(new_n370), .B1(new_n712), .B2(new_n1111), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1110), .A2(new_n728), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G150), .C2(new_n733), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(new_n798), .C2(new_n731), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n737), .A2(new_n558), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1011), .B1(G283), .B2(new_n727), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT123), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n733), .A2(G107), .B1(G116), .B2(new_n729), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT122), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n311), .B1(new_n712), .B2(new_n358), .C1(new_n495), .C2(new_n731), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n801), .B2(G77), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1209), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1206), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1199), .B(new_n1200), .C1(new_n755), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1087), .B2(new_n772), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1197), .A2(new_n1217), .ZN(G381));
  INV_X1    g1018(.A(G378), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n1182), .C1(new_n1191), .C2(new_n1189), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1220), .A2(G384), .A3(G381), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n975), .B1(new_n974), .B2(new_n990), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n992), .A2(new_n997), .A3(KEYINPUT107), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G390), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n944), .A3(new_n1225), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1226), .A2(G396), .A3(G393), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(G407));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(G343), .C2(new_n1220), .ZN(G409));
  XNOR2_X1  g1029(.A(G393), .B(G396), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1225), .B1(new_n1224), .B2(new_n944), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n944), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1233), .B(G390), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1231), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(G390), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n1226), .A3(new_n1230), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G375), .A2(G378), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n639), .A2(G213), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1098), .A2(new_n1125), .A3(new_n1160), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1190), .A2(new_n1185), .A3(new_n1196), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT124), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1190), .A2(new_n1185), .A3(new_n1244), .A4(new_n1196), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1168), .A2(new_n1176), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n772), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1241), .A2(new_n1243), .A3(new_n1245), .A4(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1239), .A2(new_n1240), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n639), .A2(G213), .A3(G2897), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1195), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1195), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n664), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1195), .A2(new_n1255), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1253), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1259), .A2(G384), .A3(new_n1217), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1259), .B2(new_n1217), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1251), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1217), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1259), .A2(G384), .A3(new_n1217), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1250), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1262), .A2(new_n1267), .ZN(new_n1268));
  AOI211_X1 g1068(.A(KEYINPUT61), .B(new_n1238), .C1(new_n1249), .C2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1239), .A2(new_n1240), .A3(new_n1248), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT126), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1271), .A2(new_n1275), .A3(new_n1272), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1269), .A2(new_n1274), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1249), .B2(new_n1268), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1271), .A2(KEYINPUT62), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G375), .A2(G378), .B1(G213), .B2(new_n639), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1248), .A4(new_n1270), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(new_n1280), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1238), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(new_n1239), .A2(new_n1220), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1238), .A2(new_n1220), .A3(new_n1239), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1270), .ZN(G402));
endmodule


