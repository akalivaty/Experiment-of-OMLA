//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G228gat), .A2(G233gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n208), .B1(G155gat), .B2(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT78), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  OR2_X1    g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT78), .A3(new_n211), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221));
  NAND2_X1  g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT22), .ZN(new_n224));
  INV_X1    g023(.A(G197gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT71), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT71), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G197gat), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n226), .A2(new_n228), .A3(G204gat), .ZN(new_n229));
  AOI21_X1  g028(.A(G204gat), .B1(new_n226), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G211gat), .A2(G218gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT72), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n222), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT72), .B1(new_n223), .B2(new_n232), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G204gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n227), .A2(G197gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT71), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n228), .A3(G204gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n244), .A2(new_n224), .B1(new_n236), .B2(new_n235), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n221), .B1(new_n238), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n220), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT29), .B1(new_n220), .B2(new_n247), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n244), .A2(new_n236), .A3(new_n235), .A4(new_n224), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n237), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n206), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G22gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n213), .A2(KEYINPUT79), .A3(new_n219), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n218), .A2(KEYINPUT78), .A3(new_n211), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n211), .B1(new_n218), .B2(KEYINPUT78), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT29), .B1(new_n250), .B2(new_n251), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n256), .B(new_n260), .C1(new_n261), .C2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT73), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n238), .B2(new_n245), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n258), .A2(new_n259), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n221), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT73), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n206), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n262), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n254), .A2(new_n255), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n255), .B1(new_n254), .B2(new_n270), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n205), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n262), .A2(new_n269), .A3(new_n268), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n265), .B1(new_n261), .B2(KEYINPUT3), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n250), .A3(new_n251), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(G22gat), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n205), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n254), .A2(new_n255), .A3(new_n270), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n273), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n274), .B1(new_n273), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT66), .B1(new_n286), .B2(G120gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(G120gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(G120gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n287), .A2(new_n290), .A3(KEYINPUT67), .A4(new_n291), .ZN(new_n295));
  INV_X1    g094(.A(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G127gat), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G134gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT1), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n294), .A2(new_n295), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n289), .A2(G113gat), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n303), .A2(new_n291), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n304), .B2(KEYINPUT1), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n260), .A3(new_n256), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n220), .A2(new_n305), .A3(new_n302), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT4), .B1(new_n306), .B2(new_n265), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n220), .A2(new_n315), .A3(new_n305), .A4(new_n302), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(KEYINPUT80), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n260), .A2(new_n256), .A3(KEYINPUT3), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n220), .A2(new_n247), .B1(new_n302), .B2(new_n305), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n311), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n308), .A2(new_n321), .A3(KEYINPUT4), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n310), .B1(new_n307), .B2(new_n308), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n313), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n314), .A2(new_n316), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n320), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G1gat), .B(G29gat), .Z(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(KEYINPUT6), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n336), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n328), .B2(new_n330), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n327), .A2(new_n323), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n325), .A2(new_n324), .A3(new_n326), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n339), .B(new_n330), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(KEYINPUT83), .A3(new_n344), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT74), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n221), .ZN(new_n352));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT27), .B(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT28), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G183gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT27), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G183gat), .ZN(new_n370));
  AND4_X1   g169(.A1(KEYINPUT28), .A2(new_n368), .A3(new_n370), .A4(new_n365), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n362), .B(new_n363), .C1(new_n366), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n359), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n357), .ZN(new_n377));
  AND3_X1   g176(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n379));
  OAI21_X1  g178(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n374), .A2(new_n375), .B1(new_n355), .B2(new_n356), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n379), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n365), .B2(new_n379), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT25), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n372), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT75), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n382), .B1(new_n377), .B2(new_n381), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT25), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n372), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n352), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n388), .A2(new_n351), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n252), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n351), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n264), .A2(new_n267), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n388), .A2(new_n221), .A3(new_n351), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT76), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT76), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n403), .A2(new_n410), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n402), .A3(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT77), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n397), .A2(new_n416), .A3(new_n402), .A4(new_n406), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT30), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n412), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n285), .B1(new_n349), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT68), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n388), .B2(new_n306), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n302), .A2(new_n305), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(KEYINPUT68), .A3(new_n392), .A4(new_n372), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n388), .A2(new_n306), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n429), .B(KEYINPUT64), .Z(new_n430));
  OR3_X1    g229(.A1(new_n428), .A2(KEYINPUT34), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n429), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT34), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT32), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n428), .B2(new_n430), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT33), .B1(new_n428), .B2(new_n430), .ZN(new_n437));
  XOR2_X1   g236(.A(G15gat), .B(G43gat), .Z(new_n438));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n436), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  AOI221_X4 g241(.A(new_n435), .B1(KEYINPUT33), .B2(new_n440), .C1(new_n428), .C2(new_n430), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n434), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n430), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT32), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n448), .A3(new_n440), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n436), .B1(new_n437), .B2(new_n441), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n433), .A4(new_n431), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n451), .A3(KEYINPUT70), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT36), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT70), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n454), .B(new_n434), .C1(new_n442), .C2(new_n443), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n444), .A2(new_n451), .A3(KEYINPUT69), .A4(KEYINPUT36), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n444), .A2(new_n451), .A3(KEYINPUT36), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n422), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n331), .A2(new_n336), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n344), .A3(new_n343), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n395), .A2(new_n252), .A3(new_n396), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT37), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n407), .A2(KEYINPUT37), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n408), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n414), .A2(new_n417), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n337), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n340), .A2(KEYINPUT86), .A3(KEYINPUT6), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n463), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  AND4_X1   g281(.A1(KEYINPUT86), .A2(new_n331), .A3(KEYINPUT6), .A4(new_n336), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT86), .B1(new_n340), .B2(KEYINPUT6), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n475), .B1(new_n473), .B2(new_n470), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n465), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n403), .A2(KEYINPUT37), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT38), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n318), .A2(new_n319), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n310), .B1(new_n329), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT39), .B1(new_n309), .B2(new_n311), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT39), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n497), .A2(KEYINPUT85), .A3(new_n339), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT85), .B1(new_n497), .B2(new_n339), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT40), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT40), .B(new_n495), .C1(new_n498), .C2(new_n499), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n409), .A2(new_n411), .B1(KEYINPUT30), .B2(new_n419), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n340), .B1(new_n506), .B2(new_n418), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n285), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n462), .B1(new_n491), .B2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n510));
  AND4_X1   g309(.A1(new_n418), .A2(new_n412), .A3(new_n420), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n452), .A2(new_n455), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n273), .A2(new_n282), .ZN(new_n513));
  INV_X1    g312(.A(new_n274), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n273), .A2(new_n274), .A3(new_n282), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n479), .A2(new_n465), .A3(new_n480), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n511), .A2(new_n512), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n444), .A2(new_n451), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT89), .B1(new_n285), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n345), .A2(new_n346), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n464), .A3(new_n348), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n421), .B1(new_n524), .B2(new_n337), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  INV_X1    g325(.A(new_n521), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n517), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n520), .B1(new_n529), .B2(KEYINPUT35), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n202), .B1(new_n509), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n519), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n491), .A2(new_n508), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n422), .A2(new_n461), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n536), .A3(KEYINPUT90), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(G1gat), .ZN(new_n539));
  AOI21_X1  g338(.A(G8gat), .B1(new_n539), .B2(KEYINPUT94), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n538), .B1(new_n541), .B2(G1gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n540), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT92), .Z(new_n546));
  INV_X1    g345(.A(G43gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n204), .ZN(new_n548));
  NOR2_X1   g347(.A1(G43gat), .A2(G50gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT15), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n546), .B(new_n550), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT93), .B(G50gat), .Z(new_n555));
  AOI211_X1 g354(.A(KEYINPUT15), .B(new_n548), .C1(new_n555), .C2(new_n547), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n553), .B1(KEYINPUT91), .B2(new_n551), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(KEYINPUT91), .B2(new_n551), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n550), .B1(new_n559), .B2(new_n546), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n544), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n554), .A2(new_n556), .ZN(new_n563));
  INV_X1    g362(.A(new_n560), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT17), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n557), .B2(new_n560), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n544), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n544), .B(new_n561), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n569), .B(KEYINPUT13), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n562), .A2(new_n568), .A3(KEYINPUT18), .A4(new_n569), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G197gat), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT11), .B(G169gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT12), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n572), .A2(new_n575), .A3(new_n582), .A4(new_n576), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n584), .A2(KEYINPUT95), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT95), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n531), .A2(new_n537), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n349), .ZN(new_n591));
  XOR2_X1   g390(.A(G57gat), .B(G64gat), .Z(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT9), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(KEYINPUT96), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G71gat), .B(G78gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n544), .B1(new_n611), .B2(new_n599), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n608), .A2(new_n614), .A3(new_n609), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  INV_X1    g422(.A(G85gat), .ZN(new_n624));
  INV_X1    g423(.A(G92gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(KEYINPUT8), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G99gat), .B(G106gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT101), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n561), .ZN(new_n633));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT99), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n633), .B1(KEYINPUT41), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n565), .A2(new_n567), .A3(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n636), .A2(KEYINPUT41), .ZN(new_n643));
  XOR2_X1   g442(.A(G134gat), .B(G162gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n641), .B2(new_n642), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n632), .A2(new_n599), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n630), .A2(new_n598), .A3(new_n631), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n653), .A2(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n651), .A2(new_n653), .ZN(new_n661));
  INV_X1    g460(.A(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  AOI21_X1  g465(.A(new_n662), .B1(new_n654), .B2(new_n655), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n660), .A2(new_n663), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n666), .ZN(new_n670));
  INV_X1    g469(.A(new_n663), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(new_n667), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n618), .A2(new_n650), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n591), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(G1gat), .Z(G1324gat));
  NAND2_X1  g477(.A1(new_n590), .A2(new_n421), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n676), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(G8gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(new_n680), .ZN(new_n684));
  MUX2_X1   g483(.A(new_n682), .B(new_n684), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g484(.A1(new_n590), .A2(new_n512), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(G15gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n675), .ZN(new_n689));
  INV_X1    g488(.A(new_n461), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n590), .A2(new_n675), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n688), .B2(new_n691), .ZN(G1326gat));
  NAND3_X1  g491(.A1(new_n590), .A2(new_n675), .A3(new_n285), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(new_n618), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n673), .B(KEYINPUT104), .Z(new_n697));
  AND3_X1   g496(.A1(new_n584), .A2(KEYINPUT103), .A3(new_n585), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT103), .B1(new_n584), .B2(new_n585), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n696), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n531), .A2(new_n537), .A3(new_n650), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n707), .A3(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n421), .A2(new_n464), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n517), .B1(new_n710), .B2(new_n504), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n486), .A2(new_n479), .A3(new_n480), .A4(new_n465), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n712), .A2(new_n463), .B1(KEYINPUT38), .B2(new_n489), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n713), .B2(new_n487), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(KEYINPUT106), .A3(new_n462), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n534), .B2(new_n535), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n533), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(new_n719), .A3(new_n650), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT106), .B1(new_n714), .B2(new_n462), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n534), .A2(new_n535), .A3(new_n716), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n649), .B1(new_n725), .B2(new_n533), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(KEYINPUT107), .A3(new_n719), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n703), .B1(new_n709), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n349), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G29gat), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n696), .A2(new_n649), .A3(new_n674), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(G29gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n591), .B2(new_n735), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n591), .A2(new_n732), .A3(new_n735), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n731), .A2(new_n736), .A3(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(G36gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT46), .B1(new_n679), .B2(new_n740), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n679), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n729), .A2(new_n421), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n739), .ZN(G1329gat));
  NOR2_X1   g543(.A1(new_n734), .A2(G43gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n687), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT47), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n547), .B1(new_n729), .B2(new_n690), .ZN(new_n749));
  INV_X1    g548(.A(new_n746), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n720), .A2(new_n721), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT107), .B1(new_n726), .B2(new_n719), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n704), .A2(new_n707), .A3(KEYINPUT44), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n707), .B1(new_n704), .B2(KEYINPUT44), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n690), .A3(new_n702), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  INV_X1    g557(.A(new_n748), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n746), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n751), .A2(new_n760), .ZN(G1330gat));
  NOR2_X1   g560(.A1(new_n517), .A2(new_n555), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n756), .A2(new_n702), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n590), .A2(new_n285), .A3(new_n733), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n555), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n763), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n765), .B1(new_n763), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(G1331gat));
  NAND4_X1  g570(.A1(new_n697), .A2(new_n696), .A3(new_n649), .A4(new_n701), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n725), .B2(new_n533), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n349), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G57gat), .ZN(G1332gat));
  INV_X1    g574(.A(new_n421), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT110), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1333gat));
  NAND3_X1  g580(.A1(new_n773), .A2(G71gat), .A3(new_n690), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT111), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n512), .B(KEYINPUT112), .Z(new_n784));
  AND2_X1   g583(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(G71gat), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n285), .ZN(new_n789));
  XNOR2_X1  g588(.A(KEYINPUT114), .B(G78gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n696), .A2(new_n700), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n726), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT51), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n673), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n624), .A3(new_n349), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n674), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n709), .B2(new_n728), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n349), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n799), .B2(new_n624), .ZN(G1336gat));
  AOI21_X1  g599(.A(new_n625), .B1(new_n798), .B2(new_n421), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n697), .A2(new_n625), .A3(new_n421), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n797), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n756), .A2(new_n421), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G92gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n794), .A2(new_n802), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n810), .ZN(G1337gat));
  INV_X1    g610(.A(G99gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n812), .A3(new_n512), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n798), .A2(new_n690), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n812), .ZN(G1338gat));
  INV_X1    g614(.A(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n798), .B2(new_n285), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n697), .A2(new_n816), .A3(new_n285), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT115), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n794), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT53), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n756), .A2(new_n285), .A3(new_n805), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n794), .A2(new_n820), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n822), .A2(new_n827), .ZN(G1339gat));
  INV_X1    g627(.A(new_n349), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n659), .B(new_n662), .C1(new_n654), .C2(new_n655), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n654), .A2(new_n655), .A3(new_n662), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n666), .B1(new_n667), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n830), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n660), .A2(new_n668), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT55), .B(new_n837), .C1(new_n840), .C2(new_n834), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n841), .A3(new_n669), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n839), .A2(new_n841), .A3(new_n844), .A4(new_n669), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n700), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n573), .A2(new_n574), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n569), .B1(new_n562), .B2(new_n568), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n581), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n585), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n674), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n650), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n649), .A2(new_n850), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n843), .A2(new_n854), .A3(new_n845), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n618), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n675), .A2(new_n701), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n829), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n522), .A2(new_n776), .A3(new_n528), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n700), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n285), .B1(new_n857), .B2(new_n858), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(new_n349), .A3(new_n776), .A4(new_n512), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n865), .A2(new_n286), .A3(new_n588), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n863), .A2(new_n866), .ZN(G1340gat));
  AOI21_X1  g666(.A(G120gat), .B1(new_n862), .B2(new_n674), .ZN(new_n868));
  INV_X1    g667(.A(new_n697), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n865), .A2(new_n289), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n868), .A2(new_n870), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n865), .B2(new_n618), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n696), .A2(new_n298), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n861), .B2(new_n873), .ZN(G1342gat));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n296), .A3(new_n650), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n865), .B2(new_n649), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n349), .A2(new_n776), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n690), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n517), .B1(new_n857), .B2(new_n858), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n842), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n839), .A2(new_n841), .A3(KEYINPUT117), .A4(new_n669), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n589), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n650), .B1(new_n889), .B2(new_n852), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n855), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n588), .B1(new_n886), .B2(new_n842), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n893), .A2(new_n888), .B1(new_n674), .B2(new_n851), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(KEYINPUT118), .A3(new_n650), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n618), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n517), .B1(new_n896), .B2(new_n858), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n885), .B1(new_n897), .B2(new_n884), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT118), .B1(new_n894), .B2(new_n650), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n890), .A2(new_n891), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n855), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n902), .A2(new_n618), .B1(new_n675), .B2(new_n701), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n517), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n885), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n906), .A3(new_n700), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n690), .A2(new_n517), .A3(new_n421), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n859), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n588), .A2(G141gat), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n907), .A2(G141gat), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n859), .A2(new_n908), .A3(new_n910), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n904), .A2(new_n589), .A3(new_n885), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(G141gat), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT120), .B(new_n914), .C1(new_n915), .C2(G141gat), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n911), .A2(new_n912), .B1(new_n918), .B2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(G148gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n909), .A2(new_n921), .A3(new_n674), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G148gat), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n899), .A2(new_n906), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n674), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n883), .A2(new_n884), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n842), .A2(new_n649), .A3(new_n850), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n618), .B1(new_n890), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n675), .A2(new_n588), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT57), .B(new_n517), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n674), .B1(new_n881), .B2(KEYINPUT121), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(KEYINPUT121), .B2(new_n881), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT122), .B(KEYINPUT59), .C1(new_n935), .C2(new_n921), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n921), .B1(new_n932), .B2(new_n934), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n923), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n922), .B1(new_n926), .B2(new_n940), .ZN(G1345gat));
  NAND4_X1  g740(.A1(new_n899), .A2(new_n906), .A3(G155gat), .A4(new_n696), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n909), .A2(new_n696), .ZN(new_n943));
  INV_X1    g742(.A(G155gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(KEYINPUT123), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1346gat));
  AOI21_X1  g749(.A(G162gat), .B1(new_n909), .B2(new_n650), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n650), .A2(G162gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n925), .B2(new_n952), .ZN(G1347gat));
  AOI21_X1  g752(.A(new_n349), .B1(new_n857), .B2(new_n858), .ZN(new_n954));
  AND4_X1   g753(.A1(new_n421), .A2(new_n954), .A3(new_n522), .A4(new_n528), .ZN(new_n955));
  AOI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n700), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n349), .A2(new_n776), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n784), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n864), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n589), .A2(G169gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(G1348gat));
  INV_X1    g761(.A(G176gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n955), .A2(new_n963), .A3(new_n674), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n960), .A2(new_n697), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n963), .ZN(G1349gat));
  AOI21_X1  g765(.A(new_n367), .B1(new_n960), .B2(new_n696), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n955), .A2(new_n696), .A3(new_n364), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT125), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n967), .A2(KEYINPUT60), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT60), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1350gat));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n365), .A3(new_n650), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  OAI21_X1  g773(.A(G190gat), .B1(new_n974), .B2(KEYINPUT126), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n960), .B2(new_n650), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT126), .A3(new_n974), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(KEYINPUT126), .B2(new_n974), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(G1351gat));
  NAND2_X1  g778(.A1(new_n461), .A2(new_n957), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n932), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n982), .A2(new_n225), .A3(new_n588), .ZN(new_n983));
  AND4_X1   g782(.A1(new_n285), .A2(new_n954), .A3(new_n421), .A4(new_n461), .ZN(new_n984));
  AOI21_X1  g783(.A(G197gat), .B1(new_n984), .B2(new_n700), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n983), .A2(new_n985), .ZN(G1352gat));
  NAND3_X1  g785(.A1(new_n984), .A2(new_n239), .A3(new_n674), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT62), .Z(new_n988));
  OAI21_X1  g787(.A(G204gat), .B1(new_n982), .B2(new_n869), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1353gat));
  INV_X1    g789(.A(G211gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n984), .A2(new_n991), .A3(new_n696), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n932), .A2(new_n696), .A3(new_n981), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n993), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1354gat));
  OAI21_X1  g796(.A(G218gat), .B1(new_n982), .B2(new_n649), .ZN(new_n998));
  INV_X1    g797(.A(G218gat), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n999), .A3(new_n650), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(G1355gat));
endmodule


