//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n548, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n466));
  OAI22_X1  g041(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n464), .B2(new_n463), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(G160));
  OAI221_X1 g051(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n472), .C2(G112), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT69), .Z(new_n478));
  INV_X1    g053(.A(new_n463), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(new_n466), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n464), .A2(new_n463), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n478), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  AND3_X1   g065(.A1(new_n461), .A2(G102), .A3(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(G126), .B1(new_n464), .B2(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n491), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n479), .A2(new_n480), .B1(new_n470), .B2(new_n471), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G138), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n467), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n495), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n497), .B1(new_n467), .B2(new_n501), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n481), .A2(new_n472), .A3(G138), .A4(new_n498), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(new_n495), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n516), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G88), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n518), .B(new_n521), .C1(new_n522), .C2(new_n513), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  XOR2_X1   g099(.A(KEYINPUT73), .B(G51), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n519), .A2(G89), .A3(new_n520), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n528), .A2(KEYINPUT74), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT74), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n526), .B(new_n527), .C1(new_n531), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n517), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n519), .A2(new_n520), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n535), .B1(new_n536), .B2(new_n537), .C1(new_n513), .C2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND3_X1  g115(.A1(new_n519), .A2(G43), .A3(G543), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT75), .B(G81), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n519), .A2(new_n520), .A3(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(new_n513), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT76), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  AND3_X1   g128(.A1(new_n515), .A2(KEYINPUT6), .A3(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT6), .B1(new_n515), .B2(G651), .ZN(new_n555));
  OAI211_X1 g130(.A(G53), .B(G543), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n517), .A2(new_n558), .A3(G53), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n557), .A2(KEYINPUT77), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT77), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n565), .A3(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(G651), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n536), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n562), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(new_n517), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n519), .A2(G87), .A3(new_n520), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n563), .A2(new_n565), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT79), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n520), .A2(new_n586), .A3(G61), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n517), .A2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n573), .A2(G86), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n517), .A2(G47), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n519), .A2(G85), .A3(new_n520), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n513), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n536), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .A4(new_n520), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n517), .A2(G54), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n513), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n597), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n597), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n576), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n576), .B2(G868), .ZN(G280));
  XNOR2_X1  g186(.A(KEYINPUT80), .B(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(G860), .B2(new_n612), .ZN(G148));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n487), .A2(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT81), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n622), .A2(KEYINPUT82), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(KEYINPUT82), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n484), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n487), .A2(G135), .ZN(new_n627));
  OAI221_X1 g202(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n472), .C2(G111), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n625), .B(new_n631), .C1(new_n623), .C2(new_n621), .ZN(G156));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n638), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT17), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n648), .B2(new_n651), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n647), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n649), .A2(new_n651), .A3(new_n647), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n630), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n630), .B1(new_n658), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n622), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n656), .A2(new_n657), .ZN(new_n665));
  INV_X1    g240(.A(new_n652), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n660), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G2096), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(G2100), .A3(new_n661), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT84), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n678), .A2(KEYINPUT85), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(KEYINPUT85), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n673), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n682), .B2(new_n673), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n675), .B(KEYINPUT19), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n677), .A2(new_n684), .A3(new_n682), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n683), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1981), .B(G1986), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n683), .A2(new_n688), .A3(new_n690), .A4(new_n687), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n672), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(new_n671), .A3(new_n696), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  XNOR2_X1  g278(.A(KEYINPUT89), .B(G16), .ZN(new_n704));
  MUX2_X1   g279(.A(G24), .B(G290), .S(new_n704), .Z(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(G1986), .Z(new_n706));
  INV_X1    g281(.A(G25), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT86), .B1(new_n707), .B2(G29), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n707), .A2(KEYINPUT86), .A3(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n487), .A2(G131), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT87), .ZN(new_n711));
  NOR2_X1   g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT88), .Z(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n484), .A2(G119), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n708), .B(new_n709), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT35), .B(G1991), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n719), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G6), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G305), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT32), .B(G1981), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n728), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  INV_X1    g309(.A(new_n704), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n735), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT94), .B(G1971), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G23), .ZN(new_n740));
  NAND2_X1  g315(.A1(G288), .A2(KEYINPUT92), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n578), .A2(new_n580), .A3(new_n742), .A4(new_n579), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n740), .B1(new_n744), .B2(G16), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT93), .B(G1976), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT33), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n733), .A2(new_n734), .A3(new_n739), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n706), .B(new_n722), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT36), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n749), .B(new_n750), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n755), .A2(new_n756), .A3(new_n706), .A4(new_n722), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n718), .A2(G26), .ZN(new_n759));
  OAI221_X1 g334(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n472), .C2(G116), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n487), .A2(G140), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n481), .A2(new_n482), .A3(G128), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(new_n718), .ZN(new_n765));
  MUX2_X1   g340(.A(new_n759), .B(new_n765), .S(KEYINPUT28), .Z(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(KEYINPUT24), .A2(G34), .ZN(new_n769));
  NOR2_X1   g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n769), .A2(new_n770), .A3(G29), .ZN(new_n771));
  INV_X1    g346(.A(G160), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2084), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT96), .B(KEYINPUT25), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n472), .A2(new_n777), .A3(G103), .A4(G2104), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G115), .A2(G2104), .ZN(new_n782));
  INV_X1    g357(.A(G127), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n486), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(new_n482), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n487), .A2(G139), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n781), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  OR2_X1    g363(.A1(G29), .A2(G33), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n788), .A2(G2072), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n775), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT26), .Z(new_n793));
  NAND3_X1  g368(.A1(new_n481), .A2(new_n482), .A3(G129), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n481), .A2(G141), .A3(new_n461), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G29), .B2(G32), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT27), .B(G1996), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n788), .A2(new_n789), .ZN(new_n804));
  INV_X1    g379(.A(G2072), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g381(.A(KEYINPUT97), .B(G2072), .C1(new_n788), .C2(new_n789), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n791), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n791), .A2(KEYINPUT99), .A3(new_n802), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n774), .A2(G2084), .ZN(new_n814));
  AND2_X1   g389(.A1(KEYINPUT30), .A2(G28), .ZN(new_n815));
  NOR2_X1   g390(.A1(KEYINPUT30), .A2(G28), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n718), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n817), .B1(new_n629), .B2(new_n718), .C1(new_n800), .C2(new_n801), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT102), .B1(G5), .B2(G16), .ZN(new_n820));
  OR3_X1    g395(.A1(KEYINPUT102), .A2(G5), .A3(G16), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n820), .B(new_n821), .C1(G301), .C2(new_n723), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT103), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(G1961), .ZN(new_n824));
  NAND2_X1  g399(.A1(G168), .A2(G16), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G16), .B2(G21), .ZN(new_n826));
  INV_X1    g401(.A(G1966), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(G1961), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n819), .A2(new_n824), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(G27), .A2(G29), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G164), .B2(G29), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2078), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n830), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT100), .B(KEYINPUT31), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G11), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n813), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT104), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n842));
  INV_X1    g417(.A(G35), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G29), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(G29), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n489), .B2(G29), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n846), .B2(new_n842), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT29), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(G2090), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(G2090), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n735), .A2(KEYINPUT23), .A3(G20), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT23), .ZN(new_n852));
  INV_X1    g427(.A(G20), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n704), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n851), .B(new_n854), .C1(new_n576), .C2(new_n723), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G1956), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n723), .A2(G4), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n606), .B2(new_n723), .ZN(new_n858));
  INV_X1    g433(.A(G1348), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n735), .A2(G19), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n546), .B2(new_n735), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT95), .B(G1341), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NOR4_X1   g440(.A1(new_n849), .A2(new_n850), .A3(new_n856), .A4(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n813), .A2(new_n837), .A3(new_n867), .A4(new_n839), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n841), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n758), .A2(new_n768), .A3(new_n869), .ZN(G311));
  NAND3_X1  g445(.A1(new_n758), .A2(new_n869), .A3(new_n768), .ZN(G150));
  OR2_X1    g446(.A1(KEYINPUT106), .A2(G93), .ZN(new_n872));
  NAND2_X1  g447(.A1(KEYINPUT106), .A2(G93), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n519), .A2(new_n520), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n519), .A2(G55), .A3(G543), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n513), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n606), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g456(.A1(G68), .A2(G543), .ZN(new_n882));
  INV_X1    g457(.A(G56), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n582), .B2(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n884), .A2(G651), .B1(G43), .B2(new_n517), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n877), .A2(new_n885), .A3(new_n543), .ZN(new_n886));
  NAND2_X1  g461(.A1(G80), .A2(G543), .ZN(new_n887));
  INV_X1    g462(.A(G67), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n582), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n889), .A2(G651), .B1(G55), .B2(new_n517), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n545), .A2(new_n890), .A3(new_n874), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT39), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n881), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n879), .B1(new_n894), .B2(G860), .ZN(G145));
  XNOR2_X1  g470(.A(new_n489), .B(new_n772), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n484), .A2(G130), .B1(G142), .B2(new_n487), .ZN(new_n897));
  OAI221_X1 g472(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n472), .C2(G118), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n619), .B(new_n899), .Z(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n787), .A2(KEYINPUT107), .A3(new_n503), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n763), .B(new_n797), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n781), .A2(KEYINPUT107), .A3(new_n785), .A4(new_n786), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n495), .A3(new_n507), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n902), .B2(new_n905), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n907), .A2(new_n908), .A3(new_n716), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n902), .A2(new_n905), .ZN(new_n910));
  INV_X1    g485(.A(new_n903), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n717), .B1(new_n912), .B2(new_n906), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n901), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n716), .B1(new_n907), .B2(new_n908), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n717), .A3(new_n906), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n900), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n629), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n914), .A2(new_n915), .A3(new_n629), .A4(new_n918), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n896), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n922), .A3(new_n896), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g503(.A1(G72), .A2(G543), .ZN(new_n929));
  INV_X1    g504(.A(G60), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(new_n582), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G651), .ZN(new_n932));
  NAND4_X1  g507(.A1(G303), .A2(new_n594), .A3(new_n932), .A4(new_n593), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n518), .A2(new_n521), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n522), .A2(new_n513), .ZN(new_n935));
  NAND3_X1  g510(.A1(G290), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n744), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n744), .B1(new_n936), .B2(new_n933), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n938), .A2(new_n939), .A3(G305), .ZN(new_n940));
  INV_X1    g515(.A(G305), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(new_n936), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n741), .A2(new_n743), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n944), .B2(new_n937), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n940), .B2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(G305), .B1(new_n938), .B2(new_n939), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n944), .A2(new_n941), .A3(new_n937), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(KEYINPUT109), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n947), .B1(KEYINPUT42), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n614), .B(new_n892), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n606), .B1(new_n562), .B2(new_n575), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n557), .A2(new_n559), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT77), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n557), .A2(KEYINPUT77), .A3(new_n559), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n575), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n955), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n956), .A2(KEYINPUT41), .A3(new_n964), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT41), .B1(new_n956), .B2(new_n964), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n955), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n954), .B(new_n970), .ZN(new_n971));
  MUX2_X1   g546(.A(new_n877), .B(new_n971), .S(G868), .Z(G295));
  MUX2_X1   g547(.A(new_n877), .B(new_n971), .S(G868), .Z(G331));
  NAND2_X1  g548(.A1(G286), .A2(G171), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n528), .A2(new_n530), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT74), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n528), .A2(KEYINPUT74), .A3(new_n530), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n979), .A2(new_n526), .A3(new_n527), .A4(G301), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n886), .B2(new_n891), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n886), .A2(new_n891), .A3(new_n982), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n981), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n892), .A2(KEYINPUT110), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(new_n984), .A3(new_n974), .A4(new_n980), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n965), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n967), .A2(KEYINPUT113), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT41), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n963), .B1(new_n961), .B2(new_n962), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n956), .A2(KEYINPUT41), .A3(new_n964), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n991), .B1(new_n997), .B2(KEYINPUT113), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n990), .B1(new_n998), .B2(new_n989), .ZN(new_n999));
  INV_X1    g574(.A(new_n953), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT111), .B1(new_n969), .B2(new_n989), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n997), .A2(new_n1003), .A3(new_n988), .A4(new_n986), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1002), .A2(new_n953), .A3(new_n990), .A4(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1005), .A2(KEYINPUT112), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(KEYINPUT112), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n925), .B(new_n1001), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n969), .A2(new_n989), .A3(KEYINPUT111), .ZN(new_n1011));
  AND4_X1   g586(.A1(new_n987), .A2(new_n984), .A3(new_n974), .A4(new_n980), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n987), .A2(new_n984), .B1(new_n980), .B2(new_n974), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1003), .B1(new_n1014), .B2(new_n997), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n953), .A4(new_n990), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1005), .A2(KEYINPUT112), .ZN(new_n1019));
  AOI21_X1  g594(.A(G37), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n990), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1000), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT43), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT44), .B1(new_n1010), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1009), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(G397));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  INV_X1    g606(.A(G40), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n469), .A2(new_n475), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n507), .B2(new_n495), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n507), .A2(new_n508), .A3(new_n495), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n508), .B1(new_n507), .B2(new_n495), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(G1384), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1031), .B(new_n1037), .C1(new_n1040), .C2(new_n1036), .ZN(new_n1041));
  INV_X1    g616(.A(G1384), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n503), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n504), .A2(new_n1042), .A3(new_n509), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT114), .B(G1971), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT55), .Z(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1030), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n589), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1035), .B2(new_n1033), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1055), .A2(G1981), .A3(new_n1059), .A4(new_n1056), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1066), .B2(new_n943), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT52), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT52), .B(new_n1067), .C1(new_n1066), .C2(G288), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1046), .A2(new_n1044), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1048), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1062), .B1(new_n1076), .B2(new_n1041), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(KEYINPUT115), .A3(new_n1052), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1054), .A2(new_n1071), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1080), .A2(G288), .B1(G1981), .B2(G305), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1063), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1033), .B1(new_n1043), .B2(KEYINPUT50), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(KEYINPUT50), .B2(new_n1046), .ZN(new_n1085));
  INV_X1    g660(.A(G2084), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1034), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n1042), .A4(new_n509), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1085), .A2(new_n1086), .B1(new_n1089), .B2(new_n827), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G286), .A2(G8), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(new_n1091), .C1(new_n1090), .C2(new_n1062), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1089), .A2(new_n827), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n1086), .A3(new_n1037), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT51), .B(G8), .C1(new_n1098), .C2(G286), .ZN(new_n1099));
  AOI211_X1 g674(.A(KEYINPUT62), .B(new_n1092), .C1(new_n1094), .C2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1048), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1034), .B1(new_n1043), .B2(KEYINPUT50), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1046), .B2(KEYINPUT50), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n1104));
  AOI21_X1  g679(.A(G2090), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1102), .B(KEYINPUT117), .C1(new_n1046), .C2(KEYINPUT50), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1053), .B1(new_n1107), .B2(new_n1062), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT115), .B1(new_n1077), .B2(new_n1052), .ZN(new_n1109));
  AND4_X1   g684(.A1(KEYINPUT115), .A2(new_n1049), .A3(G8), .A4(new_n1052), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1108), .B(new_n1071), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1100), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n1089), .B2(G2078), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  INV_X1    g689(.A(G2078), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1087), .A2(new_n1088), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1113), .A2(KEYINPUT53), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1072), .A2(new_n1115), .A3(new_n1073), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1096), .A2(new_n1037), .ZN(new_n1121));
  INV_X1    g696(.A(G1961), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G171), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1092), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(KEYINPUT62), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1083), .B1(new_n1112), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n503), .A2(new_n1042), .A3(new_n1033), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT118), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1035), .A2(new_n1133), .A3(new_n1033), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n767), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n767), .A4(new_n1134), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1121), .A2(new_n859), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  INV_X1    g717(.A(G1956), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1047), .A2(new_n1142), .B1(new_n1103), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT57), .B1(new_n557), .B2(new_n559), .ZN(new_n1145));
  AOI22_X1  g720(.A1(G299), .A2(KEYINPUT57), .B1(new_n962), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1141), .A2(new_n1147), .A3(new_n606), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1348), .B1(new_n1096), .B2(new_n1037), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n963), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1140), .A2(new_n606), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1156));
  INV_X1    g731(.A(G1996), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(new_n1073), .C1(new_n1040), .C2(KEYINPUT45), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT58), .B(G1341), .Z(new_n1159));
  INV_X1    g734(.A(new_n1134), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1133), .B1(new_n1035), .B2(new_n1033), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1156), .B1(new_n1163), .B2(new_n546), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1156), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n545), .B(new_n1165), .C1(new_n1158), .C2(new_n1162), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1139), .A2(new_n1168), .A3(new_n606), .A4(new_n1140), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1147), .A2(KEYINPUT61), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1155), .A2(new_n1167), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT121), .B1(new_n1147), .B2(KEYINPUT61), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1144), .A2(new_n1173), .A3(new_n1174), .A4(new_n1146), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1150), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1111), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n1117), .A2(new_n1124), .A3(G171), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1118), .A2(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1035), .A2(KEYINPUT45), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n469), .A2(KEYINPUT123), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT53), .B1(new_n1185), .B2(new_n1115), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1184), .A2(new_n475), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(G40), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n469), .B2(KEYINPUT123), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1182), .A2(new_n1183), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1181), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1180), .B1(new_n1191), .B2(G171), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1179), .A2(new_n1192), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1120), .A2(new_n1123), .A3(G301), .A4(new_n1190), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1181), .A2(KEYINPUT125), .A3(G301), .A4(new_n1190), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1125), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1180), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1177), .A2(new_n1178), .A3(new_n1193), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1090), .A2(new_n1062), .A3(G286), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1201), .B1(new_n1111), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1054), .A2(new_n1078), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1205), .A2(new_n1071), .A3(new_n1202), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1130), .A2(new_n1200), .A3(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1182), .A2(new_n1034), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n764), .A2(new_n767), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n763), .A2(G2067), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n797), .B(new_n1157), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n720), .B2(new_n716), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n717), .A2(new_n721), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g793(.A(G290), .B(G1986), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1210), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1209), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1210), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1222), .A2(G1986), .A3(G290), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1223), .B(KEYINPUT48), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1224), .B1(new_n1210), .B2(new_n1218), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1222), .A2(G1996), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1226), .B1(new_n1227), .B2(KEYINPUT46), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1213), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1210), .B1(new_n1229), .B2(new_n797), .ZN(new_n1230));
  XNOR2_X1  g805(.A(KEYINPUT126), .B(KEYINPUT46), .ZN(new_n1231));
  OAI211_X1 g806(.A(new_n1228), .B(new_n1230), .C1(new_n1226), .C2(new_n1231), .ZN(new_n1232));
  XOR2_X1   g807(.A(new_n1232), .B(KEYINPUT47), .Z(new_n1233));
  OAI21_X1  g808(.A(new_n1211), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1234));
  AOI211_X1 g809(.A(new_n1225), .B(new_n1233), .C1(new_n1210), .C2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1221), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g811(.A(new_n459), .B1(new_n699), .B2(new_n701), .ZN(new_n1238));
  AND3_X1   g812(.A1(new_n664), .A2(new_n645), .A3(new_n669), .ZN(new_n1239));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1240));
  AND3_X1   g814(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g815(.A(new_n1240), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1242));
  NOR2_X1   g816(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AND3_X1   g817(.A1(new_n921), .A2(new_n922), .A3(new_n896), .ZN(new_n1244));
  NOR3_X1   g818(.A1(new_n1244), .A2(new_n923), .A3(G37), .ZN(new_n1245));
  NAND2_X1  g819(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1246));
  NAND2_X1  g820(.A1(new_n1246), .A2(KEYINPUT43), .ZN(new_n1247));
  NAND3_X1  g821(.A1(new_n1020), .A2(new_n1009), .A3(new_n1001), .ZN(new_n1248));
  AOI211_X1 g822(.A(new_n1243), .B(new_n1245), .C1(new_n1247), .C2(new_n1248), .ZN(G308));
  OAI221_X1 g823(.A(new_n927), .B1(new_n1242), .B2(new_n1241), .C1(new_n1026), .C2(new_n1027), .ZN(G225));
endmodule


