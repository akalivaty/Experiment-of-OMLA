

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  NOR2_X1 U324 ( .A1(n584), .A2(n419), .ZN(n421) );
  NOR2_X1 U325 ( .A1(n531), .A2(n482), .ZN(n564) );
  XNOR2_X1 U326 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U327 ( .A(n456), .B(n455), .ZN(n507) );
  XOR2_X1 U328 ( .A(n372), .B(n371), .Z(n531) );
  XOR2_X1 U329 ( .A(G183GAT), .B(KEYINPUT18), .Z(n292) );
  XNOR2_X1 U330 ( .A(n424), .B(KEYINPUT69), .ZN(n425) );
  XNOR2_X1 U331 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U332 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U333 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U334 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U335 ( .A(n406), .B(KEYINPUT99), .ZN(n407) );
  NOR2_X1 U336 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U337 ( .A(n365), .B(n364), .ZN(n370) );
  XNOR2_X1 U338 ( .A(n408), .B(n407), .ZN(n568) );
  XNOR2_X1 U339 ( .A(KEYINPUT38), .B(KEYINPUT108), .ZN(n455) );
  XNOR2_X1 U340 ( .A(n436), .B(n435), .ZN(n574) );
  XNOR2_X1 U341 ( .A(n403), .B(n402), .ZN(n522) );
  XNOR2_X1 U342 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U343 ( .A(n461), .B(G43GAT), .ZN(n462) );
  XNOR2_X1 U344 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT3), .B(KEYINPUT89), .Z(n294) );
  XNOR2_X1 U347 ( .A(KEYINPUT88), .B(G155GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U349 ( .A(KEYINPUT2), .B(n295), .Z(n377) );
  XOR2_X1 U350 ( .A(G85GAT), .B(G162GAT), .Z(n297) );
  XNOR2_X1 U351 ( .A(G29GAT), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U353 ( .A(KEYINPUT1), .B(n298), .Z(n300) );
  NAND2_X1 U354 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n377), .B(n301), .ZN(n319) );
  XOR2_X1 U357 ( .A(KEYINPUT96), .B(KEYINPUT93), .Z(n303) );
  XNOR2_X1 U358 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U360 ( .A(G57GAT), .B(G148GAT), .Z(n305) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(G1GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n317) );
  XOR2_X1 U364 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n309) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G127GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U367 ( .A(G134GAT), .B(KEYINPUT81), .Z(n310) );
  XOR2_X1 U368 ( .A(n311), .B(n310), .Z(n371) );
  INV_X1 U369 ( .A(n371), .ZN(n315) );
  XOR2_X1 U370 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n313) );
  XNOR2_X1 U371 ( .A(KEYINPUT5), .B(KEYINPUT95), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U373 ( .A(n315), .B(n314), .Z(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U375 ( .A(n319), .B(n318), .Z(n547) );
  INV_X1 U376 ( .A(n547), .ZN(n566) );
  XNOR2_X1 U377 ( .A(KEYINPUT105), .B(KEYINPUT36), .ZN(n336) );
  XOR2_X1 U378 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n321) );
  XNOR2_X1 U379 ( .A(KEYINPUT72), .B(KEYINPUT11), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n327) );
  XOR2_X1 U381 ( .A(G29GAT), .B(G43GAT), .Z(n323) );
  XNOR2_X1 U382 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n444) );
  XOR2_X1 U384 ( .A(G92GAT), .B(n444), .Z(n325) );
  NAND2_X1 U385 ( .A1(G232GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n335) );
  XOR2_X1 U388 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n329) );
  XNOR2_X1 U389 ( .A(G134GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .ZN(n433) );
  XNOR2_X1 U392 ( .A(n330), .B(n433), .ZN(n333) );
  XOR2_X1 U393 ( .A(G50GAT), .B(G162GAT), .Z(n373) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G190GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n331), .B(G218GAT), .ZN(n396) );
  XNOR2_X1 U396 ( .A(n373), .B(n396), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U398 ( .A(n335), .B(n334), .Z(n560) );
  INV_X1 U399 ( .A(n560), .ZN(n491) );
  XOR2_X1 U400 ( .A(n336), .B(n491), .Z(n584) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XOR2_X1 U402 ( .A(G211GAT), .B(G78GAT), .Z(n338) );
  XNOR2_X1 U403 ( .A(G71GAT), .B(G155GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U405 ( .A(G127GAT), .B(G183GAT), .Z(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n358) );
  XOR2_X1 U408 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n344) );
  XNOR2_X1 U409 ( .A(KEYINPUT74), .B(KEYINPUT14), .ZN(n343) );
  XNOR2_X1 U410 ( .A(n344), .B(n343), .ZN(n356) );
  XOR2_X1 U411 ( .A(KEYINPUT79), .B(G64GAT), .Z(n346) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(G22GAT), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U414 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n348) );
  XNOR2_X1 U415 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n347) );
  XNOR2_X1 U416 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U417 ( .A(n350), .B(n349), .Z(n354) );
  XNOR2_X1 U418 ( .A(G15GAT), .B(G1GAT), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n351), .B(KEYINPUT66), .ZN(n439) );
  XNOR2_X1 U420 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n352), .B(KEYINPUT67), .ZN(n429) );
  XNOR2_X1 U422 ( .A(n439), .B(n429), .ZN(n353) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U424 ( .A(n356), .B(n355), .Z(n357) );
  XOR2_X1 U425 ( .A(n358), .B(n357), .Z(n471) );
  XOR2_X1 U426 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U427 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n359) );
  XNOR2_X1 U428 ( .A(n292), .B(n359), .ZN(n394) );
  XOR2_X1 U429 ( .A(n434), .B(n394), .Z(n365) );
  XOR2_X1 U430 ( .A(G176GAT), .B(G15GAT), .Z(n361) );
  NAND2_X1 U431 ( .A1(G227GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U432 ( .A(n361), .B(n360), .ZN(n363) );
  XNOR2_X1 U433 ( .A(G43GAT), .B(G99GAT), .ZN(n362) );
  XOR2_X1 U434 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n367) );
  XNOR2_X1 U435 ( .A(G190GAT), .B(KEYINPUT84), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U437 ( .A(G169GAT), .B(n368), .Z(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U439 ( .A(G204GAT), .B(G218GAT), .Z(n375) );
  XOR2_X1 U440 ( .A(G141GAT), .B(G22GAT), .Z(n440) );
  XNOR2_X1 U441 ( .A(n440), .B(n373), .ZN(n374) );
  XOR2_X1 U442 ( .A(n375), .B(n374), .Z(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n379) );
  AND2_X1 U444 ( .A1(G228GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U446 ( .A(G106GAT), .B(G78GAT), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n380), .B(G148GAT), .ZN(n426) );
  XNOR2_X1 U448 ( .A(n381), .B(n426), .ZN(n383) );
  XNOR2_X1 U449 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n391) );
  XOR2_X1 U451 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n385) );
  XNOR2_X1 U452 ( .A(KEYINPUT87), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U454 ( .A(G197GAT), .B(n386), .Z(n398) );
  XOR2_X1 U455 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n388) );
  XNOR2_X1 U456 ( .A(KEYINPUT85), .B(KEYINPUT24), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n398), .B(n389), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n479) );
  XOR2_X1 U460 ( .A(n479), .B(KEYINPUT28), .Z(n527) );
  XOR2_X1 U461 ( .A(G64GAT), .B(G92GAT), .Z(n393) );
  XNOR2_X1 U462 ( .A(G176GAT), .B(G204GAT), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n393), .B(n392), .ZN(n430) );
  XNOR2_X1 U464 ( .A(n394), .B(n430), .ZN(n403) );
  XOR2_X1 U465 ( .A(G169GAT), .B(G8GAT), .Z(n447) );
  XOR2_X1 U466 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n395) );
  XOR2_X1 U467 ( .A(n447), .B(n399), .Z(n401) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U470 ( .A(n522), .B(KEYINPUT27), .Z(n405) );
  NAND2_X1 U471 ( .A1(n527), .A2(n405), .ZN(n404) );
  NOR2_X1 U472 ( .A1(n566), .A2(n404), .ZN(n533) );
  NAND2_X1 U473 ( .A1(n531), .A2(n533), .ZN(n417) );
  INV_X1 U474 ( .A(n405), .ZN(n409) );
  AND2_X1 U475 ( .A1(n479), .A2(n531), .ZN(n408) );
  XNOR2_X1 U476 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n406) );
  NOR2_X1 U477 ( .A1(n409), .A2(n568), .ZN(n548) );
  XNOR2_X1 U478 ( .A(n548), .B(KEYINPUT101), .ZN(n414) );
  NOR2_X1 U479 ( .A1(n531), .A2(n522), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n410), .B(KEYINPUT102), .ZN(n411) );
  NOR2_X1 U481 ( .A1(n479), .A2(n411), .ZN(n412) );
  XNOR2_X1 U482 ( .A(KEYINPUT25), .B(n412), .ZN(n413) );
  NAND2_X1 U483 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U484 ( .A1(n415), .A2(n566), .ZN(n416) );
  NAND2_X1 U485 ( .A1(n417), .A2(n416), .ZN(n494) );
  NAND2_X1 U486 ( .A1(n471), .A2(n494), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n418), .B(KEYINPUT106), .ZN(n419) );
  XNOR2_X1 U488 ( .A(KEYINPUT37), .B(KEYINPUT107), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n520) );
  XOR2_X1 U490 ( .A(KEYINPUT68), .B(KEYINPUT33), .Z(n423) );
  XNOR2_X1 U491 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n422) );
  XNOR2_X1 U492 ( .A(n423), .B(n422), .ZN(n428) );
  AND2_X1 U493 ( .A1(G230GAT), .A2(G233GAT), .ZN(n424) );
  XOR2_X1 U494 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U497 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n438) );
  XNOR2_X1 U498 ( .A(G113GAT), .B(G197GAT), .ZN(n437) );
  XOR2_X1 U499 ( .A(n438), .B(n437), .Z(n452) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n443), .B(KEYINPUT64), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n444), .B(KEYINPUT30), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U507 ( .A(G50GAT), .B(G36GAT), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n464) );
  INV_X1 U510 ( .A(n464), .ZN(n453) );
  INV_X1 U511 ( .A(n453), .ZN(n570) );
  NAND2_X1 U512 ( .A1(n574), .A2(n570), .ZN(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT70), .B(n454), .Z(n496) );
  NAND2_X1 U514 ( .A1(n520), .A2(n496), .ZN(n456) );
  NOR2_X1 U515 ( .A1(n566), .A2(n507), .ZN(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT109), .B(KEYINPUT39), .ZN(n458) );
  INV_X1 U517 ( .A(G29GAT), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  NOR2_X1 U520 ( .A1(n531), .A2(n507), .ZN(n463) );
  INV_X1 U521 ( .A(KEYINPUT40), .ZN(n461) );
  INV_X1 U522 ( .A(n471), .ZN(n579) );
  XOR2_X1 U523 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n466) );
  XOR2_X1 U524 ( .A(KEYINPUT41), .B(n574), .Z(n509) );
  INV_X1 U525 ( .A(n509), .ZN(n483) );
  NAND2_X1 U526 ( .A1(n483), .A2(n464), .ZN(n465) );
  XOR2_X1 U527 ( .A(n466), .B(n465), .Z(n467) );
  NOR2_X1 U528 ( .A1(n579), .A2(n467), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT114), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n469), .A2(n491), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT47), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n584), .A2(n471), .ZN(n472) );
  XNOR2_X1 U533 ( .A(KEYINPUT45), .B(n472), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n473), .A2(n574), .ZN(n474) );
  NOR2_X1 U535 ( .A1(n474), .A2(n570), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT48), .ZN(n550) );
  NOR2_X1 U537 ( .A1(n522), .A2(n550), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT54), .B(n478), .ZN(n567) );
  NOR2_X1 U539 ( .A1(n479), .A2(n547), .ZN(n480) );
  AND2_X1 U540 ( .A1(n567), .A2(n480), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n564), .A2(n483), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G176GAT), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1349GAT) );
  NAND2_X1 U546 ( .A1(n564), .A2(n560), .ZN(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n488) );
  XNOR2_X1 U548 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n487) );
  XOR2_X1 U549 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n493) );
  NAND2_X1 U550 ( .A1(n579), .A2(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n495) );
  AND2_X1 U552 ( .A1(n495), .A2(n494), .ZN(n510) );
  NAND2_X1 U553 ( .A1(n510), .A2(n496), .ZN(n504) );
  NOR2_X1 U554 ( .A1(n566), .A2(n504), .ZN(n498) );
  XNOR2_X1 U555 ( .A(KEYINPUT34), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  NOR2_X1 U558 ( .A1(n522), .A2(n504), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(n500), .Z(n501) );
  XNOR2_X1 U560 ( .A(G8GAT), .B(n501), .ZN(G1325GAT) );
  NOR2_X1 U561 ( .A1(n531), .A2(n504), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  NOR2_X1 U564 ( .A1(n527), .A2(n504), .ZN(n505) );
  XOR2_X1 U565 ( .A(G22GAT), .B(n505), .Z(G1327GAT) );
  NOR2_X1 U566 ( .A1(n522), .A2(n507), .ZN(n506) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U568 ( .A1(n527), .A2(n507), .ZN(n508) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NOR2_X1 U570 ( .A1(n570), .A2(n509), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n519), .A2(n510), .ZN(n516) );
  NOR2_X1 U572 ( .A1(n566), .A2(n516), .ZN(n511) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n516), .ZN(n513) );
  XOR2_X1 U576 ( .A(KEYINPUT110), .B(n513), .Z(n514) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n531), .A2(n516), .ZN(n515) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n515), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n527), .A2(n516), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U584 ( .A1(n566), .A2(n526), .ZN(n521) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n526), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n531), .A2(n526), .ZN(n525) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  INV_X1 U595 ( .A(n531), .ZN(n532) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U597 ( .A1(n550), .A2(n534), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n570), .A2(n543), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U601 ( .A1(n543), .A2(n483), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n542) );
  XOR2_X1 U605 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U606 ( .A1(n543), .A2(n579), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U610 ( .A1(n543), .A2(n560), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n570), .A2(n559), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n553) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(n554), .Z(n556) );
  NAND2_X1 U621 ( .A1(n559), .A2(n483), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT121), .Z(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n579), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n570), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n579), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n569) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n580) );
  NAND2_X1 U636 ( .A1(n580), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  INV_X1 U639 ( .A(n580), .ZN(n583) );
  NOR2_X1 U640 ( .A1(n583), .A2(n574), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT127), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

