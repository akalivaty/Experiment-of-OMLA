//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  INV_X1    g036(.A(G2106), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n455), .B2(new_n462), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT68), .Z(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n468), .B1(new_n471), .B2(G137), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n465), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n467), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n478), .A2(KEYINPUT69), .B1(G113), .B2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G125), .C1(new_n473), .C2(new_n474), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n465), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n477), .A2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n471), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n465), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n484), .B1(new_n485), .B2(new_n486), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT71), .ZN(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n473), .B2(new_n474), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT72), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(new_n495), .C1(new_n473), .C2(new_n474), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n465), .C1(new_n473), .C2(new_n474), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n488), .A2(new_n503), .A3(G138), .A4(new_n465), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT73), .B(G651), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n511), .A2(new_n512), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G88), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n521), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(G543), .B1(new_n530), .B2(new_n519), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n518), .B(new_n524), .C1(new_n525), .C2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n522), .A2(G89), .A3(new_n523), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n522), .A2(G51), .A3(G543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G168));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n547), .B(new_n548), .C1(new_n513), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n549), .B1(new_n511), .B2(new_n512), .ZN(new_n551));
  INV_X1    g126(.A(new_n548), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT75), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n517), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n522), .A2(G90), .A3(new_n523), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n531), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT76), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n531), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G52), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n561), .A2(new_n554), .A3(new_n562), .A4(new_n556), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G171));
  AOI22_X1  g139(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n516), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n522), .A2(G81), .A3(new_n523), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n522), .A2(G43), .A3(G543), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  OAI211_X1 g151(.A(G91), .B(new_n523), .C1(new_n530), .C2(new_n519), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n522), .A2(new_n579), .A3(G91), .A4(new_n523), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g156(.A(G53), .B(G543), .C1(new_n530), .C2(new_n519), .ZN(new_n582));
  XOR2_X1   g157(.A(KEYINPUT78), .B(KEYINPUT9), .Z(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT9), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n522), .A2(G53), .A3(G543), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G78), .A2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT80), .ZN(new_n590));
  INV_X1    g165(.A(G65), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n513), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n581), .A2(new_n588), .A3(new_n593), .ZN(G299));
  INV_X1    g169(.A(G171), .ZN(G301));
  NAND2_X1  g170(.A1(new_n545), .A2(KEYINPUT81), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n542), .A2(new_n543), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n597), .A2(new_n598), .A3(new_n544), .A4(new_n541), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G286));
  NAND3_X1  g176(.A1(new_n522), .A2(G49), .A3(G543), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n522), .A2(G87), .A3(new_n523), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G288));
  OAI211_X1 g180(.A(G48), .B(G543), .C1(new_n530), .C2(new_n519), .ZN(new_n606));
  OAI211_X1 g181(.A(G86), .B(new_n523), .C1(new_n530), .C2(new_n519), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n511), .B2(new_n512), .ZN(new_n609));
  AND2_X1   g184(.A1(G73), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n517), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(G305));
  NAND3_X1  g187(.A1(new_n522), .A2(G85), .A3(new_n523), .ZN(new_n613));
  INV_X1    g188(.A(G47), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n531), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT82), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(new_n516), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(G290));
  OAI211_X1 g194(.A(G92), .B(new_n523), .C1(new_n530), .C2(new_n519), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  INV_X1    g198(.A(G66), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n513), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n560), .A2(G54), .B1(G651), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G868), .B2(G171), .ZN(G284));
  XNOR2_X1  g204(.A(G284), .B(KEYINPUT83), .ZN(G321));
  NOR2_X1   g205(.A1(G299), .A2(G868), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n600), .ZN(G297));
  AOI21_X1  g207(.A(new_n631), .B1(G868), .B2(new_n600), .ZN(G280));
  INV_X1    g208(.A(new_n627), .ZN(new_n634));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G860), .ZN(G148));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n569), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n627), .A2(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(new_n637), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n488), .A2(new_n466), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT13), .Z(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT84), .B(G2100), .ZN(new_n645));
  INV_X1    g220(.A(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n471), .A2(G135), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  INV_X1    g225(.A(G111), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(G2105), .ZN(new_n652));
  INV_X1    g227(.A(new_n489), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(G123), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI22_X1  g231(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(G2096), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n657), .B(new_n658), .C1(new_n645), .C2(new_n644), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT86), .Z(G156));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n662), .B(new_n664), .Z(new_n665));
  INV_X1    g240(.A(KEYINPUT14), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT87), .B(G2438), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2427), .B(G2430), .Z(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n670), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n665), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(G14), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT89), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G401));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT17), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT90), .B(G2100), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2072), .B(G2078), .Z(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n683), .B2(KEYINPUT18), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(new_n646), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1971), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n696), .B2(new_n702), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT92), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(new_n708), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n712), .B1(new_n709), .B2(new_n713), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n694), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n718), .A2(new_n693), .A3(new_n714), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n717), .A2(new_n719), .ZN(G229));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G33), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT25), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n488), .A2(G127), .ZN(new_n725));
  NAND2_X1  g300(.A1(G115), .A2(G2104), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n465), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n724), .B(new_n727), .C1(G139), .C2(new_n471), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n722), .B1(new_n728), .B2(new_n721), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G2072), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT102), .Z(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G28), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT104), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(new_n721), .C1(new_n733), .C2(G28), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n732), .B(new_n736), .C1(new_n655), .C2(new_n721), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n729), .B2(G2072), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n471), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  INV_X1    g316(.A(G129), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n741), .C1(new_n742), .C2(new_n489), .ZN(new_n743));
  MUX2_X1   g318(.A(G32), .B(new_n743), .S(G29), .Z(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT103), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n744), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n731), .A2(new_n738), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n634), .A2(G16), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G4), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(G1348), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n748), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n721), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT100), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n653), .A2(G128), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT99), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n465), .A2(G116), .ZN(new_n761));
  OAI21_X1  g336(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n471), .A2(G140), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT98), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n758), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT101), .B(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G160), .A2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(KEYINPUT24), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n721), .A2(G27), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n721), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2078), .ZN(new_n781));
  INV_X1    g356(.A(G16), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n782), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1966), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n781), .B(new_n785), .C1(new_n776), .C2(new_n775), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n755), .A2(new_n778), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G5), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G171), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1961), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G19), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n570), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT97), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1341), .ZN(new_n795));
  INV_X1    g370(.A(G2090), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n721), .A2(G35), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT105), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G162), .B2(new_n721), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT29), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n782), .A2(G20), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT23), .Z(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G299), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1956), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n801), .B2(new_n796), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT106), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n791), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n811));
  NAND2_X1  g386(.A1(G303), .A2(G16), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n782), .A2(G22), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT94), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G23), .B(G288), .S(G16), .Z(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT33), .B(G1976), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n812), .A2(new_n814), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G1971), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n817), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(G305), .A2(new_n782), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n828));
  OR2_X1    g403(.A1(G6), .A2(G16), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g406(.A(G1981), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT32), .ZN(new_n834));
  INV_X1    g409(.A(G1981), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n811), .B1(new_n826), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n817), .A2(new_n820), .A3(new_n825), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n832), .A2(new_n837), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT95), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n810), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n782), .A2(G24), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT93), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n616), .A2(new_n618), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n782), .ZN(new_n848));
  INV_X1    g423(.A(G1986), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n721), .A2(G25), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n653), .A2(G119), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n471), .A2(G131), .ZN(new_n853));
  OR2_X1    g428(.A1(G95), .A2(G2105), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n854), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n851), .B1(new_n857), .B2(new_n721), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G1991), .Z(new_n859));
  XOR2_X1   g434(.A(new_n858), .B(new_n859), .Z(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n850), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n843), .A2(new_n844), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n826), .A2(new_n811), .A3(new_n838), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT95), .B1(new_n840), .B2(new_n841), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT34), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n850), .A2(new_n861), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT96), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT34), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT36), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT36), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n809), .B1(new_n872), .B2(new_n874), .ZN(G311));
  AND3_X1   g450(.A1(new_n791), .A2(new_n802), .A3(new_n808), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n869), .A2(new_n873), .A3(new_n870), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n869), .B2(new_n870), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(G150));
  NOR2_X1   g454(.A1(new_n627), .A2(new_n635), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n522), .A2(G93), .A3(new_n523), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT107), .B(G55), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n882), .B1(new_n516), .B2(new_n883), .C1(new_n531), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n569), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n881), .B(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(G860), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(G860), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT37), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n890), .A2(new_n892), .ZN(G145));
  NAND2_X1  g468(.A1(new_n471), .A2(G142), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n897));
  INV_X1    g472(.A(G118), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(G2105), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(new_n653), .B2(G130), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT109), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n643), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n901), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n643), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n728), .B(new_n743), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n903), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n764), .A2(G164), .A3(new_n766), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G164), .B1(new_n764), .B2(new_n766), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n857), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(new_n856), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G162), .B(G160), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(new_n656), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n910), .A2(new_n917), .A3(new_n919), .A4(new_n912), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n923), .B1(new_n921), .B2(new_n924), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(KEYINPUT110), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n930), .B(new_n923), .C1(new_n921), .C2(new_n924), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g508(.A1(new_n847), .A2(G305), .ZN(new_n934));
  XNOR2_X1  g509(.A(G303), .B(G288), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n616), .A2(G305), .A3(new_n618), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n935), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n847), .A2(G305), .ZN(new_n939));
  INV_X1    g514(.A(new_n936), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n570), .B(new_n885), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(new_n639), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n634), .A2(G299), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n584), .A2(new_n587), .B1(G651), .B2(new_n592), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n627), .A2(new_n581), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n634), .A2(KEYINPUT111), .A3(G299), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT41), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n945), .A2(new_n947), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n952), .A2(KEYINPUT41), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n944), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n949), .A2(new_n950), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n886), .B(new_n639), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n954), .A2(new_n957), .A3(KEYINPUT42), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n951), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n956), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n949), .A2(new_n950), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n944), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n959), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n942), .B1(new_n958), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT42), .B1(new_n954), .B2(new_n957), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n959), .A3(new_n963), .ZN(new_n967));
  INV_X1    g542(.A(new_n942), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G868), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n885), .A2(new_n637), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n637), .B1(new_n965), .B2(new_n969), .ZN(new_n975));
  INV_X1    g550(.A(new_n973), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT112), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(G295));
  NAND2_X1  g553(.A1(new_n971), .A2(new_n973), .ZN(G331));
  AOI22_X1  g554(.A1(new_n596), .A2(new_n599), .B1(new_n559), .B2(new_n563), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n559), .A2(new_n545), .A3(new_n563), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n886), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n600), .A2(G171), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n559), .A2(new_n545), .A3(new_n563), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n943), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n984), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT113), .A3(new_n886), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n952), .A2(KEYINPUT41), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT114), .B(new_n886), .C1(new_n980), .C2(new_n981), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n985), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT114), .B1(new_n988), .B2(new_n886), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n962), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT41), .B(new_n991), .C1(new_n993), .C2(new_n994), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n968), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n987), .A2(new_n951), .A3(new_n953), .A4(new_n989), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n982), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n955), .A2(new_n1002), .A3(new_n985), .A4(new_n992), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n942), .A3(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1004), .A2(new_n926), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n999), .A2(new_n1005), .A3(KEYINPUT43), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n926), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n942), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT44), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n999), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1017), .ZN(G397));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G1384), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n506), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT117), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1022), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n500), .B2(new_n505), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1384), .B1(new_n500), .B2(new_n505), .ZN(new_n1030));
  OAI211_X1 g605(.A(G160), .B(G40), .C1(KEYINPUT45), .C2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n813), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1384), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n506), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G113), .A2(G2104), .ZN(new_n1037));
  INV_X1    g612(.A(G125), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n469), .B2(new_n470), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1039), .B2(new_n480), .ZN(new_n1040));
  INV_X1    g615(.A(new_n481), .ZN(new_n1041));
  OAI21_X1  g616(.A(G2105), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n471), .A2(new_n468), .A3(G137), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1043), .A2(new_n1044), .B1(G101), .B2(new_n466), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1042), .A2(new_n1045), .A3(G40), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1030), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1036), .A2(new_n796), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1020), .B1(new_n1032), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1019), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1020), .B1(new_n1046), .B2(new_n1030), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n606), .A2(new_n607), .A3(new_n835), .A4(new_n611), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1057), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1046), .A2(new_n1030), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n602), .A2(new_n603), .A3(G1976), .A4(new_n604), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1063), .A2(G8), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1042), .A2(new_n1045), .A3(G40), .ZN(new_n1068));
  OAI211_X1 g643(.A(G8), .B(new_n1064), .C1(new_n1068), .C2(new_n1034), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT52), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1062), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  AOI211_X1 g646(.A(G1384), .B(new_n1035), .C1(new_n500), .C2(new_n505), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n1068), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1034), .A2(KEYINPUT50), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n796), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1020), .B1(new_n1032), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1071), .B1(new_n1076), .B2(new_n1053), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1027), .B1(new_n506), .B2(new_n1022), .ZN(new_n1078));
  AOI211_X1 g653(.A(KEYINPUT117), .B(new_n1025), .C1(new_n500), .C2(new_n505), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT45), .B1(new_n506), .B2(new_n1033), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n1068), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1971), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1049), .ZN(new_n1084));
  OAI21_X1  g659(.A(G8), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(KEYINPUT119), .A3(new_n1052), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1966), .B1(new_n1082), .B2(new_n1023), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1030), .A2(new_n1047), .ZN(new_n1088));
  NOR4_X1   g663(.A1(new_n1088), .A2(new_n1072), .A3(new_n1068), .A4(G2084), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n600), .A2(G8), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1054), .A2(new_n1077), .A3(new_n1086), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT120), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1090), .A2(new_n1094), .A3(new_n1091), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1077), .B(new_n1099), .C1(new_n1053), .C2(new_n1076), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1076), .A2(new_n1053), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1055), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1057), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G288), .A2(G1976), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1062), .B2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1102), .A2(new_n1071), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n545), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1035), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1030), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1074), .A2(new_n776), .A3(new_n1046), .A4(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1081), .A2(new_n1068), .A3(new_n1026), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1112), .B(G168), .C1(new_n1113), .C2(G1966), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1109), .A2(G8), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1114), .A2(new_n1117), .A3(G8), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1108), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G2078), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1080), .A2(new_n1082), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1124));
  INV_X1    g699(.A(G1961), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1113), .A2(KEYINPUT53), .A3(new_n1121), .ZN(new_n1127));
  AOI21_X1  g702(.A(G301), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1054), .A2(new_n1077), .A3(new_n1086), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1120), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1118), .B1(KEYINPUT51), .B2(new_n1115), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1108), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1107), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT121), .B(G1956), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(G160), .B(G40), .C1(new_n1030), .C2(new_n1110), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1048), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT56), .B(G2072), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1080), .A2(new_n1082), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT57), .B1(new_n588), .B2(KEYINPUT122), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G299), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n584), .B2(new_n587), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n946), .B(new_n581), .C1(new_n1144), .C2(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1138), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1138), .A2(new_n1140), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1152));
  INV_X1    g727(.A(G2067), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1068), .A2(new_n1034), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1124), .A2(new_n751), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1152), .A2(new_n1146), .B1(new_n627), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1156), .A3(KEYINPUT124), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1146), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1151), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(KEYINPUT126), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1148), .A2(new_n1150), .B1(new_n1163), .B2(new_n1162), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1169), .B2(KEYINPUT61), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(G1996), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1080), .A2(new_n1082), .A3(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(KEYINPUT58), .B(G1341), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1154), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n570), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(KEYINPUT125), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n627), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1177), .A2(KEYINPUT125), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1175), .A2(new_n570), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n627), .B1(new_n1155), .B2(KEYINPUT60), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(KEYINPUT60), .B2(new_n1155), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1164), .A2(KEYINPUT61), .A3(new_n1147), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1161), .B1(new_n1171), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT54), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1068), .A2(new_n1123), .A3(G2078), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT115), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1021), .B1(new_n1030), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1080), .B(new_n1192), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  AND4_X1   g771(.A1(G301), .A2(new_n1190), .A3(new_n1191), .A4(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1189), .B1(new_n1197), .B2(new_n1128), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(KEYINPUT127), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1200), .B(new_n1189), .C1(new_n1197), .C2(new_n1128), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1190), .A2(new_n1191), .A3(new_n1196), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(G171), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1126), .A2(G301), .A3(new_n1127), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1204), .A2(KEYINPUT54), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1054), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1206), .A2(new_n1207), .A3(new_n1131), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1101), .B(new_n1133), .C1(new_n1188), .C2(new_n1209), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1195), .A2(new_n1194), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1211), .A2(new_n1068), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n767), .A2(G2067), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n764), .A2(new_n1153), .A3(new_n766), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n743), .B(new_n1172), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n856), .B(new_n859), .Z(new_n1217));
  OAI21_X1  g792(.A(new_n1212), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1212), .ZN(new_n1219));
  XNOR2_X1  g794(.A(G290), .B(new_n849), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT116), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1210), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1212), .B1(new_n1224), .B2(new_n743), .ZN(new_n1225));
  NOR3_X1   g800(.A1(new_n1219), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT46), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1227), .B1(new_n1212), .B2(new_n1172), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1225), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1229), .B(KEYINPUT47), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1219), .A2(G1986), .A3(G290), .ZN(new_n1231));
  OR2_X1    g806(.A1(new_n1231), .A2(KEYINPUT48), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(KEYINPUT48), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1232), .A2(new_n1218), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n857), .A2(new_n859), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1214), .B1(new_n1216), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1212), .ZN(new_n1237));
  AND3_X1   g812(.A1(new_n1230), .A2(new_n1234), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1223), .A2(new_n1238), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g814(.A1(G227), .A2(new_n463), .ZN(new_n1241));
  NAND2_X1  g815(.A1(new_n678), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g816(.A(new_n1242), .B1(new_n717), .B2(new_n719), .ZN(new_n1243));
  NAND3_X1  g817(.A1(new_n1243), .A2(new_n1015), .A3(new_n932), .ZN(G225));
  INV_X1    g818(.A(G225), .ZN(G308));
endmodule


