

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G651), .A2(n539), .ZN(n649) );
  INV_X1 U554 ( .A(n719), .ZN(n720) );
  NAND2_X1 U555 ( .A1(n688), .A2(n781), .ZN(n719) );
  BUF_X1 U556 ( .A(n562), .Z(n523) );
  NOR2_X2 U557 ( .A1(n736), .A2(n735), .ZN(n741) );
  NOR2_X1 U558 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U559 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U560 ( .A(n752), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U561 ( .A1(G8), .A2(n719), .ZN(n775) );
  NOR2_X2 U562 ( .A1(n536), .A2(n539), .ZN(n590) );
  XOR2_X1 U563 ( .A(n729), .B(KEYINPUT28), .Z(n521) );
  NOR2_X1 U564 ( .A1(n775), .A2(n757), .ZN(n522) );
  XNOR2_X2 U565 ( .A(n570), .B(KEYINPUT65), .ZN(G160) );
  INV_X1 U566 ( .A(n1001), .ZN(n707) );
  XNOR2_X1 U567 ( .A(KEYINPUT30), .B(KEYINPUT100), .ZN(n692) );
  XNOR2_X1 U568 ( .A(n693), .B(n692), .ZN(n694) );
  INV_X1 U569 ( .A(KEYINPUT13), .ZN(n594) );
  XNOR2_X1 U570 ( .A(n594), .B(KEYINPUT71), .ZN(n595) );
  XNOR2_X1 U571 ( .A(n596), .B(n595), .ZN(n597) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n651) );
  INV_X1 U573 ( .A(KEYINPUT104), .ZN(n815) );
  XOR2_X1 U574 ( .A(KEYINPUT15), .B(n610), .Z(n1004) );
  AND2_X1 U575 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U576 ( .A(G2104), .ZN(n526) );
  NOR2_X1 U577 ( .A1(G2105), .A2(n526), .ZN(n562) );
  NAND2_X1 U578 ( .A1(G99), .A2(n523), .ZN(n525) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n981) );
  NAND2_X1 U580 ( .A1(G111), .A2(n981), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n525), .A2(n524), .ZN(n529) );
  AND2_X1 U582 ( .A1(n526), .A2(G2105), .ZN(n980) );
  NAND2_X1 U583 ( .A1(n980), .A2(G123), .ZN(n527) );
  XOR2_X1 U584 ( .A(KEYINPUT18), .B(n527), .Z(n528) );
  NOR2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n532) );
  NOR2_X2 U586 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XOR2_X2 U587 ( .A(KEYINPUT17), .B(n530), .Z(n984) );
  NAND2_X1 U588 ( .A1(n984), .A2(G135), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n974) );
  XNOR2_X1 U590 ( .A(G2096), .B(n974), .ZN(n533) );
  OR2_X1 U591 ( .A1(G2100), .A2(n533), .ZN(G156) );
  INV_X1 U592 ( .A(G651), .ZN(n536) );
  NOR2_X1 U593 ( .A1(G543), .A2(n536), .ZN(n534) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n534), .Z(n650) );
  NAND2_X1 U595 ( .A1(G65), .A2(n650), .ZN(n538) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n535) );
  XNOR2_X1 U597 ( .A(KEYINPUT68), .B(n535), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G78), .A2(n590), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G91), .A2(n651), .ZN(n541) );
  NAND2_X1 U601 ( .A1(G53), .A2(n649), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n727) );
  INV_X1 U604 ( .A(n727), .ZN(G299) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  INV_X1 U606 ( .A(G132), .ZN(G219) );
  INV_X1 U607 ( .A(G82), .ZN(G220) );
  NAND2_X1 U608 ( .A1(G52), .A2(n649), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n544), .B(KEYINPUT69), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G77), .A2(n590), .ZN(n546) );
  NAND2_X1 U611 ( .A1(G90), .A2(n651), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NAND2_X1 U614 ( .A1(G64), .A2(n650), .ZN(n548) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(G171) );
  INV_X1 U617 ( .A(G171), .ZN(G301) );
  NAND2_X1 U618 ( .A1(G114), .A2(n981), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G126), .A2(n980), .ZN(n553) );
  NAND2_X1 U620 ( .A1(G138), .A2(n984), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n562), .A2(G102), .ZN(n554) );
  XOR2_X1 U623 ( .A(KEYINPUT88), .B(n554), .Z(n555) );
  NOR2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT89), .ZN(G164) );
  NAND2_X1 U627 ( .A1(G125), .A2(n980), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n984), .A2(G137), .ZN(n560) );
  AND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT23), .B(KEYINPUT67), .Z(n564) );
  NAND2_X1 U631 ( .A1(G101), .A2(n562), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(KEYINPUT66), .ZN(n567) );
  AND2_X1 U634 ( .A1(n981), .A2(G113), .ZN(n566) );
  NOR2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n650), .A2(G63), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT77), .B(n571), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n649), .A2(G51), .ZN(n572) );
  XOR2_X1 U640 ( .A(n572), .B(KEYINPUT78), .Z(n573) );
  NOR2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT6), .B(n575), .Z(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(KEYINPUT79), .ZN(n584) );
  XOR2_X1 U644 ( .A(KEYINPUT4), .B(KEYINPUT76), .Z(n578) );
  NAND2_X1 U645 ( .A1(G89), .A2(n651), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U647 ( .A(KEYINPUT75), .B(n579), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n590), .A2(G76), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT5), .B(n582), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n585), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U653 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U654 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U656 ( .A(G223), .ZN(n845) );
  NAND2_X1 U657 ( .A1(n845), .A2(G567), .ZN(n587) );
  XOR2_X1 U658 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  NAND2_X1 U659 ( .A1(n650), .A2(G56), .ZN(n588) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n588), .Z(n598) );
  NAND2_X1 U661 ( .A1(n651), .A2(G81), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT12), .B(n589), .Z(n593) );
  NAND2_X1 U663 ( .A1(n590), .A2(G68), .ZN(n591) );
  XOR2_X1 U664 ( .A(n591), .B(KEYINPUT70), .Z(n592) );
  NOR2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U667 ( .A(n599), .B(KEYINPUT72), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G43), .A2(n649), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n1001) );
  INV_X1 U670 ( .A(G860), .ZN(n616) );
  OR2_X1 U671 ( .A1(n1001), .A2(n616), .ZN(n602) );
  XOR2_X1 U672 ( .A(KEYINPUT73), .B(n602), .Z(G153) );
  NAND2_X1 U673 ( .A1(G868), .A2(G301), .ZN(n612) );
  NAND2_X1 U674 ( .A1(n649), .A2(G54), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G79), .A2(n590), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G92), .A2(n651), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n650), .A2(G66), .ZN(n605) );
  XOR2_X1 U679 ( .A(KEYINPUT74), .B(n605), .Z(n606) );
  NOR2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n610) );
  INV_X1 U682 ( .A(G868), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n1004), .A2(n613), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(G284) );
  NOR2_X1 U685 ( .A1(G286), .A2(n613), .ZN(n615) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n616), .A2(G559), .ZN(n617) );
  INV_X1 U689 ( .A(n1004), .ZN(n661) );
  NAND2_X1 U690 ( .A1(n617), .A2(n661), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G868), .A2(n1001), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n661), .A2(G868), .ZN(n619) );
  NOR2_X1 U694 ( .A1(G559), .A2(n619), .ZN(n620) );
  NOR2_X1 U695 ( .A1(n621), .A2(n620), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G75), .A2(n590), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G88), .A2(n651), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n650), .A2(G62), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT84), .B(n624), .Z(n625) );
  NOR2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n649), .A2(G50), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(G303) );
  INV_X1 U704 ( .A(G303), .ZN(G166) );
  NAND2_X1 U705 ( .A1(G73), .A2(n590), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U707 ( .A1(G61), .A2(n650), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G48), .A2(n649), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G86), .A2(n651), .ZN(n632) );
  XNOR2_X1 U711 ( .A(KEYINPUT83), .B(n632), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(G305) );
  AND2_X1 U714 ( .A1(n650), .A2(G60), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G72), .A2(n590), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G85), .A2(n651), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n649), .A2(G47), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U721 ( .A1(n539), .A2(G87), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n643), .B(KEYINPUT82), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G49), .A2(n649), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U726 ( .A1(n650), .A2(n646), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U728 ( .A1(G55), .A2(n649), .ZN(n658) );
  NAND2_X1 U729 ( .A1(G67), .A2(n650), .ZN(n653) );
  NAND2_X1 U730 ( .A1(G93), .A2(n651), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n590), .A2(G80), .ZN(n654) );
  XOR2_X1 U733 ( .A(KEYINPUT80), .B(n654), .Z(n655) );
  NOR2_X1 U734 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n659), .B(KEYINPUT81), .ZN(n970) );
  NOR2_X1 U737 ( .A1(G868), .A2(n970), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n660), .B(KEYINPUT87), .ZN(n672) );
  NAND2_X1 U739 ( .A1(G559), .A2(n661), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n1001), .B(n662), .ZN(n969) );
  XOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n664) );
  XNOR2_X1 U742 ( .A(G166), .B(KEYINPUT85), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n727), .B(n665), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(G305), .ZN(n668) );
  XOR2_X1 U746 ( .A(G290), .B(G288), .Z(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n970), .B(n669), .ZN(n1002) );
  XOR2_X1 U749 ( .A(n969), .B(n1002), .Z(n670) );
  NAND2_X1 U750 ( .A1(G868), .A2(n670), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U760 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G96), .A2(n679), .ZN(n967) );
  NAND2_X1 U762 ( .A1(n967), .A2(G2106), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U764 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U765 ( .A1(G108), .A2(n681), .ZN(n968) );
  NAND2_X1 U766 ( .A1(n968), .A2(G567), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n972) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U769 ( .A1(n972), .A2(n684), .ZN(n848) );
  NAND2_X1 U770 ( .A1(n848), .A2(G36), .ZN(G176) );
  NOR2_X1 U771 ( .A1(G1971), .A2(G303), .ZN(n685) );
  XNOR2_X1 U772 ( .A(n685), .B(KEYINPUT103), .ZN(n756) );
  NOR2_X1 U773 ( .A1(G1976), .A2(G288), .ZN(n912) );
  NAND2_X1 U774 ( .A1(G40), .A2(G160), .ZN(n686) );
  XNOR2_X1 U775 ( .A(KEYINPUT90), .B(n686), .ZN(n780) );
  XNOR2_X1 U776 ( .A(n780), .B(KEYINPUT95), .ZN(n688) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n687) );
  XNOR2_X1 U778 ( .A(KEYINPUT64), .B(n687), .ZN(n781) );
  NOR2_X1 U779 ( .A1(G2084), .A2(n719), .ZN(n690) );
  NAND2_X1 U780 ( .A1(G8), .A2(n690), .ZN(n689) );
  XOR2_X1 U781 ( .A(KEYINPUT96), .B(n689), .Z(n740) );
  NOR2_X1 U782 ( .A1(G1966), .A2(n775), .ZN(n737) );
  NOR2_X1 U783 ( .A1(n737), .A2(n690), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G8), .A2(n691), .ZN(n693) );
  NOR2_X1 U785 ( .A1(n694), .A2(G168), .ZN(n699) );
  INV_X1 U786 ( .A(n719), .ZN(n722) );
  XOR2_X1 U787 ( .A(G1961), .B(KEYINPUT97), .Z(n945) );
  NOR2_X1 U788 ( .A1(n722), .A2(n945), .ZN(n695) );
  XNOR2_X1 U789 ( .A(n695), .B(KEYINPUT98), .ZN(n697) );
  XOR2_X1 U790 ( .A(G2078), .B(KEYINPUT25), .Z(n895) );
  NOR2_X1 U791 ( .A1(n719), .A2(n895), .ZN(n696) );
  NOR2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n732) );
  AND2_X1 U793 ( .A1(G301), .A2(n732), .ZN(n698) );
  XNOR2_X1 U794 ( .A(n700), .B(KEYINPUT31), .ZN(n736) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n719), .ZN(n702) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n722), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n1004), .A2(n703), .ZN(n718) );
  NAND2_X1 U799 ( .A1(n1004), .A2(G2067), .ZN(n705) );
  XOR2_X1 U800 ( .A(KEYINPUT26), .B(KEYINPUT99), .Z(n714) );
  NAND2_X1 U801 ( .A1(G1996), .A2(n714), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n706), .A2(n722), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U805 ( .A1(G1348), .A2(n1004), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n714), .A2(n709), .ZN(n710) );
  NOR2_X1 U807 ( .A1(G1341), .A2(n710), .ZN(n711) );
  NOR2_X1 U808 ( .A1(n722), .A2(n711), .ZN(n712) );
  OR2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n714), .ZN(n715) );
  NOR2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n720), .A2(G2072), .ZN(n721) );
  XNOR2_X1 U814 ( .A(n721), .B(KEYINPUT27), .ZN(n724) );
  INV_X1 U815 ( .A(G1956), .ZN(n936) );
  NOR2_X1 U816 ( .A1(n936), .A2(n722), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n521), .ZN(n731) );
  XNOR2_X1 U821 ( .A(n731), .B(KEYINPUT29), .ZN(n734) );
  NOR2_X1 U822 ( .A1(G301), .A2(n732), .ZN(n733) );
  NOR2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U824 ( .A1(n737), .A2(n741), .ZN(n738) );
  XNOR2_X1 U825 ( .A(n738), .B(KEYINPUT101), .ZN(n739) );
  NOR2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n754) );
  INV_X1 U827 ( .A(n741), .ZN(n743) );
  AND2_X1 U828 ( .A1(G286), .A2(G8), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n751) );
  INV_X1 U830 ( .A(G8), .ZN(n749) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n775), .ZN(n745) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n719), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n746), .A2(G303), .ZN(n747) );
  XNOR2_X1 U835 ( .A(n747), .B(KEYINPUT102), .ZN(n748) );
  OR2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U838 ( .A1(n754), .A2(n753), .ZN(n763) );
  NOR2_X1 U839 ( .A1(n912), .A2(n763), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n756), .A2(n755), .ZN(n762) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n913) );
  INV_X1 U842 ( .A(n913), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n912), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U844 ( .A1(n758), .A2(n775), .ZN(n760) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n929) );
  INV_X1 U846 ( .A(n929), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n765) );
  AND2_X1 U848 ( .A1(n522), .A2(n765), .ZN(n761) );
  AND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n779) );
  INV_X1 U850 ( .A(n763), .ZN(n768) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G8), .A2(n764), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n765), .A2(KEYINPUT33), .ZN(n769) );
  AND2_X1 U854 ( .A1(n766), .A2(n769), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n772) );
  INV_X1 U856 ( .A(n769), .ZN(n770) );
  OR2_X1 U857 ( .A1(n770), .A2(n775), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n777) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n773) );
  XOR2_X1 U860 ( .A(n773), .B(KEYINPUT24), .Z(n774) );
  OR2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n814) );
  NOR2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n830) );
  INV_X1 U865 ( .A(n830), .ZN(n812) );
  NAND2_X1 U866 ( .A1(G119), .A2(n980), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G131), .A2(n984), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G95), .A2(n523), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G107), .A2(n981), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n995) );
  NAND2_X1 U873 ( .A1(G1991), .A2(n995), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(KEYINPUT92), .ZN(n799) );
  NAND2_X1 U875 ( .A1(G141), .A2(n984), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n789), .B(KEYINPUT94), .ZN(n797) );
  NAND2_X1 U877 ( .A1(n523), .A2(G105), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n790), .B(KEYINPUT38), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G129), .A2(n980), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G117), .A2(n981), .ZN(n793) );
  XNOR2_X1 U882 ( .A(KEYINPUT93), .B(n793), .ZN(n794) );
  NOR2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n977) );
  NAND2_X1 U885 ( .A1(G1996), .A2(n977), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n860) );
  XOR2_X1 U887 ( .A(G1986), .B(G290), .Z(n918) );
  NAND2_X1 U888 ( .A1(G128), .A2(n980), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G116), .A2(n981), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n802), .B(KEYINPUT35), .ZN(n808) );
  XNOR2_X1 U892 ( .A(KEYINPUT91), .B(KEYINPUT34), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G104), .A2(n523), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G140), .A2(n984), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U896 ( .A(n806), .B(n805), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U898 ( .A(KEYINPUT36), .B(n809), .ZN(n998) );
  XOR2_X1 U899 ( .A(G2067), .B(KEYINPUT37), .Z(n817) );
  NAND2_X1 U900 ( .A1(n998), .A2(n817), .ZN(n818) );
  NAND2_X1 U901 ( .A1(n918), .A2(n818), .ZN(n810) );
  NOR2_X1 U902 ( .A1(n860), .A2(n810), .ZN(n811) );
  NOR2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U905 ( .A(n816), .B(n815), .ZN(n833) );
  NOR2_X1 U906 ( .A1(n998), .A2(n817), .ZN(n861) );
  INV_X1 U907 ( .A(n818), .ZN(n879) );
  XOR2_X1 U908 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n819) );
  XNOR2_X1 U909 ( .A(KEYINPUT108), .B(n819), .ZN(n826) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n977), .ZN(n820) );
  XOR2_X1 U911 ( .A(KEYINPUT105), .B(n820), .Z(n858) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n995), .ZN(n876) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n876), .A2(n821), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT106), .ZN(n823) );
  NOR2_X1 U916 ( .A1(n860), .A2(n823), .ZN(n824) );
  NOR2_X1 U917 ( .A1(n858), .A2(n824), .ZN(n825) );
  XOR2_X1 U918 ( .A(n826), .B(n825), .Z(n827) );
  NOR2_X1 U919 ( .A1(n879), .A2(n827), .ZN(n828) );
  NOR2_X1 U920 ( .A1(n861), .A2(n828), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT109), .B(n829), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U924 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U925 ( .A(G2443), .B(G1348), .ZN(n843) );
  XNOR2_X1 U926 ( .A(G2430), .B(G2435), .ZN(n841) );
  XOR2_X1 U927 ( .A(KEYINPUT110), .B(G2454), .Z(n836) );
  XNOR2_X1 U928 ( .A(G2427), .B(G2451), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U930 ( .A(n837), .B(G2446), .Z(n839) );
  XNOR2_X1 U931 ( .A(G1341), .B(G2438), .ZN(n838) );
  XNOR2_X1 U932 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U933 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U934 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U935 ( .A1(n844), .A2(G14), .ZN(n1028) );
  XNOR2_X1 U936 ( .A(KEYINPUT111), .B(n1028), .ZN(G401) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U939 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(G188) );
  NAND2_X1 U943 ( .A1(G124), .A2(n980), .ZN(n849) );
  XNOR2_X1 U944 ( .A(n849), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U945 ( .A1(G112), .A2(n981), .ZN(n850) );
  XOR2_X1 U946 ( .A(KEYINPUT115), .B(n850), .Z(n851) );
  NAND2_X1 U947 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U948 ( .A1(G100), .A2(n523), .ZN(n854) );
  NAND2_X1 U949 ( .A1(G136), .A2(n984), .ZN(n853) );
  NAND2_X1 U950 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U951 ( .A1(n856), .A2(n855), .ZN(G162) );
  XOR2_X1 U952 ( .A(G2090), .B(G162), .Z(n857) );
  NOR2_X1 U953 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT51), .B(n859), .Z(n863) );
  NOR2_X1 U955 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U956 ( .A1(n863), .A2(n862), .ZN(n884) );
  XNOR2_X1 U957 ( .A(KEYINPUT50), .B(KEYINPUT121), .ZN(n874) );
  NAND2_X1 U958 ( .A1(G103), .A2(n523), .ZN(n865) );
  NAND2_X1 U959 ( .A1(G139), .A2(n984), .ZN(n864) );
  NAND2_X1 U960 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U961 ( .A1(G127), .A2(n980), .ZN(n867) );
  NAND2_X1 U962 ( .A1(G115), .A2(n981), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U964 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U965 ( .A1(n870), .A2(n869), .ZN(n975) );
  XNOR2_X1 U966 ( .A(G2072), .B(n975), .ZN(n872) );
  XNOR2_X1 U967 ( .A(G164), .B(G2078), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n874), .B(n873), .ZN(n882) );
  XOR2_X1 U970 ( .A(G160), .B(G2084), .Z(n875) );
  NOR2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n877) );
  NAND2_X1 U972 ( .A1(n877), .A2(n974), .ZN(n878) );
  NOR2_X1 U973 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U974 ( .A(n880), .B(KEYINPUT120), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U976 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U977 ( .A(KEYINPUT52), .B(n885), .ZN(n886) );
  INV_X1 U978 ( .A(KEYINPUT55), .ZN(n908) );
  NAND2_X1 U979 ( .A1(n886), .A2(n908), .ZN(n887) );
  NAND2_X1 U980 ( .A1(n887), .A2(G29), .ZN(n965) );
  XNOR2_X1 U981 ( .A(G2084), .B(KEYINPUT54), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n888), .B(G34), .ZN(n903) );
  XNOR2_X1 U983 ( .A(G1991), .B(G25), .ZN(n893) );
  XNOR2_X1 U984 ( .A(G2067), .B(G26), .ZN(n890) );
  XNOR2_X1 U985 ( .A(G2072), .B(G33), .ZN(n889) );
  NOR2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(KEYINPUT123), .B(n891), .ZN(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G28), .A2(n894), .ZN(n900) );
  XNOR2_X1 U990 ( .A(G1996), .B(G32), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n895), .B(G27), .ZN(n896) );
  NOR2_X1 U992 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U993 ( .A(KEYINPUT124), .B(n898), .Z(n899) );
  NOR2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(KEYINPUT53), .ZN(n902) );
  NOR2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n906) );
  XOR2_X1 U997 ( .A(G2090), .B(KEYINPUT122), .Z(n904) );
  XNOR2_X1 U998 ( .A(G35), .B(n904), .ZN(n905) );
  NAND2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n910) );
  INV_X1 U1001 ( .A(G29), .ZN(n909) );
  NAND2_X1 U1002 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(G11), .A2(n911), .ZN(n963) );
  XNOR2_X1 U1004 ( .A(G16), .B(KEYINPUT56), .ZN(n935) );
  INV_X1 U1005 ( .A(n912), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(n914), .A2(n913), .ZN(n920) );
  XNOR2_X1 U1007 ( .A(G299), .B(G1956), .ZN(n916) );
  XNOR2_X1 U1008 ( .A(G303), .B(G1971), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(n920), .A2(n919), .ZN(n924) );
  XNOR2_X1 U1012 ( .A(G301), .B(G1961), .ZN(n922) );
  XNOR2_X1 U1013 ( .A(n1004), .B(G1348), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1016 ( .A(G1341), .B(n1001), .Z(n925) );
  XNOR2_X1 U1017 ( .A(KEYINPUT125), .B(n925), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(KEYINPUT126), .B(n928), .ZN(n933) );
  XNOR2_X1 U1020 ( .A(G1966), .B(G168), .ZN(n930) );
  NAND2_X1 U1021 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1022 ( .A(KEYINPUT57), .B(n931), .ZN(n932) );
  NAND2_X1 U1023 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1024 ( .A1(n935), .A2(n934), .ZN(n961) );
  INV_X1 U1025 ( .A(G16), .ZN(n959) );
  XNOR2_X1 U1026 ( .A(G20), .B(n936), .ZN(n940) );
  XNOR2_X1 U1027 ( .A(G1341), .B(G19), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(G1981), .B(G6), .ZN(n937) );
  NOR2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1030 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1031 ( .A(KEYINPUT59), .B(G1348), .Z(n941) );
  XNOR2_X1 U1032 ( .A(G4), .B(n941), .ZN(n942) );
  NOR2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1034 ( .A(KEYINPUT60), .B(n944), .ZN(n949) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G21), .ZN(n947) );
  XNOR2_X1 U1036 ( .A(n945), .B(G5), .ZN(n946) );
  NOR2_X1 U1037 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1038 ( .A1(n949), .A2(n948), .ZN(n956) );
  XNOR2_X1 U1039 ( .A(G1986), .B(G24), .ZN(n951) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G22), .ZN(n950) );
  NOR2_X1 U1041 ( .A1(n951), .A2(n950), .ZN(n953) );
  XOR2_X1 U1042 ( .A(G1976), .B(G23), .Z(n952) );
  NAND2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(KEYINPUT58), .B(n954), .ZN(n955) );
  NOR2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1046 ( .A(KEYINPUT61), .B(n957), .ZN(n958) );
  NAND2_X1 U1047 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1048 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1049 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1050 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1051 ( .A(KEYINPUT62), .B(n966), .Z(G311) );
  XNOR2_X1 U1052 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1053 ( .A(G120), .ZN(G236) );
  INV_X1 U1054 ( .A(G96), .ZN(G221) );
  INV_X1 U1055 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1056 ( .A1(n968), .A2(n967), .ZN(G325) );
  INV_X1 U1057 ( .A(G325), .ZN(G261) );
  NOR2_X1 U1058 ( .A1(n969), .A2(G860), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(n971), .B(n970), .ZN(G145) );
  INV_X1 U1060 ( .A(n972), .ZN(G319) );
  XOR2_X1 U1061 ( .A(G164), .B(G162), .Z(n973) );
  XNOR2_X1 U1062 ( .A(n974), .B(n973), .ZN(n979) );
  XOR2_X1 U1063 ( .A(G160), .B(n975), .Z(n976) );
  XNOR2_X1 U1064 ( .A(n977), .B(n976), .ZN(n978) );
  XNOR2_X1 U1065 ( .A(n979), .B(n978), .ZN(n997) );
  XOR2_X1 U1066 ( .A(KEYINPUT117), .B(KEYINPUT48), .Z(n993) );
  NAND2_X1 U1067 ( .A1(G130), .A2(n980), .ZN(n983) );
  NAND2_X1 U1068 ( .A1(G118), .A2(n981), .ZN(n982) );
  NAND2_X1 U1069 ( .A1(n983), .A2(n982), .ZN(n990) );
  NAND2_X1 U1070 ( .A1(G106), .A2(n523), .ZN(n986) );
  NAND2_X1 U1071 ( .A1(G142), .A2(n984), .ZN(n985) );
  NAND2_X1 U1072 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1073 ( .A(KEYINPUT116), .B(n987), .Z(n988) );
  XNOR2_X1 U1074 ( .A(KEYINPUT45), .B(n988), .ZN(n989) );
  NOR2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1076 ( .A(n991), .B(KEYINPUT46), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(n993), .B(n992), .ZN(n994) );
  XNOR2_X1 U1078 ( .A(n995), .B(n994), .ZN(n996) );
  XNOR2_X1 U1079 ( .A(n997), .B(n996), .ZN(n999) );
  XNOR2_X1 U1080 ( .A(n999), .B(n998), .ZN(n1000) );
  NOR2_X1 U1081 ( .A1(G37), .A2(n1000), .ZN(G395) );
  XNOR2_X1 U1082 ( .A(G286), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1083 ( .A(n1003), .B(n1002), .ZN(n1006) );
  XOR2_X1 U1084 ( .A(n1004), .B(G171), .Z(n1005) );
  XNOR2_X1 U1085 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1086 ( .A1(G37), .A2(n1007), .ZN(G397) );
  XOR2_X1 U1087 ( .A(G2096), .B(KEYINPUT43), .Z(n1009) );
  XNOR2_X1 U1088 ( .A(G2067), .B(G2072), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(n1009), .B(n1008), .ZN(n1010) );
  XOR2_X1 U1090 ( .A(n1010), .B(G2678), .Z(n1012) );
  XNOR2_X1 U1091 ( .A(G2090), .B(KEYINPUT42), .ZN(n1011) );
  XNOR2_X1 U1092 ( .A(n1012), .B(n1011), .ZN(n1016) );
  XOR2_X1 U1093 ( .A(KEYINPUT112), .B(G2100), .Z(n1014) );
  XNOR2_X1 U1094 ( .A(G2078), .B(G2084), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(n1016), .B(n1015), .ZN(G227) );
  XOR2_X1 U1097 ( .A(G2474), .B(G1976), .Z(n1018) );
  XNOR2_X1 U1098 ( .A(G1991), .B(G1956), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(n1018), .B(n1017), .ZN(n1019) );
  XOR2_X1 U1100 ( .A(n1019), .B(KEYINPUT41), .Z(n1021) );
  XNOR2_X1 U1101 ( .A(G1996), .B(G1961), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(n1021), .B(n1020), .ZN(n1025) );
  XOR2_X1 U1103 ( .A(KEYINPUT113), .B(G1971), .Z(n1023) );
  XNOR2_X1 U1104 ( .A(G1986), .B(G1966), .ZN(n1022) );
  XNOR2_X1 U1105 ( .A(n1023), .B(n1022), .ZN(n1024) );
  XOR2_X1 U1106 ( .A(n1025), .B(n1024), .Z(n1027) );
  XNOR2_X1 U1107 ( .A(G1981), .B(KEYINPUT114), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1027), .B(n1026), .ZN(G229) );
  NAND2_X1 U1109 ( .A1(n1028), .A2(G319), .ZN(n1029) );
  XNOR2_X1 U1110 ( .A(n1029), .B(KEYINPUT118), .ZN(n1032) );
  NOR2_X1 U1111 ( .A1(G395), .A2(G397), .ZN(n1030) );
  XNOR2_X1 U1112 ( .A(n1030), .B(KEYINPUT119), .ZN(n1031) );
  NOR2_X1 U1113 ( .A1(n1032), .A2(n1031), .ZN(n1035) );
  NOR2_X1 U1114 ( .A1(G227), .A2(G229), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(KEYINPUT49), .B(n1033), .Z(n1034) );
  NAND2_X1 U1116 ( .A1(n1035), .A2(n1034), .ZN(G225) );
  INV_X1 U1117 ( .A(G225), .ZN(G308) );
  INV_X1 U1118 ( .A(G108), .ZN(G238) );
endmodule

