//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  NAND2_X1  g001(.A1(G29gat), .A2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT91), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n214), .A3(KEYINPUT15), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(KEYINPUT90), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n206), .A2(new_n213), .A3(new_n218), .A4(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n210), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n212), .B1(new_n210), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n205), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT92), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(G1gat), .B2(new_n230), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI221_X1 g035(.A(new_n232), .B1(new_n233), .B2(new_n229), .C1(G1gat), .C2(new_n230), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n228), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n228), .B(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n241), .B2(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT93), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n202), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n238), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n228), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n244), .B(KEYINPUT13), .Z(new_n248));
  OR2_X1    g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n228), .B(KEYINPUT17), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n246), .ZN(new_n251));
  INV_X1    g050(.A(new_n244), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n251), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n245), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n255));
  XNOR2_X1  g054(.A(G169gat), .B(G197gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n245), .A2(new_n260), .A3(new_n249), .A4(new_n253), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(KEYINPUT94), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT94), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n254), .A2(new_n265), .A3(new_n261), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT95), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(KEYINPUT95), .A3(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G141gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT76), .B1(new_n272), .B2(G148gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n274));
  INV_X1    g073(.A(G148gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(G141gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n273), .B(new_n276), .C1(G141gat), .C2(new_n275), .ZN(new_n277));
  XNOR2_X1  g076(.A(G155gat), .B(G162gat), .ZN(new_n278));
  INV_X1    g077(.A(G155gat), .ZN(new_n279));
  INV_X1    g078(.A(G162gat), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT2), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n278), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(KEYINPUT2), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT22), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n291), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n292), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n290), .B(new_n291), .ZN(new_n301));
  INV_X1    g100(.A(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n289), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT83), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n282), .A2(new_n285), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n303), .B2(new_n300), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n304), .B2(new_n305), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n286), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n303), .A2(new_n315), .A3(new_n300), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n298), .B1(new_n292), .B2(new_n299), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n317), .B2(KEYINPUT81), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n307), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n304), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n310), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(KEYINPUT82), .A3(new_n310), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G22gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n321), .A2(KEYINPUT82), .A3(new_n310), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT82), .B1(new_n321), .B2(new_n310), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n312), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G22gat), .ZN(new_n332));
  XOR2_X1   g131(.A(G78gat), .B(G106gat), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT31), .ZN(new_n334));
  INV_X1    g133(.A(G50gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT84), .A4(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT84), .B1(new_n331), .B2(G22gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n336), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n331), .A2(G22gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n327), .B1(new_n341), .B2(new_n312), .ZN(new_n342));
  OAI22_X1  g141(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G120gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G113gat), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G120gat), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT1), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G134gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G127gat), .ZN(new_n354));
  INV_X1    g153(.A(G127gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n307), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(new_n354), .A3(new_n356), .A4(new_n287), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n357), .A2(KEYINPUT4), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n356), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n355), .B1(new_n350), .B2(new_n352), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n320), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n358), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n356), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n320), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n372), .A2(new_n374), .A3(new_n364), .A4(new_n361), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n373), .A2(new_n320), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n365), .B1(new_n376), .B2(new_n357), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(KEYINPUT5), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n378), .ZN(new_n387));
  INV_X1    g186(.A(new_n383), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n367), .A2(new_n378), .A3(KEYINPUT80), .A4(new_n383), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n386), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n388), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n395));
  INV_X1    g194(.A(G183gat), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT27), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT28), .ZN(new_n398));
  INV_X1    g197(.A(G190gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT27), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT64), .A3(G183gat), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n397), .A2(new_n398), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(KEYINPUT27), .B(G183gat), .Z(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(G190gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n404), .B2(new_n398), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT65), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G169gat), .ZN(new_n408));
  INV_X1    g207(.A(G176gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT66), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(KEYINPUT65), .B(new_n402), .C1(new_n404), .C2(new_n398), .ZN(new_n413));
  INV_X1    g212(.A(new_n410), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n414), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n407), .A2(new_n412), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(KEYINPUT24), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT23), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n408), .A3(new_n409), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n396), .A2(new_n399), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(KEYINPUT24), .A3(new_n417), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n422), .B(new_n424), .C1(new_n408), .C2(new_n409), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT25), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT74), .ZN(new_n429));
  INV_X1    g228(.A(G226gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n303), .A2(new_n300), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n432), .A2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n416), .A2(new_n427), .A3(new_n433), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n433), .B1(new_n416), .B2(new_n427), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n416), .A2(new_n427), .A3(new_n432), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT75), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT75), .ZN(new_n447));
  INV_X1    g246(.A(new_n443), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n434), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n437), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n446), .B(new_n447), .C1(new_n450), .C2(new_n436), .ZN(new_n451));
  XNOR2_X1  g250(.A(G8gat), .B(G36gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G64gat), .B(G92gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n445), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n446), .B1(new_n450), .B2(new_n436), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(KEYINPUT30), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n439), .B2(new_n444), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n337), .B(new_n343), .C1(new_n394), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n368), .A2(new_n369), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n416), .A2(new_n466), .A3(new_n427), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n416), .B2(new_n427), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n464), .B(new_n465), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT70), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n428), .A2(new_n373), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT70), .A3(new_n467), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n465), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT71), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT34), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n475), .B2(KEYINPUT34), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n473), .A2(G227gat), .A3(G233gat), .A4(new_n467), .ZN(new_n480));
  XNOR2_X1  g279(.A(G15gat), .B(G43gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G99gat), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT68), .B(G71gat), .Z(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT33), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(KEYINPUT32), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT69), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT69), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n480), .A2(new_n488), .A3(KEYINPUT32), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n480), .B1(KEYINPUT32), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n484), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n475), .A2(KEYINPUT34), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT71), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT34), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n487), .A2(new_n489), .B1(new_n492), .B2(new_n484), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n470), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n495), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n495), .B2(new_n501), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n463), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n364), .B1(new_n362), .B2(new_n363), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT39), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n388), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n363), .A2(new_n361), .A3(new_n359), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n365), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n376), .A2(new_n365), .A3(new_n357), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT39), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n514), .A2(KEYINPUT40), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT40), .B1(new_n514), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n462), .A2(new_n389), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n343), .A2(new_n337), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n457), .B1(new_n456), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n450), .A2(new_n436), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n435), .A2(new_n438), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(KEYINPUT37), .C1(new_n436), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(new_n459), .A3(new_n392), .A4(new_n393), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n445), .A2(new_n451), .A3(KEYINPUT37), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n526), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n522), .B(new_n523), .C1(new_n531), .C2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n463), .B(KEYINPUT85), .C1(new_n504), .C2(new_n508), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n511), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n337), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT84), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n326), .B2(new_n327), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n539), .A2(new_n336), .B1(new_n328), .B2(new_n332), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n495), .B(new_n501), .C1(new_n537), .C2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n455), .A2(new_n458), .A3(new_n461), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n392), .A2(new_n393), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n542), .A2(KEYINPUT35), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n523), .A2(new_n543), .A3(new_n495), .A4(new_n501), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n394), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n271), .B1(new_n536), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(G71gat), .A2(G78gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G57gat), .B(G64gat), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G64gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(G57gat), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G64gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n557), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n558), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n238), .B1(KEYINPUT21), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G183gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G211gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n572), .A2(new_n574), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n578), .B1(new_n575), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n552), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(new_n551), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(KEYINPUT97), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT8), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n590), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n592), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n593), .ZN(new_n599));
  NOR2_X1   g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g402(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n589), .B2(new_n590), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n601), .A2(new_n604), .A3(new_n592), .A4(new_n597), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n222), .B2(new_n227), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n250), .B2(new_n606), .ZN(new_n608));
  NAND3_X1  g407(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n588), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(KEYINPUT98), .A3(new_n611), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT96), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n614), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n588), .B(new_n622), .C1(new_n612), .C2(new_n613), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n587), .A2(KEYINPUT99), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n586), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n567), .A2(new_n603), .A3(new_n605), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT100), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n598), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n631), .A2(new_n604), .A3(new_n592), .A4(new_n597), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n567), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT101), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n634), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT101), .B1(new_n638), .B2(new_n568), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n606), .A2(new_n637), .A3(new_n567), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n567), .A2(new_n603), .A3(new_n605), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n598), .B(new_n631), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n567), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n639), .B1(new_n650), .B2(KEYINPUT101), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n651), .A2(new_n646), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n647), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n642), .B1(new_n651), .B2(new_n637), .ZN(new_n658));
  INV_X1    g457(.A(new_n646), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT103), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n661), .A3(new_n646), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n652), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n655), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n550), .A2(new_n629), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n544), .B(KEYINPUT104), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n462), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n673), .B2(new_n229), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n229), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  MUX2_X1   g476(.A(KEYINPUT42), .B(new_n674), .S(new_n677), .Z(G1325gat));
  NOR2_X1   g477(.A1(new_n479), .A2(new_n494), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n500), .B1(new_n499), .B2(new_n470), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(G15gat), .B1(new_n667), .B2(new_n681), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n679), .A2(new_n680), .B1(new_n505), .B2(new_n506), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n495), .A2(new_n501), .A3(new_n503), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n682), .B1(new_n667), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT106), .ZN(G1326gat));
  INV_X1    g488(.A(new_n523), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n667), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NOR3_X1   g492(.A1(new_n587), .A2(new_n624), .A3(new_n665), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n550), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n208), .A3(new_n669), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(new_n267), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n587), .A2(new_n665), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n545), .A2(new_n548), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  INV_X1    g503(.A(new_n534), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n509), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n543), .A2(new_n544), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n683), .A2(new_n684), .B1(new_n707), .B2(new_n690), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n534), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n703), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n621), .A2(KEYINPUT109), .A3(new_n623), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT109), .B1(new_n621), .B2(new_n623), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n536), .A2(new_n549), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n627), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n701), .B(new_n702), .C1(new_n715), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT110), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n509), .A3(new_n704), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n708), .B2(new_n534), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n549), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n716), .A3(new_n713), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n624), .B1(new_n536), .B2(new_n549), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n701), .A4(new_n702), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n668), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n700), .B1(new_n208), .B2(new_n729), .ZN(G1328gat));
  NAND3_X1  g529(.A1(new_n698), .A2(new_n209), .A3(new_n462), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT46), .Z(new_n732));
  AOI21_X1  g531(.A(new_n543), .B1(new_n720), .B2(new_n728), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n209), .B2(new_n733), .ZN(G1329gat));
  AND3_X1   g533(.A1(new_n696), .A2(new_n681), .A3(new_n697), .ZN(new_n735));
  INV_X1    g534(.A(G43gat), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT47), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n685), .B1(new_n720), .B2(new_n728), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n736), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  OAI21_X1  g539(.A(G43gat), .B1(new_n719), .B2(new_n685), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n735), .A2(new_n736), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n739), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n740), .B1(new_n739), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1330gat));
  OAI21_X1  g546(.A(G50gat), .B1(new_n719), .B2(new_n523), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n698), .A2(new_n335), .A3(new_n690), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT48), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n720), .A2(new_n728), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n690), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G50gat), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n749), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n750), .B1(new_n754), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g554(.A1(new_n267), .A2(new_n723), .A3(new_n629), .A4(new_n665), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n669), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n462), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n756), .A2(new_n763), .A3(new_n681), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n756), .A2(new_n686), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n763), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g566(.A1(new_n756), .A2(new_n690), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n587), .A2(new_n701), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n723), .A2(new_n627), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT51), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n666), .ZN(new_n773));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n669), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n665), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT112), .Z(new_n776));
  AND2_X1   g575(.A1(new_n726), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n668), .A2(new_n589), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n773), .A2(new_n590), .A3(new_n462), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n462), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n771), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT51), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n543), .A2(new_n666), .A3(G92gat), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n781), .A2(G92gat), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n784), .B1(new_n789), .B2(new_n783), .ZN(G1337gat));
  INV_X1    g589(.A(G99gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n791), .A3(new_n681), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n686), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n791), .B2(new_n794), .ZN(G1338gat));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n690), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n523), .A2(G106gat), .A3(new_n666), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n797), .B(new_n798), .C1(new_n772), .C2(new_n800), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n796), .A2(G106gat), .B1(new_n787), .B2(new_n799), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n798), .ZN(G1339gat));
  NAND2_X1  g602(.A1(new_n658), .A2(new_n659), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT54), .B1(new_n660), .B2(new_n662), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n656), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n661), .B1(new_n644), .B2(new_n646), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT103), .B(new_n659), .C1(new_n641), .C2(new_n643), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT114), .B1(new_n812), .B2(new_n655), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n805), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n805), .B(KEYINPUT55), .C1(new_n808), .C2(new_n813), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n657), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n816), .A2(new_n820), .A3(new_n657), .A4(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n701), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n247), .A2(new_n248), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT116), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n252), .B1(new_n251), .B2(new_n239), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n259), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n263), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n665), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n713), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n713), .A2(new_n819), .A3(new_n821), .A4(new_n827), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n586), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n625), .A2(new_n267), .A3(new_n628), .A4(new_n666), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n832), .A2(KEYINPUT117), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT117), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n668), .ZN(new_n836));
  INV_X1    g635(.A(new_n547), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n271), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n701), .A2(new_n346), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(G1340gat));
  NOR2_X1   g640(.A1(new_n838), .A2(new_n666), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(new_n344), .ZN(G1341gat));
  NOR2_X1   g642(.A1(new_n838), .A2(new_n586), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT67), .B(G127gat), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(KEYINPUT118), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(KEYINPUT118), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n844), .B2(new_n847), .ZN(G1342gat));
  NOR3_X1   g647(.A1(new_n838), .A2(G134gat), .A3(new_n624), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n838), .B2(new_n624), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n850), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n832), .A2(new_n833), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n832), .A2(KEYINPUT117), .A3(new_n833), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n690), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n271), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n685), .A2(new_n669), .A3(new_n543), .ZN(new_n862));
  INV_X1    g661(.A(new_n833), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n828), .B1(new_n271), .B2(new_n818), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n624), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n587), .B1(new_n865), .B2(new_n830), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n690), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n860), .A2(new_n861), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT122), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n860), .A2(new_n868), .A3(new_n871), .A4(new_n861), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(G141gat), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n690), .A3(new_n859), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n862), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n272), .A3(new_n861), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT121), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NOR4_X1   g677(.A1(new_n874), .A2(G141gat), .A3(new_n271), .A4(new_n862), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n873), .A2(new_n877), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n860), .A2(new_n701), .A3(new_n868), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(G141gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n883), .B2(G141gat), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(new_n879), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(new_n878), .ZN(G1344gat));
  NAND3_X1  g687(.A1(new_n875), .A2(new_n275), .A3(new_n665), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(new_n862), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n629), .A2(new_n271), .A3(new_n666), .ZN(new_n893));
  INV_X1    g692(.A(new_n827), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n818), .A2(new_n894), .A3(new_n624), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n587), .B1(new_n865), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n858), .B(new_n690), .C1(new_n893), .C2(new_n896), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n891), .A2(new_n665), .A3(new_n892), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n890), .B1(new_n898), .B2(G148gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n860), .A2(new_n868), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n890), .B1(new_n900), .B2(new_n666), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n275), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n889), .B1(new_n899), .B2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(G155gat), .B1(new_n900), .B2(new_n586), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n875), .A2(new_n279), .A3(new_n587), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n900), .B2(new_n714), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n875), .A2(new_n280), .A3(new_n627), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1347gat));
  NAND4_X1  g708(.A1(new_n857), .A2(new_n542), .A3(new_n668), .A4(new_n859), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n543), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n408), .A3(new_n701), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n861), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT123), .B1(new_n913), .B2(G169gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(G1348gat));
  NAND2_X1  g715(.A1(new_n911), .A2(new_n665), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g717(.A(new_n396), .B1(new_n911), .B2(new_n587), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n911), .A2(new_n587), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n920), .B(new_n921), .C1(new_n403), .C2(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n403), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT60), .B1(new_n924), .B2(new_n919), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n399), .A3(new_n713), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n543), .A3(new_n624), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT124), .B1(new_n928), .B2(new_n399), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n834), .A2(new_n835), .A3(new_n669), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n931), .A2(new_n542), .A3(new_n462), .A4(new_n627), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n933), .A3(G190gat), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n929), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n930), .B1(new_n929), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n927), .B1(new_n935), .B2(new_n936), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n686), .A2(new_n523), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n931), .A2(new_n462), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n701), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n891), .A2(new_n897), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n686), .A2(new_n669), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n462), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n891), .A2(KEYINPUT125), .A3(new_n897), .ZN(new_n948));
  AND4_X1   g747(.A1(new_n861), .A2(new_n944), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n941), .B1(new_n949), .B2(new_n940), .ZN(G1352gat));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n931), .A2(new_n951), .A3(new_n462), .A4(new_n938), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(new_n666), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n944), .A2(new_n665), .A3(new_n947), .A4(new_n948), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G204gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  NOR2_X1   g756(.A1(new_n946), .A2(new_n586), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n891), .A2(new_n897), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(new_n295), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n962), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n964), .B(new_n965), .C1(new_n959), .C2(new_n295), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n939), .A2(new_n295), .A3(new_n587), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(G1354gat));
  AOI21_X1  g767(.A(G218gat), .B1(new_n939), .B2(new_n713), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n624), .A2(new_n296), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT127), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n969), .B1(new_n970), .B2(new_n972), .ZN(G1355gat));
endmodule


