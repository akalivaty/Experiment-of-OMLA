//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(G183gat), .B(G211gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT98), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT19), .Z(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G155gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT20), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n204), .B(new_n206), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G71gat), .B(G78gat), .Z(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT97), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n213), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n212), .B(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT97), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT21), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT99), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT93), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G8gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n222), .B(new_n227), .C1(new_n225), .C2(G1gat), .ZN(new_n230));
  OR3_X1    g029(.A1(new_n222), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n229), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n232), .A2(G8gat), .B1(new_n233), .B2(new_n223), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n220), .A2(new_n221), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n218), .A2(KEYINPUT97), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n214), .A2(new_n215), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(G8gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n223), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT99), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G231gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n235), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n235), .B2(new_n243), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n237), .A2(new_n238), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT21), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n243), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n244), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(new_n246), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n208), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n247), .B2(new_n248), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n252), .A3(new_n246), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n207), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT41), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G162gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(G29gat), .A2(G36gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT14), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT14), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(G29gat), .B2(G36gat), .ZN(new_n268));
  OAI211_X1 g067(.A(KEYINPUT89), .B(new_n266), .C1(new_n268), .C2(new_n265), .ZN(new_n269));
  AND2_X1   g068(.A1(G43gat), .A2(G50gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(G43gat), .A2(G50gat), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT15), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n269), .B(new_n272), .Z(new_n273));
  MUX2_X1   g072(.A(new_n268), .B(new_n267), .S(new_n265), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT15), .ZN(new_n275));
  INV_X1    g074(.A(new_n270), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT90), .B(G43gat), .Z(new_n277));
  INV_X1    g076(.A(G50gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT91), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT91), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT17), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(KEYINPUT91), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n273), .A2(new_n280), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT100), .B(KEYINPUT7), .Z(new_n289));
  INV_X1    g088(.A(G85gat), .ZN(new_n290));
  INV_X1    g089(.A(G92gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G99gat), .A2(G106gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n289), .A2(new_n292), .B1(KEYINPUT8), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n291), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n290), .B2(new_n291), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G99gat), .B(G106gat), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n298), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n288), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n281), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n301), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n261), .A2(KEYINPUT41), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G134gat), .ZN(new_n308));
  INV_X1    g107(.A(G134gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n303), .A2(new_n309), .A3(new_n305), .A4(new_n306), .ZN(new_n310));
  XNOR2_X1  g109(.A(G190gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n308), .B2(new_n310), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n264), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n311), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n263), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT102), .ZN(new_n320));
  NAND2_X1  g119(.A1(G230gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n298), .A2(new_n299), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n298), .A2(new_n299), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n214), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(new_n326), .C1(new_n249), .C2(new_n301), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n249), .A2(KEYINPUT10), .A3(new_n301), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n322), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n249), .A2(new_n301), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n321), .B1(new_n330), .B2(new_n325), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n320), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G120gat), .B(G148gat), .ZN(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n335), .B(G204gat), .Z(new_n336));
  XNOR2_X1  g135(.A(new_n332), .B(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n260), .A2(new_n315), .A3(new_n319), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G227gat), .ZN(new_n339));
  INV_X1    g138(.A(G233gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G183gat), .ZN(new_n343));
  INV_X1    g142(.A(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT66), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT65), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n345), .A2(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT64), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT64), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT24), .ZN(new_n354));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT66), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n349), .A2(new_n350), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n361), .A2(new_n362), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT25), .ZN(new_n365));
  AND2_X1   g164(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n344), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT67), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n369), .A2(KEYINPUT67), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT68), .B1(new_n359), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n373), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT68), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n374), .A2(new_n375), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT27), .B(G183gat), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(KEYINPUT67), .A3(new_n369), .A4(new_n344), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n372), .A2(new_n379), .A3(new_n381), .A4(new_n355), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n355), .A2(new_n351), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(new_n347), .A3(new_n345), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n388), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n389));
  INV_X1    g188(.A(G127gat), .ZN(new_n390));
  INV_X1    g189(.A(G120gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G113gat), .ZN(new_n392));
  INV_X1    g191(.A(G113gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G120gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT1), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n309), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(G127gat), .B1(new_n388), .B2(KEYINPUT1), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n396), .A3(new_n390), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(G134gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n383), .B1(new_n358), .B2(new_n363), .ZN(new_n404));
  INV_X1    g203(.A(new_n386), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n399), .A2(new_n400), .A3(G134gat), .ZN(new_n407));
  AOI21_X1  g206(.A(G134gat), .B1(new_n399), .B2(new_n400), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n409), .A3(new_n382), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n342), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G71gat), .ZN(new_n415));
  INV_X1    g214(.A(G99gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n410), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n409), .B1(new_n406), .B2(new_n382), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n341), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT32), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT34), .B1(new_n411), .B2(new_n424), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n419), .A2(new_n420), .A3(new_n341), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n423), .B2(new_n425), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n418), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n423), .A2(new_n425), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n426), .ZN(new_n432));
  INV_X1    g231(.A(new_n418), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(new_n278), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT83), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n439), .B(KEYINPUT31), .Z(new_n440));
  INV_X1    g239(.A(KEYINPUT73), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT72), .B(G211gat), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT22), .B1(new_n442), .B2(G218gat), .ZN(new_n443));
  AND2_X1   g242(.A1(G197gat), .A2(G204gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(G197gat), .A2(G204gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n441), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G211gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT72), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G211gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n451), .A3(G218gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT22), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n446), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G211gat), .B(G218gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n446), .B1(new_n452), .B2(new_n453), .ZN(new_n460));
  INV_X1    g259(.A(new_n457), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT73), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT2), .ZN(new_n467));
  INV_X1    g266(.A(G141gat), .ZN(new_n468));
  INV_X1    g267(.A(G148gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G141gat), .A2(G148gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473));
  XNOR2_X1  g272(.A(G155gat), .B(G162gat), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n465), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G228gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n458), .A2(KEYINPUT74), .A3(new_n462), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT74), .B1(new_n458), .B2(new_n462), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n464), .B1(new_n475), .B2(new_n476), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT80), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT80), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n464), .C1(new_n475), .C2(new_n476), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT29), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n478), .B(new_n480), .C1(new_n483), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n485), .A2(new_n487), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n490), .A2(new_n459), .B1(new_n462), .B2(new_n458), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n473), .ZN(new_n492));
  INV_X1    g291(.A(new_n474), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n463), .B2(new_n464), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n479), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n499));
  INV_X1    g298(.A(G22gat), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n489), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n489), .A2(new_n498), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT84), .B1(new_n502), .B2(G22gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n489), .A2(new_n498), .A3(new_n500), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n440), .B(new_n501), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n500), .B1(new_n489), .B2(new_n498), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n504), .B1(new_n509), .B2(KEYINPUT84), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(KEYINPUT85), .A3(new_n440), .A4(new_n501), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n505), .A2(new_n509), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n440), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n436), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G226gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n340), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n387), .B2(new_n459), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n406), .B2(new_n382), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n483), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n457), .B1(new_n460), .B2(KEYINPUT73), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n443), .A2(new_n441), .A3(new_n446), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n462), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n387), .A2(new_n518), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT29), .B1(new_n406), .B2(new_n382), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n528), .B(new_n529), .C1(new_n530), .C2(new_n518), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533));
  XOR2_X1   g332(.A(G8gat), .B(G36gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G64gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n291), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT75), .ZN(new_n537));
  OR3_X1    g336(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n533), .B1(new_n532), .B2(new_n537), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n522), .B2(new_n531), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n538), .A2(new_n539), .B1(KEYINPUT30), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT78), .ZN(new_n542));
  INV_X1    g341(.A(new_n536), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n525), .B2(new_n526), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n458), .A2(KEYINPUT74), .A3(new_n462), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n382), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n548), .A2(new_n404), .A3(new_n405), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n520), .B1(new_n549), .B2(KEYINPUT29), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n547), .B1(new_n550), .B2(new_n529), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n519), .A2(new_n527), .A3(new_n521), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n543), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT77), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n542), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT78), .B(KEYINPUT30), .C1(new_n554), .C2(new_n556), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n541), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G1gat), .B(G29gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT0), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G57gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n290), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n477), .A2(KEYINPUT3), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n486), .B1(new_n496), .B2(new_n464), .ZN(new_n569));
  INV_X1    g368(.A(new_n487), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n402), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n496), .A2(new_n398), .A3(new_n401), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT4), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT4), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n496), .A2(new_n398), .A3(new_n574), .A4(new_n401), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G225gat), .A2(G233gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT5), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n402), .A2(new_n477), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n577), .B1(new_n581), .B2(new_n572), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n409), .B1(new_n485), .B2(new_n487), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n583), .A2(new_n568), .B1(new_n573), .B2(new_n575), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n582), .B1(new_n584), .B2(new_n577), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n567), .B(new_n580), .C1(new_n585), .C2(new_n579), .ZN(new_n586));
  INV_X1    g385(.A(new_n582), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n579), .B1(new_n578), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT5), .B1(new_n584), .B2(new_n577), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n566), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT87), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n587), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT5), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(new_n567), .A3(new_n580), .A4(new_n591), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n597), .A2(new_n594), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n516), .A2(new_n562), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n586), .A2(new_n590), .A3(KEYINPUT82), .A4(new_n592), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n597), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n555), .B1(new_n532), .B2(new_n543), .ZN(new_n608));
  AOI211_X1 g407(.A(KEYINPUT77), .B(new_n536), .C1(new_n522), .C2(new_n531), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n558), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT78), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n557), .A2(new_n542), .A3(new_n558), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n613), .A3(new_n541), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n514), .B1(new_n508), .B2(new_n511), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n614), .A2(new_n615), .A3(new_n436), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n603), .B1(new_n616), .B2(new_n599), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT71), .B1(new_n430), .B2(new_n435), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n618), .A2(KEYINPUT70), .A3(KEYINPUT36), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n436), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT70), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n436), .B2(KEYINPUT70), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n619), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n581), .A2(new_n577), .A3(new_n572), .ZN(new_n627));
  OAI211_X1 g426(.A(KEYINPUT39), .B(new_n627), .C1(new_n584), .C2(new_n577), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n584), .A2(new_n577), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n566), .B(new_n628), .C1(new_n629), .C2(KEYINPUT39), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n586), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n561), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n598), .A2(new_n600), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n550), .A2(new_n547), .A3(new_n529), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n527), .B1(new_n519), .B2(new_n521), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT37), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n537), .B1(new_n638), .B2(KEYINPUT86), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT38), .B1(new_n532), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n639), .B(new_n641), .C1(KEYINPUT86), .C2(new_n638), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n543), .B1(new_n532), .B2(new_n640), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n640), .B2(new_n532), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT38), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n635), .A2(new_n557), .A3(new_n642), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n512), .A2(new_n515), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n634), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n614), .A2(new_n615), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n626), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n338), .B1(new_n617), .B2(new_n650), .ZN(new_n651));
  AOI211_X1 g450(.A(new_n284), .B(KEYINPUT17), .C1(new_n273), .C2(new_n280), .ZN(new_n652));
  AND4_X1   g451(.A1(new_n273), .A2(new_n280), .A3(new_n285), .A4(new_n286), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n234), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G229gat), .A2(G233gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n234), .A2(new_n281), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n656), .B1(new_n288), .B2(new_n234), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(KEYINPUT18), .A3(new_n655), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT94), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n304), .B2(new_n242), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n234), .A2(new_n281), .A3(KEYINPUT94), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n657), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n655), .B(KEYINPUT13), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n670));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(G169gat), .B(G197gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT12), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n660), .A2(new_n662), .A3(new_n675), .A4(new_n668), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT95), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(KEYINPUT95), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n651), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n607), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  INV_X1    g488(.A(G8gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n686), .B2(new_n561), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n225), .A2(new_n690), .ZN(new_n693));
  NOR4_X1   g492(.A1(new_n685), .A2(new_n562), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT42), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(KEYINPUT42), .B2(new_n694), .ZN(G1325gat));
  NAND2_X1  g495(.A1(new_n623), .A2(new_n625), .ZN(new_n697));
  INV_X1    g496(.A(new_n619), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n686), .A2(G15gat), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n436), .ZN(new_n701));
  AOI21_X1  g500(.A(G15gat), .B1(new_n686), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n685), .A2(new_n647), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NAND3_X1  g505(.A1(new_n649), .A2(new_n697), .A3(new_n698), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n634), .A2(new_n646), .A3(new_n647), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n607), .A2(new_n613), .A3(new_n541), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n599), .B1(new_n516), .B2(new_n709), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n615), .A2(new_n561), .A3(new_n601), .A4(new_n436), .ZN(new_n711));
  OAI22_X1  g510(.A1(new_n707), .A2(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n315), .A2(new_n319), .ZN(new_n713));
  INV_X1    g512(.A(new_n336), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n332), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n260), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n712), .A2(new_n684), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(G29gat), .A3(new_n607), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT45), .Z(new_n719));
  INV_X1    g518(.A(new_n713), .ZN(new_n720));
  AOI211_X1 g519(.A(KEYINPUT44), .B(new_n720), .C1(new_n617), .C2(new_n650), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n712), .B2(new_n713), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n679), .B(new_n716), .C1(new_n721), .C2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724), .B2(new_n607), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(new_n725), .ZN(G1328gat));
  OR3_X1    g525(.A1(new_n717), .A2(G36gat), .A3(new_n562), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n728));
  OAI21_X1  g527(.A(G36gat), .B1(new_n724), .B2(new_n562), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(new_n277), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n724), .B2(new_n626), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n717), .A2(new_n732), .A3(new_n436), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1330gat));
  AOI21_X1  g538(.A(new_n720), .B1(new_n617), .B2(new_n650), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n722), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n647), .A2(new_n278), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n679), .A3(new_n716), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n740), .A2(new_n745), .A3(new_n684), .A4(new_n716), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n615), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n278), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n743), .A2(new_n748), .A3(new_n750), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1331gat));
  INV_X1    g553(.A(new_n260), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n713), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n679), .A2(new_n337), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n712), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT105), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n712), .A2(new_n760), .A3(new_n756), .A4(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n607), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT106), .B(G57gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1332gat));
  OAI22_X1  g564(.A1(new_n762), .A2(new_n562), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT49), .B(G64gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n759), .A2(new_n561), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n762), .B2(new_n626), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n436), .A2(G71gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n761), .A3(new_n775), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n774), .B1(new_n773), .B2(new_n776), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(G1334gat));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n647), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g580(.A1(new_n260), .A2(new_n679), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n712), .A2(new_n713), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n607), .A2(new_n337), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n290), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n741), .A2(new_n782), .A3(new_n788), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n791), .B2(new_n290), .ZN(G1336gat));
  OAI211_X1 g591(.A(new_n715), .B(new_n782), .C1(new_n721), .C2(new_n723), .ZN(new_n793));
  OAI21_X1  g592(.A(G92gat), .B1(new_n793), .B2(new_n562), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n562), .A2(new_n337), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n787), .A2(new_n291), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n291), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n783), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n800), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n741), .A2(new_n561), .A3(new_n715), .A4(new_n782), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(G92gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n798), .B1(new_n805), .B2(new_n795), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n793), .B2(new_n626), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n416), .A3(new_n701), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n337), .B2(new_n808), .ZN(G1338gat));
  NOR2_X1   g608(.A1(new_n647), .A2(new_n337), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n782), .B(new_n810), .C1(new_n721), .C2(new_n723), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(G106gat), .ZN(new_n812));
  INV_X1    g611(.A(G106gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n801), .B2(new_n802), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT53), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n741), .A2(new_n817), .A3(new_n782), .A4(new_n810), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n818), .A2(G106gat), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n822));
  INV_X1    g621(.A(new_n814), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n787), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g623(.A(KEYINPUT110), .B(new_n814), .C1(new_n785), .C2(new_n786), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n816), .B1(new_n820), .B2(new_n826), .ZN(G1339gat));
  NAND2_X1  g626(.A1(new_n654), .A2(new_n657), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(KEYINPUT113), .A3(G229gat), .A4(G233gat), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n661), .B2(new_n655), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n829), .B(new_n831), .C1(new_n667), .C2(new_n666), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n674), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n715), .A2(new_n833), .A3(new_n678), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n329), .A2(new_n331), .A3(new_n336), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n327), .A2(new_n328), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n321), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n327), .A2(new_n322), .A3(new_n328), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n714), .B1(new_n329), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n836), .B1(new_n843), .B2(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n842), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n679), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n715), .A2(new_n833), .A3(new_n849), .A4(new_n678), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n720), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n844), .A2(new_n847), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n833), .A2(new_n678), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n713), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n260), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n338), .A2(new_n857), .A3(new_n679), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n338), .B2(new_n679), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n562), .A2(new_n687), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n516), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT116), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n393), .A3(new_n679), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n862), .A2(KEYINPUT115), .A3(new_n516), .A4(new_n864), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n683), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n872), .ZN(G1340gat));
  NAND3_X1  g672(.A1(new_n866), .A2(new_n391), .A3(new_n715), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n715), .A3(new_n870), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(G120gat), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n875), .B2(G120gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(G1341gat));
  NOR3_X1   g678(.A1(new_n871), .A2(new_n390), .A3(new_n755), .ZN(new_n880));
  INV_X1    g679(.A(new_n865), .ZN(new_n881));
  AOI21_X1  g680(.A(G127gat), .B1(new_n881), .B2(new_n260), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(G1342gat));
  OAI21_X1  g682(.A(G134gat), .B1(new_n871), .B2(new_n720), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n881), .A2(new_n885), .A3(new_n309), .A4(new_n713), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n862), .A2(new_n309), .A3(new_n516), .A4(new_n864), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT118), .B1(new_n888), .B2(new_n720), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n887), .B1(new_n886), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n884), .B1(new_n890), .B2(new_n891), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n699), .A2(new_n863), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n862), .A2(new_n615), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(G141gat), .A3(new_n683), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n845), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n840), .A2(KEYINPUT119), .A3(new_n842), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n846), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n681), .A2(new_n682), .A3(new_n844), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n713), .B1(new_n900), .B2(new_n834), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n853), .A2(new_n713), .A3(new_n854), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n755), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND4_X1   g702(.A1(new_n260), .A2(new_n315), .A3(new_n319), .A4(new_n337), .ZN(new_n904));
  INV_X1    g703(.A(new_n679), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT112), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n858), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n615), .A2(KEYINPUT57), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n615), .B1(new_n856), .B2(new_n861), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n908), .A2(new_n916), .A3(new_n910), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n912), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n679), .A3(new_n893), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n895), .B1(new_n919), .B2(G141gat), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT58), .ZN(new_n921));
  INV_X1    g720(.A(new_n893), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n908), .B2(new_n910), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT120), .B(new_n909), .C1(new_n903), .C2(new_n907), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n925), .B2(new_n915), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n468), .B1(new_n926), .B2(new_n684), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n895), .A2(KEYINPUT58), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n920), .A2(new_n921), .B1(new_n927), .B2(new_n928), .ZN(G1344gat));
  INV_X1    g728(.A(new_n894), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n469), .A3(new_n715), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n918), .A2(new_n715), .A3(new_n893), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(G148gat), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n935));
  XOR2_X1   g734(.A(new_n893), .B(KEYINPUT122), .Z(new_n936));
  NAND2_X1  g735(.A1(new_n913), .A2(KEYINPUT57), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n904), .A2(new_n683), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n903), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n914), .A3(new_n615), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n936), .A2(new_n937), .A3(new_n715), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n935), .B1(new_n941), .B2(G148gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n931), .B1(new_n934), .B2(new_n942), .ZN(G1345gat));
  INV_X1    g742(.A(G155gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n944), .A3(new_n260), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n926), .A2(new_n260), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n944), .ZN(G1346gat));
  AOI21_X1  g746(.A(G162gat), .B1(new_n930), .B2(new_n713), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n713), .A2(G162gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n926), .B2(new_n949), .ZN(G1347gat));
  AND2_X1   g749(.A1(new_n862), .A2(new_n647), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n561), .A2(new_n607), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(new_n436), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n683), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n951), .A2(new_n953), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n905), .A2(G169gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(G1348gat));
  NOR3_X1   g758(.A1(new_n955), .A2(new_n334), .A3(new_n337), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n334), .B1(new_n957), .B2(new_n337), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n963), .B(new_n334), .C1(new_n957), .C2(new_n337), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n960), .B1(new_n962), .B2(new_n964), .ZN(G1349gat));
  NAND3_X1  g764(.A1(new_n951), .A2(new_n260), .A3(new_n954), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G183gat), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n951), .A2(new_n380), .A3(new_n260), .A4(new_n953), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT60), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n967), .B(new_n968), .C1(KEYINPUT125), .C2(new_n970), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1350gat));
  NAND3_X1  g773(.A1(new_n951), .A2(new_n713), .A3(new_n954), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n975), .A2(new_n976), .A3(G190gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n975), .B2(G190gat), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n713), .A2(new_n344), .ZN(new_n979));
  OAI22_X1  g778(.A1(new_n977), .A2(new_n978), .B1(new_n957), .B2(new_n979), .ZN(G1351gat));
  AND2_X1   g779(.A1(new_n937), .A2(new_n940), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n699), .A2(new_n952), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(G197gat), .B1(new_n983), .B2(new_n683), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n862), .A2(new_n615), .A3(new_n982), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n905), .A2(G197gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  NOR4_X1   g786(.A1(new_n699), .A2(G204gat), .A3(new_n562), .A4(new_n337), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n862), .A2(new_n607), .A3(new_n615), .A4(new_n988), .ZN(new_n989));
  XOR2_X1   g788(.A(new_n989), .B(KEYINPUT62), .Z(new_n990));
  NAND3_X1  g789(.A1(new_n981), .A2(new_n715), .A3(new_n982), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(G204gat), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1353gat));
  NAND4_X1  g792(.A1(new_n937), .A2(new_n260), .A3(new_n940), .A4(new_n982), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(G211gat), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT63), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n994), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(KEYINPUT127), .A3(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(new_n985), .ZN(new_n1000));
  INV_X1    g799(.A(new_n442), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1000), .A2(new_n1001), .A3(new_n260), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n1000), .A2(KEYINPUT126), .A3(new_n1001), .A4(new_n260), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n995), .A2(new_n1007), .A3(new_n996), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n999), .A2(new_n1006), .A3(new_n1008), .ZN(G1354gat));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n983), .A2(new_n1010), .A3(new_n720), .ZN(new_n1011));
  AOI21_X1  g810(.A(G218gat), .B1(new_n1000), .B2(new_n713), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1355gat));
endmodule


