//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT88), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT88), .B1(new_n203), .B2(KEYINPUT15), .ZN(new_n209));
  OAI221_X1 g008(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n204), .C2(new_n209), .ZN(new_n210));
  NOR3_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n202), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n209), .A2(new_n204), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n207), .A2(new_n208), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n219), .A2(KEYINPUT89), .A3(new_n214), .A4(new_n206), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n212), .A2(KEYINPUT87), .A3(new_n213), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(new_n207), .B2(new_n208), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n213), .B1(new_n212), .B2(KEYINPUT87), .ZN(new_n224));
  OAI211_X1 g023(.A(KEYINPUT15), .B(new_n203), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(G1gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(G1gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT16), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(new_n233), .C1(G1gat), .C2(new_n231), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(G8gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT94), .B1(new_n226), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n235), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n235), .B(KEYINPUT92), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n225), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT93), .A4(new_n245), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n248), .A2(new_n239), .A3(new_n237), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n241), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n251), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(KEYINPUT95), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n250), .A2(new_n255), .A3(new_n251), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  INV_X1    g056(.A(G197gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT11), .B(G169gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT12), .Z(new_n262));
  AND2_X1   g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n250), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT18), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(new_n253), .A3(new_n241), .ZN(new_n266));
  INV_X1    g065(.A(new_n262), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n254), .A2(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT2), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT75), .ZN(new_n271));
  OR2_X1    g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n269), .ZN(new_n273));
  INV_X1    g072(.A(G148gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G141gat), .ZN(new_n275));
  INV_X1    g074(.A(G141gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G148gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT75), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n269), .A2(new_n279), .A3(KEYINPUT2), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n271), .A2(new_n273), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G141gat), .B(G148gat), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n269), .B(new_n272), .C1(new_n282), .C2(KEYINPUT2), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G120gat), .ZN(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G113gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT1), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G127gat), .ZN(new_n295));
  INV_X1    g094(.A(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G127gat), .A2(G134gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n289), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(G127gat), .A2(G134gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G127gat), .A2(G134gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(KEYINPUT68), .C1(new_n304), .C2(KEYINPUT1), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n290), .B2(G120gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n292), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n309), .A2(new_n291), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n315));
  OAI22_X1  g114(.A1(new_n313), .A2(new_n315), .B1(new_n302), .B2(new_n301), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n307), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(KEYINPUT1), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(new_n297), .B2(new_n298), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n309), .A2(new_n291), .A3(new_n310), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(KEYINPUT71), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n306), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT76), .B1(new_n288), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(new_n322), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n300), .A2(new_n305), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n287), .A4(new_n285), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n281), .A2(new_n283), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n334), .C1(KEYINPUT4), .C2(new_n332), .ZN(new_n335));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OR3_X1    g136(.A1(new_n335), .A2(KEYINPUT5), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n331), .B1(new_n325), .B2(new_n326), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT79), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n320), .A2(KEYINPUT71), .A3(new_n321), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT71), .B1(new_n320), .B2(new_n321), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n284), .B1(new_n345), .B2(new_n306), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n337), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n339), .B1(new_n342), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n333), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n347), .A2(KEYINPUT78), .A3(new_n333), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n337), .B1(new_n324), .B2(new_n329), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n351), .A2(KEYINPUT80), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT80), .B1(new_n351), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n338), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT85), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n358), .A2(new_n359), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n349), .B1(new_n348), .B2(new_n337), .ZN(new_n368));
  AOI211_X1 g167(.A(KEYINPUT79), .B(new_n336), .C1(new_n346), .C2(new_n347), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT5), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n351), .A2(KEYINPUT80), .A3(new_n360), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT85), .A3(new_n338), .ZN(new_n374));
  XNOR2_X1  g173(.A(G57gat), .B(G85gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  NAND3_X1  g178(.A1(new_n365), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT86), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n365), .A2(new_n374), .A3(new_n382), .A4(new_n379), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n379), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n338), .C1(new_n361), .C2(new_n362), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n379), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G226gat), .ZN(new_n396));
  INV_X1    g195(.A(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT24), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(G183gat), .A3(G190gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT24), .ZN(new_n402));
  NOR2_X1   g201(.A1(G183gat), .A2(G190gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT65), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT23), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT65), .B(new_n400), .C1(new_n402), .C2(new_n403), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n407), .A2(KEYINPUT23), .ZN(new_n410));
  NAND2_X1  g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n406), .A2(new_n408), .A3(new_n409), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT25), .ZN(new_n415));
  INV_X1    g214(.A(new_n404), .ZN(new_n416));
  INV_X1    g215(.A(G169gat), .ZN(new_n417));
  INV_X1    g216(.A(G176gat), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n418), .A2(KEYINPUT64), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(KEYINPUT64), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT23), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT25), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n416), .A2(new_n421), .A3(new_n413), .A4(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n411), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT67), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT26), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT67), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n429), .A3(new_n411), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT27), .B(G183gat), .ZN(new_n432));
  INV_X1    g231(.A(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT28), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT66), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(KEYINPUT66), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n432), .A2(new_n438), .A3(new_n433), .A4(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n431), .A2(new_n437), .A3(new_n401), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n415), .A2(new_n423), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT29), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n398), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n398), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n441), .A2(new_n423), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(new_n415), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G197gat), .B(G204gat), .ZN(new_n449));
  INV_X1    g248(.A(G211gat), .ZN(new_n450));
  INV_X1    g249(.A(G218gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n449), .B1(KEYINPUT22), .B2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G211gat), .B(G218gat), .Z(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT74), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n445), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n398), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT29), .B1(new_n446), .B2(new_n415), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(new_n398), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n457), .B1(new_n464), .B2(new_n456), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n395), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n456), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n469), .B(KEYINPUT37), .C1(new_n456), .C2(new_n448), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n458), .B1(new_n444), .B2(new_n447), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT74), .B1(new_n462), .B2(new_n398), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n456), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n463), .A2(new_n455), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n395), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n465), .A2(new_n466), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n468), .B1(new_n478), .B2(new_n467), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n390), .A2(new_n391), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G228gat), .A2(G233gat), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n287), .A2(new_n443), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n455), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n484), .B2(KEYINPUT83), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(G22gat), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT3), .B1(new_n455), .B2(new_n443), .ZN(new_n487));
  OAI22_X1  g286(.A1(new_n487), .A2(new_n331), .B1(new_n455), .B2(new_n483), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n486), .B(new_n488), .Z(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G50gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT84), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(KEYINPUT84), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n335), .A2(new_n337), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(KEYINPUT39), .C1(new_n337), .C2(new_n348), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n498), .B(new_n385), .C1(KEYINPUT39), .C2(new_n497), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT40), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(KEYINPUT40), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n381), .A2(new_n383), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n457), .B(new_n394), .C1(new_n464), .C2(new_n456), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n476), .A3(KEYINPUT30), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n465), .A2(new_n505), .A3(new_n395), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n496), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n481), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n363), .A2(new_n379), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n387), .A3(new_n386), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n510), .B(new_n507), .C1(new_n512), .C2(new_n391), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n385), .B1(new_n373), .B2(new_n338), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n391), .B1(new_n388), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n507), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT82), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n496), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G43gat), .ZN(new_n519));
  INV_X1    g318(.A(G71gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G99gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(G227gat), .A2(G233gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n442), .A2(new_n327), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n446), .A2(new_n323), .A3(new_n415), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n526), .B2(KEYINPUT33), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT32), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n527), .A2(new_n529), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(new_n525), .A3(new_n523), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT34), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n523), .B2(KEYINPUT72), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n534), .B(new_n536), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(new_n531), .B2(new_n532), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n538), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n533), .A2(KEYINPUT73), .A3(new_n537), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n547), .B2(KEYINPUT36), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n509), .A2(new_n518), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n515), .A2(new_n516), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n510), .ZN(new_n552));
  INV_X1    g351(.A(new_n541), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n515), .A2(KEYINPUT82), .A3(new_n516), .ZN(new_n554));
  INV_X1    g353(.A(new_n496), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n557));
  NOR4_X1   g356(.A1(new_n547), .A2(new_n496), .A3(KEYINPUT35), .A4(new_n507), .ZN(new_n558));
  INV_X1    g357(.A(new_n391), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n388), .B1(new_n381), .B2(new_n383), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n268), .B1(new_n550), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566));
  AND2_X1   g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT98), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT97), .ZN(new_n573));
  OAI221_X1 g372(.A(new_n566), .B1(KEYINPUT9), .B2(new_n567), .C1(new_n570), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n572), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n566), .B1(KEYINPUT9), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n574), .A2(KEYINPUT99), .A3(new_n578), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n585));
  INV_X1    g384(.A(G183gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n235), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n588), .B(new_n590), .C1(KEYINPUT21), .C2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(KEYINPUT21), .ZN(new_n593));
  INV_X1    g392(.A(new_n588), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n594), .B2(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G231gat), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n596), .B1(new_n597), .B2(new_n397), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G211gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n592), .A2(G231gat), .A3(G233gat), .A4(new_n595), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(new_n598), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n565), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(new_n564), .A3(new_n603), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(KEYINPUT100), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(KEYINPUT100), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(G85gat), .A3(G92gat), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT8), .A2(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT100), .B(new_n610), .C1(new_n615), .C2(new_n616), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G99gat), .B(G106gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n221), .B2(new_n225), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n243), .A2(new_n245), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n626), .B2(new_n624), .ZN(new_n627));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n629), .B1(new_n627), .B2(new_n630), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n632), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n632), .B2(new_n637), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n563), .A2(new_n609), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n623), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n619), .A2(KEYINPUT102), .A3(new_n621), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n591), .A2(new_n643), .A3(new_n622), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n580), .A2(new_n624), .A3(KEYINPUT101), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT101), .B1(new_n580), .B2(new_n624), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n584), .A2(KEYINPUT10), .A3(new_n623), .A4(new_n622), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662));
  AOI211_X1 g461(.A(new_n662), .B(new_n655), .C1(new_n649), .C2(new_n650), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT103), .B1(new_n651), .B2(new_n652), .ZN(new_n664));
  AOI211_X1 g463(.A(new_n663), .B(new_n664), .C1(new_n655), .C2(new_n654), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n665), .B2(new_n660), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n641), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n515), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(G1gat), .Z(G1324gat));
  INV_X1    g469(.A(KEYINPUT16), .ZN(new_n671));
  INV_X1    g470(.A(G8gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n641), .A2(new_n667), .A3(new_n507), .A4(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G8gat), .B1(new_n668), .B2(new_n516), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n674), .B2(new_n676), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT104), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n677), .A2(new_n682), .A3(new_n678), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1325gat));
  XOR2_X1   g483(.A(new_n548), .B(KEYINPUT105), .Z(new_n685));
  OAI21_X1  g484(.A(G15gat), .B1(new_n668), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n547), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n668), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT106), .Z(G1326gat));
  NOR2_X1   g488(.A1(new_n668), .A2(new_n555), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NAND2_X1  g491(.A1(new_n501), .A2(new_n500), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n384), .A2(new_n507), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n555), .ZN(new_n695));
  INV_X1    g494(.A(new_n480), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n560), .A2(new_n696), .A3(new_n559), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n549), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n518), .A2(KEYINPUT108), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n700), .B(new_n496), .C1(new_n513), .C2(new_n517), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n562), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n640), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n252), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n253), .A2(KEYINPUT95), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n263), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n266), .A2(new_n267), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n609), .A2(new_n666), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n550), .A2(new_n562), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(KEYINPUT44), .A3(new_n704), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n707), .A2(new_n712), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT109), .B1(new_n716), .B2(new_n515), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT44), .B1(new_n703), .B2(new_n704), .ZN(new_n718));
  AOI211_X1 g517(.A(new_n706), .B(new_n640), .C1(new_n550), .C2(new_n562), .ZN(new_n719));
  INV_X1    g518(.A(new_n713), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722));
  INV_X1    g521(.A(new_n515), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(new_n712), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n717), .A2(G29gat), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n720), .B2(new_n640), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n704), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n563), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n207), .A3(new_n723), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(KEYINPUT45), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(KEYINPUT45), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT110), .B1(new_n725), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n724), .A3(G29gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n736), .B(new_n737), .C1(new_n732), .C2(new_n733), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(G1328gat));
  NOR3_X1   g538(.A1(new_n729), .A2(G36gat), .A3(new_n516), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n716), .B2(new_n516), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1329gat));
  OAI21_X1  g542(.A(G43gat), .B1(new_n716), .B2(new_n549), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n729), .A2(G43gat), .A3(new_n547), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n685), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n721), .A2(new_n712), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n750), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g550(.A(G50gat), .B1(new_n716), .B2(new_n555), .ZN(new_n752));
  OR3_X1    g551(.A1(new_n729), .A2(G50gat), .A3(new_n555), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT48), .Z(G1331gat));
  NAND4_X1  g554(.A1(new_n509), .A2(new_n549), .A3(new_n699), .A4(new_n701), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n667), .B1(new_n756), .B2(new_n562), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n606), .A2(new_n608), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n758), .A2(new_n712), .A3(new_n704), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n515), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n571), .ZN(G1332gat));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n516), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  OAI21_X1  g566(.A(new_n520), .B1(new_n760), .B2(new_n547), .ZN(new_n768));
  INV_X1    g567(.A(new_n760), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(G71gat), .A3(new_n748), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n768), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n769), .A2(new_n496), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n609), .A2(new_n712), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n707), .A2(new_n666), .A3(new_n715), .A4(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n779), .A2(new_n615), .A3(new_n515), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n704), .A4(new_n778), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n640), .B1(new_n756), .B2(new_n562), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n778), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n703), .A2(new_n704), .A3(new_n778), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(KEYINPUT113), .A3(new_n788), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n786), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n723), .A3(new_n666), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n780), .B1(new_n794), .B2(new_n615), .ZN(G1336gat));
  NOR2_X1   g594(.A1(new_n516), .A2(G92gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n666), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  INV_X1    g599(.A(new_n779), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n616), .B1(new_n801), .B2(new_n507), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n793), .A2(KEYINPUT114), .A3(new_n666), .A4(new_n796), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n799), .A2(new_n800), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n781), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n666), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(G92gat), .A3(new_n516), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n808), .B2(new_n802), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n809), .ZN(G1337gat));
  OAI21_X1  g609(.A(G99gat), .B1(new_n779), .B2(new_n685), .ZN(new_n811));
  INV_X1    g610(.A(new_n793), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n667), .A2(new_n547), .A3(G99gat), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT115), .Z(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(G1338gat));
  NOR3_X1   g614(.A1(new_n807), .A2(G106gat), .A3(new_n555), .ZN(new_n816));
  INV_X1    g615(.A(G106gat), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n801), .B2(new_n496), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT53), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n812), .A2(G106gat), .A3(new_n667), .A4(new_n555), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(G1339gat));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n664), .B2(new_n663), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n649), .A2(new_n655), .A3(new_n650), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n659), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n659), .A4(new_n826), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n661), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n712), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n261), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n248), .A2(new_n249), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n239), .B1(new_n835), .B2(new_n237), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n238), .A2(new_n240), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n710), .A2(new_n666), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n704), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n710), .A2(new_n838), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n640), .A3(new_n831), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n758), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n609), .A2(new_n667), .A3(new_n268), .A4(new_n640), .ZN(new_n844));
  AOI211_X1 g643(.A(new_n496), .B(new_n547), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n723), .A3(new_n516), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n268), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n541), .B1(new_n843), .B2(new_n844), .ZN(new_n848));
  AND4_X1   g647(.A1(new_n723), .A2(new_n848), .A3(new_n516), .A4(new_n555), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n290), .A3(new_n712), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT116), .ZN(G1340gat));
  OAI21_X1  g651(.A(G120gat), .B1(new_n846), .B2(new_n667), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n292), .A3(new_n666), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1341gat));
  NOR3_X1   g654(.A1(new_n846), .A2(new_n295), .A3(new_n758), .ZN(new_n856));
  AOI21_X1  g655(.A(G127gat), .B1(new_n849), .B2(new_n609), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  NAND3_X1  g657(.A1(new_n849), .A2(new_n296), .A3(new_n704), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT56), .Z(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n846), .B2(new_n640), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  AND3_X1   g661(.A1(new_n710), .A2(new_n666), .A3(new_n838), .ZN(new_n863));
  XOR2_X1   g662(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n864));
  NAND2_X1  g663(.A1(new_n827), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n661), .A3(new_n830), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n711), .B2(new_n710), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n640), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n704), .A2(new_n710), .A3(new_n838), .A4(new_n832), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n609), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR4_X1   g669(.A1(new_n758), .A2(new_n666), .A3(new_n712), .A4(new_n704), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n496), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT57), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n831), .B1(new_n711), .B2(new_n710), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n640), .B1(new_n863), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n609), .B1(new_n876), .B2(new_n869), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n874), .B(new_n496), .C1(new_n877), .C2(new_n871), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n723), .A2(new_n516), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n548), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n873), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G141gat), .B1(new_n881), .B2(new_n268), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n555), .B1(new_n843), .B2(new_n844), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n685), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n879), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n276), .A3(new_n712), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n878), .A2(new_n880), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n839), .B1(new_n268), .B2(new_n866), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n842), .B1(new_n640), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n844), .B1(new_n892), .B2(new_n609), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n874), .B1(new_n893), .B2(new_n496), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n889), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n873), .A2(KEYINPUT118), .A3(new_n878), .A4(new_n880), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n268), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n886), .B1(new_n897), .B2(new_n276), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n898), .A2(KEYINPUT119), .A3(KEYINPUT58), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT119), .B1(new_n898), .B2(KEYINPUT58), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n888), .B1(new_n899), .B2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  INV_X1    g701(.A(new_n866), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n712), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n704), .B1(new_n904), .B2(new_n839), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n758), .B1(new_n905), .B2(new_n842), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n555), .B1(new_n906), .B2(new_n844), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n883), .A2(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n872), .A2(KEYINPUT120), .A3(new_n874), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(KEYINPUT59), .A3(new_n666), .A4(new_n880), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n667), .B1(new_n895), .B2(new_n896), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(KEYINPUT59), .ZN(new_n914));
  AOI21_X1  g713(.A(G148gat), .B1(new_n885), .B2(new_n666), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n914), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n915), .ZN(G1345gat));
  AOI21_X1  g715(.A(G155gat), .B1(new_n885), .B2(new_n609), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n758), .B1(new_n895), .B2(new_n896), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g718(.A(G162gat), .B1(new_n885), .B2(new_n704), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n640), .B1(new_n895), .B2(new_n896), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n723), .A2(new_n516), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n845), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n268), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n848), .A2(new_n555), .A3(new_n923), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n417), .A3(new_n712), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(G1348gat));
  OAI21_X1  g728(.A(new_n418), .B1(new_n926), .B2(new_n667), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT121), .ZN(new_n931));
  NOR4_X1   g730(.A1(new_n924), .A2(new_n667), .A3(new_n419), .A4(new_n420), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n432), .A3(new_n609), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n924), .B2(new_n758), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n845), .A2(KEYINPUT122), .A3(new_n609), .A4(new_n923), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n938), .B2(new_n586), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n924), .B2(new_n640), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n433), .A3(new_n704), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1351gat));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  INV_X1    g744(.A(new_n923), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n884), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n883), .A2(KEYINPUT123), .A3(new_n685), .A4(new_n923), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n258), .A3(new_n712), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n748), .A2(new_n946), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n911), .A2(new_n712), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n258), .B2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n883), .A2(new_n954), .A3(new_n685), .A4(new_n923), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT62), .B1(new_n955), .B2(new_n667), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n955), .A2(KEYINPUT62), .A3(new_n667), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n911), .A2(new_n666), .A3(new_n951), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n956), .B(new_n957), .C1(new_n958), .C2(new_n954), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT124), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n911), .A2(new_n609), .A3(new_n951), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G211gat), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(KEYINPUT126), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n947), .A2(new_n450), .A3(new_n609), .A4(new_n948), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT125), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n962), .A2(new_n969), .A3(new_n963), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n968), .A3(new_n970), .ZN(G1354gat));
  NAND3_X1  g770(.A1(new_n949), .A2(new_n451), .A3(new_n704), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n911), .A2(new_n704), .A3(new_n951), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n451), .B2(new_n973), .ZN(G1355gat));
endmodule


