//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n546, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT64), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n460), .B2(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n459), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G101), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n461), .A2(new_n463), .A3(G137), .A4(new_n459), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT66), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(new_n461), .A2(new_n463), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n461), .A2(new_n463), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(new_n459), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G124), .B1(G136), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n484));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(new_n459), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n459), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT68), .A2(KEYINPUT4), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT68), .A2(KEYINPUT4), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n461), .A2(new_n463), .A3(new_n491), .A4(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n459), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n495), .A2(new_n498), .A3(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT69), .B1(new_n503), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT6), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n504), .A2(new_n507), .B1(new_n503), .B2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n516), .A2(new_n506), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n504), .A2(new_n507), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n503), .A2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(G543), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n515), .A2(new_n517), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n514), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND3_X1  g106(.A1(new_n508), .A2(G90), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n508), .A2(G52), .A3(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n511), .B2(new_n512), .ZN(new_n535));
  AND2_X1   g110(.A1(G77), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(G651), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n514), .A2(G81), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n506), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n521), .A2(G43), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  XOR2_X1   g122(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n548));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(G188));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n520), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n508), .A2(G91), .A3(new_n513), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n511), .B2(new_n512), .ZN(new_n557));
  AND2_X1   g132(.A1(G78), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n508), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n554), .A2(new_n555), .A3(new_n559), .A4(new_n560), .ZN(G299));
  NAND2_X1  g136(.A1(new_n514), .A2(G87), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n521), .A2(G49), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  NAND2_X1  g140(.A1(new_n514), .A2(G86), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n506), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n521), .A2(G48), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(G305));
  NAND2_X1  g145(.A1(new_n514), .A2(G85), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n506), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n521), .A2(G47), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n508), .A2(G92), .A3(new_n513), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT10), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n506), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G54), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n520), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n579), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT72), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n578), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n576), .B1(new_n589), .B2(G868), .ZN(G284));
  OAI21_X1  g165(.A(new_n576), .B1(new_n589), .B2(G868), .ZN(G321));
  NAND2_X1  g166(.A1(G286), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(G299), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(G868), .B2(new_n593), .ZN(G297));
  OAI21_X1  g169(.A(new_n592), .B1(G868), .B2(new_n593), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g176(.A1(new_n468), .A2(new_n469), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n476), .ZN(new_n603));
  XOR2_X1   g178(.A(KEYINPUT73), .B(KEYINPUT12), .Z(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2100), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n481), .A2(G123), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n482), .A2(G135), .ZN(new_n609));
  OR2_X1    g184(.A1(G99), .A2(G2105), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2096), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n607), .A2(new_n613), .ZN(G156));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n616));
  XOR2_X1   g191(.A(G2427), .B(G2430), .Z(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT76), .ZN(new_n620));
  INV_X1    g195(.A(G2438), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n620), .A2(new_n621), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n618), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n620), .A2(new_n621), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n626), .A2(new_n617), .A3(new_n622), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT77), .ZN(new_n629));
  INV_X1    g204(.A(G2451), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n625), .A2(new_n627), .A3(new_n631), .A4(KEYINPUT14), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n630), .B1(new_n629), .B2(new_n632), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n616), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n635), .ZN(new_n637));
  INV_X1    g212(.A(new_n616), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(new_n638), .A3(new_n633), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT75), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2454), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n636), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n636), .B2(new_n639), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n615), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G14), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n645), .B2(new_n647), .ZN(new_n650));
  OAI211_X1 g225(.A(KEYINPUT78), .B(new_n646), .C1(new_n643), .C2(new_n644), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2100), .Z(new_n660));
  AND2_X1   g235(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  AOI21_X1  g237(.A(KEYINPUT18), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n670), .A3(new_n672), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n674), .C2(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(G1986), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT22), .B(G1981), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  AND2_X1   g259(.A1(KEYINPUT79), .A2(G29), .ZN(new_n685));
  NOR2_X1   g260(.A1(KEYINPUT79), .A2(G29), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G35), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G162), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT29), .B(G2090), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(G29), .A2(G32), .ZN(new_n692));
  NAND3_X1  g267(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT26), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n602), .A2(G105), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n694), .B(new_n695), .C1(G141), .C2(new_n482), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n481), .A2(new_n697), .A3(G129), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n481), .B2(G129), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n692), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT27), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT88), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n544), .A2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G16), .B2(G19), .ZN(new_n707));
  INV_X1    g282(.A(G1341), .ZN(new_n708));
  OAI22_X1  g283(.A1(new_n702), .A2(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n691), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n482), .A2(G139), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n712), .B(new_n713), .C1(new_n714), .C2(new_n459), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n701), .A2(G33), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(KEYINPUT84), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(KEYINPUT84), .ZN(new_n720));
  INV_X1    g295(.A(G2072), .ZN(new_n721));
  OR3_X1    g296(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n687), .B1(new_n726), .B2(G34), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT85), .Z(new_n728));
  INV_X1    g303(.A(G34), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(KEYINPUT24), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2084), .C1(new_n474), .C2(new_n701), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n702), .A2(new_n705), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n725), .A2(KEYINPUT89), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n733), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n724), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n740), .A2(KEYINPUT23), .A3(G20), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n742));
  INV_X1    g317(.A(G20), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G16), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n744), .C1(new_n593), .C2(new_n740), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(G1956), .Z(new_n746));
  OAI21_X1  g321(.A(new_n730), .B1(new_n474), .B2(new_n701), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  NAND2_X1  g324(.A1(G171), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G5), .B2(G16), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  AND4_X1   g327(.A1(new_n710), .A2(new_n739), .A3(new_n746), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n740), .A2(G4), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n589), .B2(new_n740), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1348), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n687), .A2(KEYINPUT28), .A3(G26), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n481), .A2(G128), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT81), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT82), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n761), .A2(G104), .A3(G2105), .ZN(new_n762));
  INV_X1    g337(.A(G104), .ZN(new_n763));
  AOI21_X1  g338(.A(KEYINPUT82), .B1(new_n763), .B2(new_n459), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n459), .A2(G116), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n762), .A2(new_n764), .A3(new_n765), .A4(new_n460), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G140), .B2(new_n482), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n481), .A2(KEYINPUT81), .A3(G128), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n760), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n757), .B1(new_n770), .B2(new_n701), .ZN(new_n771));
  AOI21_X1  g346(.A(KEYINPUT28), .B1(new_n687), .B2(G26), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT83), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n707), .A2(new_n708), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n753), .A2(new_n756), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n740), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n740), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G1971), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G1971), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G16), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT33), .B(G1976), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G305), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n740), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G6), .B2(new_n740), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT34), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n792), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n791), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT34), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n796), .A2(new_n797), .A3(new_n782), .A4(new_n787), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n740), .A2(G24), .ZN(new_n799));
  INV_X1    g374(.A(G290), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n740), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT80), .B(G1986), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n687), .A2(G25), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n481), .A2(G119), .B1(G131), .B2(new_n482), .ZN(new_n805));
  OR2_X1    g380(.A1(G95), .A2(G2105), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n806), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n804), .B1(new_n809), .B2(new_n687), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT35), .B(G1991), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n794), .A2(new_n798), .A3(new_n803), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n740), .A2(G21), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G168), .B2(new_n740), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1966), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT31), .B(G11), .Z(new_n820));
  INV_X1    g395(.A(KEYINPUT30), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(G28), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(G28), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n822), .A2(new_n823), .A3(new_n701), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n819), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n825), .B1(new_n749), .B2(new_n751), .C1(new_n826), .C2(new_n687), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT90), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n687), .A2(G27), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G164), .B2(new_n687), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT91), .Z(new_n831));
  INV_X1    g406(.A(G2078), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n777), .A2(new_n816), .A3(new_n828), .A4(new_n834), .ZN(G311));
  INV_X1    g410(.A(new_n777), .ZN(new_n836));
  INV_X1    g411(.A(new_n828), .ZN(new_n837));
  INV_X1    g412(.A(new_n816), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n833), .ZN(G150));
  NAND2_X1  g414(.A1(new_n508), .A2(new_n513), .ZN(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n840), .A2(new_n841), .B1(new_n520), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT92), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(new_n506), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n589), .A2(G559), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT38), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT39), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n540), .A2(new_n542), .A3(KEYINPUT93), .A4(new_n543), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n843), .A2(KEYINPUT92), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n843), .A2(KEYINPUT92), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n854), .B(new_n846), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n844), .A2(new_n860), .A3(new_n846), .A4(new_n854), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n853), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n850), .B1(new_n865), .B2(G860), .ZN(G145));
  NAND2_X1  g441(.A1(new_n499), .A2(new_n500), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G2105), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n496), .A2(new_n497), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n868), .B(new_n494), .C1(new_n869), .C2(G2105), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n769), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n700), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n808), .B(new_n605), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n482), .A2(G142), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT94), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n481), .A2(G130), .ZN(new_n878));
  OR2_X1    g453(.A1(G106), .A2(G2105), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n875), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n474), .B(new_n826), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G162), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n474), .B(new_n612), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n488), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n875), .B(new_n881), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n885), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT96), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n891), .A3(new_n715), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n715), .B1(new_n891), .B2(new_n888), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n874), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n888), .A2(new_n891), .ZN(new_n896));
  INV_X1    g471(.A(new_n715), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n873), .A3(new_n892), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT95), .B(G37), .Z(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(G166), .A2(G288), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n784), .A2(G303), .ZN(new_n904));
  AOI21_X1  g479(.A(G305), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(G305), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n800), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(G290), .B1(new_n909), .B2(new_n905), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT98), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n910), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT97), .B1(new_n914), .B2(KEYINPUT42), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n916));
  AOI211_X1 g491(.A(new_n916), .B(new_n911), .C1(new_n910), .C2(new_n908), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n864), .B(new_n598), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n588), .A2(G299), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n578), .B(new_n593), .C1(new_n586), .C2(new_n587), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT41), .B1(new_n920), .B2(new_n921), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  OAI221_X1 g504(.A(new_n913), .B1(new_n917), .B2(new_n915), .C1(new_n923), .C2(new_n927), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n930), .A3(G868), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT99), .B1(new_n847), .B2(G868), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT99), .A4(G868), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n934), .ZN(G331));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  OR2_X1    g512(.A1(G301), .A2(KEYINPUT100), .ZN(new_n938));
  NAND2_X1  g513(.A1(G301), .A2(KEYINPUT100), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(G168), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(G286), .A3(new_n939), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n862), .A2(new_n863), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n862), .A2(new_n863), .B1(new_n941), .B2(new_n942), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n922), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n864), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n948), .B(new_n943), .C1(new_n924), .C2(new_n925), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n946), .A2(new_n949), .A3(new_n914), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n914), .B1(new_n946), .B2(new_n949), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n937), .B(new_n900), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(new_n949), .ZN(new_n953));
  INV_X1    g528(.A(new_n914), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n946), .A2(new_n949), .A3(new_n914), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n952), .B1(new_n957), .B2(new_n937), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT101), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n962), .A3(new_n959), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n937), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT102), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n900), .B1(new_n950), .B2(new_n951), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n957), .A2(new_n968), .A3(new_n937), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n965), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(new_n963), .A3(new_n970), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G164), .B2(G1384), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT103), .B(G40), .Z(new_n974));
  NOR3_X1   g549(.A1(new_n466), .A2(new_n472), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1996), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT104), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT125), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n983), .B(new_n986), .Z(new_n987));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n769), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n872), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n990), .A2(new_n977), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n989), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n983), .A2(new_n872), .B1(new_n995), .B2(new_n977), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n808), .A2(new_n811), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n700), .A2(new_n977), .A3(G1996), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT105), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n988), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n973), .B(new_n976), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n809), .A2(new_n812), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n977), .B1(new_n1003), .B2(new_n997), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n977), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT48), .ZN(new_n1007));
  AND4_X1   g582(.A1(new_n1004), .A2(new_n996), .A3(new_n999), .A4(new_n1007), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n994), .A2(new_n1002), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(G164), .B2(G1384), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n870), .A2(KEYINPUT50), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n976), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G2090), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT106), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n973), .A2(new_n975), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n1022), .A3(new_n1015), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT107), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT55), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1017), .A2(new_n1029), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1025), .A2(G8), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT108), .B(G8), .Z(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1027), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1014), .A2(new_n748), .ZN(new_n1037));
  INV_X1    g612(.A(G1966), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1019), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1034), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1035), .A2(new_n1036), .A3(G168), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1031), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n870), .A2(new_n1012), .A3(new_n975), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(new_n1033), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n784), .A2(G1976), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n784), .A2(G1976), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT111), .B(G86), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n568), .B(new_n569), .C1(new_n840), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G1981), .ZN(new_n1055));
  INV_X1    g630(.A(G1981), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n566), .A2(new_n568), .A3(new_n1056), .A4(new_n569), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1055), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(KEYINPUT112), .A2(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g638(.A(new_n1055), .B1(KEYINPUT112), .B2(KEYINPUT49), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n1045), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT109), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1052), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1069), .A3(new_n784), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1042), .A2(new_n1068), .B1(new_n1071), .B2(new_n1045), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1040), .A2(G168), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1025), .A2(G8), .A3(new_n1030), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1073), .B(new_n1067), .C1(new_n1074), .C2(new_n1027), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1075), .B2(new_n1036), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G286), .A3(new_n1033), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1040), .A2(KEYINPUT119), .A3(G286), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G286), .A2(new_n1033), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT120), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n748), .A2(new_n1014), .B1(new_n1019), .B2(new_n1038), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1040), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT51), .B1(G286), .B2(new_n1033), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1087), .A2(KEYINPUT51), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT62), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1014), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n973), .A2(new_n832), .A3(new_n1018), .A4(new_n975), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1092), .A2(new_n749), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1087), .A2(KEYINPUT51), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1098), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1091), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n554), .A2(new_n1104), .A3(new_n560), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n593), .ZN(new_n1108));
  NAND3_X1  g683(.A1(G299), .A2(new_n1106), .A3(new_n1105), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n973), .A2(new_n975), .A3(new_n1018), .A4(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT113), .B(G1956), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n1112), .C1(new_n1014), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1014), .A2(G1348), .B1(G2067), .B2(new_n1044), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n589), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1112), .B1(new_n1014), .B2(new_n1113), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1110), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1115), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT58), .B(G1341), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n1044), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n973), .A2(new_n978), .A3(new_n1018), .A4(new_n975), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1044), .A2(KEYINPUT115), .A3(new_n1122), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(KEYINPUT117), .A3(new_n544), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1120), .A2(new_n1133), .A3(new_n1114), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1120), .B2(new_n1114), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1128), .A2(KEYINPUT116), .A3(new_n544), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1137), .A2(KEYINPUT59), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g715(.A(KEYINPUT60), .B1(G2067), .B2(new_n1044), .C1(new_n1014), .C2(G1348), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1141), .A2(KEYINPUT118), .A3(new_n588), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n588), .B1(new_n1141), .B2(KEYINPUT118), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1142), .A2(new_n1143), .B1(KEYINPUT118), .B2(new_n1141), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1116), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1121), .B1(new_n1140), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n472), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n973), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n472), .A2(new_n1150), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G40), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n464), .A2(new_n465), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n459), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1152), .A2(KEYINPUT123), .A3(new_n1154), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n973), .A2(new_n1160), .A3(new_n1151), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(new_n1153), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1018), .A2(KEYINPUT53), .A3(new_n832), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1095), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1149), .B1(new_n1167), .B2(G171), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1095), .A2(G301), .A3(new_n1096), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT124), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1095), .A2(new_n1096), .A3(new_n1171), .A4(G301), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1167), .A2(G171), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1149), .B1(new_n1174), .B2(new_n1097), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1103), .B1(new_n1148), .B2(new_n1177), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1068), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1076), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(G290), .A2(G1986), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n977), .B1(new_n1181), .B2(new_n1005), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n996), .A2(new_n1004), .A3(new_n999), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1009), .B1(new_n1180), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(G319), .ZN(new_n1186));
  OR2_X1    g760(.A1(G227), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1187), .A2(KEYINPUT127), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n652), .A2(new_n958), .A3(new_n1188), .ZN(new_n1189));
  OR2_X1    g763(.A1(new_n1187), .A2(KEYINPUT127), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n901), .A2(new_n683), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1191), .ZN(G308));
  AND3_X1   g766(.A1(new_n901), .A2(new_n683), .A3(new_n1190), .ZN(new_n1193));
  NAND4_X1  g767(.A1(new_n1193), .A2(new_n652), .A3(new_n958), .A4(new_n1188), .ZN(G225));
endmodule


