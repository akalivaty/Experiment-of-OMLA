

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  XOR2_X1 U325 ( .A(n479), .B(KEYINPUT28), .Z(n538) );
  XOR2_X1 U326 ( .A(n421), .B(n420), .Z(n293) );
  XOR2_X1 U327 ( .A(KEYINPUT97), .B(n412), .Z(n294) );
  XNOR2_X1 U328 ( .A(n473), .B(KEYINPUT48), .ZN(n474) );
  XNOR2_X1 U329 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n359) );
  XNOR2_X1 U330 ( .A(n475), .B(n474), .ZN(n486) );
  XNOR2_X1 U331 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X1 U332 ( .A(n476), .B(KEYINPUT122), .ZN(n477) );
  XNOR2_X1 U333 ( .A(n478), .B(n477), .ZN(n575) );
  XOR2_X1 U334 ( .A(n432), .B(n431), .Z(n561) );
  XNOR2_X1 U335 ( .A(n366), .B(n365), .ZN(n532) );
  XNOR2_X1 U336 ( .A(KEYINPUT38), .B(n457), .ZN(n512) );
  XNOR2_X1 U337 ( .A(n483), .B(KEYINPUT58), .ZN(n484) );
  XNOR2_X1 U338 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U339 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XNOR2_X1 U341 ( .A(G1GAT), .B(G8GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n295), .B(KEYINPUT68), .ZN(n439) );
  XOR2_X1 U343 ( .A(G113GAT), .B(G15GAT), .Z(n372) );
  XOR2_X1 U344 ( .A(n439), .B(n372), .Z(n297) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G50GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n302) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n298), .B(KEYINPUT8), .ZN(n420) );
  XOR2_X1 U349 ( .A(n420), .B(KEYINPUT69), .Z(n300) );
  NAND2_X1 U350 ( .A1(G229GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U352 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U353 ( .A(G22GAT), .B(G141GAT), .Z(n304) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G36GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U356 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n306) );
  XNOR2_X1 U357 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n578) );
  XOR2_X1 U361 ( .A(G85GAT), .B(KEYINPUT72), .Z(n417) );
  XOR2_X1 U362 ( .A(G71GAT), .B(G120GAT), .Z(n312) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G176GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n369) );
  INV_X1 U365 ( .A(KEYINPUT70), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n369), .B(n313), .ZN(n314) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  NAND2_X1 U368 ( .A1(n314), .A2(n315), .ZN(n319) );
  INV_X1 U369 ( .A(n314), .ZN(n317) );
  INV_X1 U370 ( .A(n315), .ZN(n316) );
  NAND2_X1 U371 ( .A1(n317), .A2(n316), .ZN(n318) );
  NAND2_X1 U372 ( .A1(n319), .A2(n318), .ZN(n323) );
  XOR2_X1 U373 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n321) );
  XNOR2_X1 U374 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n320) );
  XOR2_X1 U375 ( .A(n321), .B(n320), .Z(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n327) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G78GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n324), .B(G148GAT), .ZN(n394) );
  XNOR2_X1 U379 ( .A(G204GAT), .B(G92GAT), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n325), .B(G64GAT), .ZN(n354) );
  XNOR2_X1 U381 ( .A(n394), .B(n354), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U383 ( .A(n417), .B(n328), .Z(n329) );
  XOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT13), .Z(n435) );
  XNOR2_X1 U385 ( .A(n329), .B(n435), .ZN(n466) );
  NOR2_X1 U386 ( .A1(n578), .A2(n466), .ZN(n499) );
  XOR2_X1 U387 ( .A(KEYINPUT101), .B(KEYINPUT37), .Z(n455) );
  XOR2_X1 U388 ( .A(G85GAT), .B(G162GAT), .Z(n331) );
  XNOR2_X1 U389 ( .A(G113GAT), .B(G120GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U391 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n333) );
  XNOR2_X1 U392 ( .A(G148GAT), .B(G155GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U394 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U395 ( .A(KEYINPUT92), .B(G57GAT), .Z(n337) );
  NAND2_X1 U396 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U398 ( .A(KEYINPUT6), .B(n338), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n349) );
  XOR2_X1 U400 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n342) );
  XNOR2_X1 U401 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n347) );
  XNOR2_X1 U403 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n343), .B(KEYINPUT2), .ZN(n392) );
  XOR2_X1 U405 ( .A(KEYINPUT0), .B(G127GAT), .Z(n376) );
  XOR2_X1 U406 ( .A(n392), .B(n376), .Z(n345) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(G134GAT), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U409 ( .A(n347), .B(n346), .Z(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n530) );
  XOR2_X1 U411 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n351) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U414 ( .A(G190GAT), .B(KEYINPUT19), .Z(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n383) );
  INV_X1 U416 ( .A(n383), .ZN(n358) );
  XOR2_X1 U417 ( .A(KEYINPUT94), .B(n354), .Z(n356) );
  NAND2_X1 U418 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n366) );
  XOR2_X1 U421 ( .A(G36GAT), .B(KEYINPUT74), .Z(n416) );
  XNOR2_X1 U422 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n360) );
  XOR2_X1 U423 ( .A(G197GAT), .B(G218GAT), .Z(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n395) );
  XNOR2_X1 U425 ( .A(n416), .B(n395), .ZN(n364) );
  XOR2_X1 U426 ( .A(G8GAT), .B(G176GAT), .Z(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U428 ( .A(KEYINPUT85), .B(KEYINPUT80), .Z(n368) );
  XNOR2_X1 U429 ( .A(KEYINPUT81), .B(KEYINPUT83), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n381) );
  XOR2_X1 U431 ( .A(G43GAT), .B(G134GAT), .Z(n421) );
  XNOR2_X1 U432 ( .A(n421), .B(n369), .ZN(n371) );
  AND2_X1 U433 ( .A1(G227GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n379) );
  XOR2_X1 U436 ( .A(KEYINPUT65), .B(KEYINPUT84), .Z(n375) );
  XNOR2_X1 U437 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U439 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U441 ( .A(n381), .B(n380), .Z(n382) );
  XNOR2_X2 U442 ( .A(n383), .B(n382), .ZN(n535) );
  NAND2_X1 U443 ( .A1(n532), .A2(n535), .ZN(n398) );
  XOR2_X1 U444 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n385) );
  XNOR2_X1 U445 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U447 ( .A(KEYINPUT24), .B(G204GAT), .Z(n387) );
  XOR2_X1 U448 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U449 ( .A(G22GAT), .B(G155GAT), .Z(n440) );
  XNOR2_X1 U450 ( .A(n428), .B(n440), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U452 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U453 ( .A1(G228GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n393) );
  XOR2_X1 U455 ( .A(n393), .B(n392), .Z(n397) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n479) );
  NAND2_X1 U458 ( .A1(n398), .A2(n479), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n399), .B(KEYINPUT98), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n400), .B(KEYINPUT25), .ZN(n404) );
  NOR2_X1 U461 ( .A1(n535), .A2(n479), .ZN(n401) );
  XNOR2_X1 U462 ( .A(KEYINPUT26), .B(n401), .ZN(n576) );
  XNOR2_X1 U463 ( .A(n532), .B(KEYINPUT95), .ZN(n402) );
  XOR2_X1 U464 ( .A(n402), .B(KEYINPUT27), .Z(n407) );
  AND2_X1 U465 ( .A1(n576), .A2(n407), .ZN(n403) );
  OR2_X1 U466 ( .A1(n404), .A2(n403), .ZN(n405) );
  XNOR2_X1 U467 ( .A(KEYINPUT99), .B(n405), .ZN(n406) );
  NOR2_X1 U468 ( .A1(n530), .A2(n406), .ZN(n413) );
  INV_X1 U469 ( .A(KEYINPUT96), .ZN(n409) );
  NAND2_X1 U470 ( .A1(n530), .A2(n407), .ZN(n487) );
  NOR2_X1 U471 ( .A1(n538), .A2(n487), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n535), .B(KEYINPUT86), .ZN(n410) );
  NOR2_X1 U474 ( .A1(n411), .A2(n410), .ZN(n412) );
  NOR2_X1 U475 ( .A1(n413), .A2(n294), .ZN(n498) );
  XOR2_X1 U476 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n415) );
  XNOR2_X1 U477 ( .A(G190GAT), .B(G99GAT), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n432) );
  XOR2_X1 U479 ( .A(n417), .B(n416), .Z(n419) );
  XNOR2_X1 U480 ( .A(G218GAT), .B(G106GAT), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n424) );
  NAND2_X1 U482 ( .A1(G232GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n293), .B(n422), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U485 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n426) );
  XNOR2_X1 U486 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U488 ( .A(n428), .B(n427), .Z(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n561), .B(KEYINPUT36), .ZN(n590) );
  NOR2_X1 U491 ( .A1(n498), .A2(n590), .ZN(n453) );
  XOR2_X1 U492 ( .A(G78GAT), .B(G211GAT), .Z(n434) );
  XNOR2_X1 U493 ( .A(G71GAT), .B(G127GAT), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U495 ( .A(n436), .B(n435), .Z(n438) );
  XNOR2_X1 U496 ( .A(G15GAT), .B(G183GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U498 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U499 ( .A1(G231GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U501 ( .A(n444), .B(n443), .Z(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n446) );
  XNOR2_X1 U503 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U505 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n448) );
  XNOR2_X1 U506 ( .A(KEYINPUT15), .B(KEYINPUT75), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n586) );
  NAND2_X1 U510 ( .A1(n453), .A2(n586), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n529) );
  NAND2_X1 U512 ( .A1(n499), .A2(n529), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT102), .B(n456), .Z(n457) );
  NAND2_X1 U514 ( .A1(n512), .A2(n535), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n459) );
  INV_X1 U516 ( .A(G43GAT), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n586), .A2(n590), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT45), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n463), .A2(n578), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n466), .A2(n464), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT113), .B(n465), .Z(n472) );
  NAND2_X1 U522 ( .A1(n561), .A2(n586), .ZN(n469) );
  XNOR2_X1 U523 ( .A(KEYINPUT41), .B(n466), .ZN(n565) );
  NOR2_X1 U524 ( .A1(n578), .A2(n565), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT46), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT47), .B(n470), .Z(n471) );
  NOR2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n475) );
  XOR2_X1 U529 ( .A(KEYINPUT64), .B(KEYINPUT114), .Z(n473) );
  NAND2_X1 U530 ( .A1(n486), .A2(n532), .ZN(n478) );
  INV_X1 U531 ( .A(KEYINPUT54), .ZN(n476) );
  INV_X1 U532 ( .A(n530), .ZN(n574) );
  AND2_X1 U533 ( .A1(n574), .A2(n479), .ZN(n480) );
  NAND2_X1 U534 ( .A1(n575), .A2(n480), .ZN(n481) );
  XNOR2_X1 U535 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  NAND2_X1 U536 ( .A1(n482), .A2(n535), .ZN(n571) );
  NOR2_X1 U537 ( .A1(n561), .A2(n571), .ZN(n485) );
  INV_X1 U538 ( .A(G190GAT), .ZN(n483) );
  INV_X1 U539 ( .A(n486), .ZN(n488) );
  NOR2_X1 U540 ( .A1(n488), .A2(n487), .ZN(n489) );
  XOR2_X1 U541 ( .A(KEYINPUT115), .B(n489), .Z(n552) );
  INV_X1 U542 ( .A(n552), .ZN(n490) );
  NOR2_X1 U543 ( .A1(n538), .A2(n490), .ZN(n491) );
  NAND2_X1 U544 ( .A1(n535), .A2(n491), .ZN(n548) );
  NOR2_X1 U545 ( .A1(n548), .A2(n578), .ZN(n492) );
  XNOR2_X1 U546 ( .A(KEYINPUT116), .B(n492), .ZN(n493) );
  XOR2_X1 U547 ( .A(G113GAT), .B(n493), .Z(G1340GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n496) );
  INV_X1 U549 ( .A(n586), .ZN(n494) );
  NAND2_X1 U550 ( .A1(n561), .A2(n494), .ZN(n495) );
  XNOR2_X1 U551 ( .A(n496), .B(n495), .ZN(n497) );
  NOR2_X1 U552 ( .A1(n498), .A2(n497), .ZN(n515) );
  AND2_X1 U553 ( .A1(n499), .A2(n515), .ZN(n506) );
  NAND2_X1 U554 ( .A1(n506), .A2(n530), .ZN(n500) );
  XNOR2_X1 U555 ( .A(KEYINPUT34), .B(n500), .ZN(n501) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U557 ( .A1(n506), .A2(n532), .ZN(n502) );
  XNOR2_X1 U558 ( .A(n502), .B(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U559 ( .A(G8GAT), .B(n503), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U561 ( .A1(n506), .A2(n535), .ZN(n504) );
  XNOR2_X1 U562 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n506), .A2(n538), .ZN(n507) );
  XNOR2_X1 U564 ( .A(n507), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .Z(n509) );
  NAND2_X1 U566 ( .A1(n512), .A2(n530), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  XOR2_X1 U568 ( .A(G36GAT), .B(KEYINPUT103), .Z(n511) );
  NAND2_X1 U569 ( .A1(n512), .A2(n532), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n511), .B(n510), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n512), .A2(n538), .ZN(n513) );
  XNOR2_X1 U572 ( .A(n513), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n517) );
  INV_X1 U574 ( .A(n578), .ZN(n514) );
  NOR2_X1 U575 ( .A1(n565), .A2(n514), .ZN(n528) );
  AND2_X1 U576 ( .A1(n528), .A2(n515), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n523), .A2(n530), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U581 ( .A1(n523), .A2(n532), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U583 ( .A(G64GAT), .B(n521), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n523), .A2(n535), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U587 ( .A1(n523), .A2(n538), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n527) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT108), .Z(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  AND2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n530), .A2(n539), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n539), .A2(n532), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n533), .B(KEYINPUT110), .ZN(n534) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  XOR2_X1 U597 ( .A(G99GAT), .B(KEYINPUT111), .Z(n537) );
  NAND2_X1 U598 ( .A1(n539), .A2(n535), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(G1338GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n541) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U603 ( .A(G106GAT), .B(n542), .Z(G1339GAT) );
  NOR2_X1 U604 ( .A1(n565), .A2(n548), .ZN(n544) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n548), .A2(n586), .ZN(n546) );
  XNOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  NOR2_X1 U611 ( .A1(n548), .A2(n561), .ZN(n550) );
  XNOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n576), .A2(n552), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n578), .A2(n560), .ZN(n554) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n558) );
  NOR2_X1 U622 ( .A1(n565), .A2(n560), .ZN(n557) );
  XOR2_X1 U623 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NOR2_X1 U624 ( .A1(n586), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n578), .A2(n571), .ZN(n564) );
  XOR2_X1 U630 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n571), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n567) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT56), .B(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NOR2_X1 U637 ( .A1(n586), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  AND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n589) );
  NOR2_X1 U642 ( .A1(n578), .A2(n589), .ZN(n582) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT126), .B(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U648 ( .A(n589), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n583), .A2(n466), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n589), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

