

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780;

  XNOR2_X1 U373 ( .A(G107), .B(G116), .ZN(n457) );
  XNOR2_X1 U374 ( .A(G122), .B(G140), .ZN(n464) );
  XNOR2_X2 U375 ( .A(n395), .B(n765), .ZN(n659) );
  XNOR2_X2 U376 ( .A(n435), .B(G902), .ZN(n632) );
  XNOR2_X2 U377 ( .A(n436), .B(KEYINPUT92), .ZN(n437) );
  NOR2_X2 U378 ( .A1(n393), .A2(G952), .ZN(n732) );
  XNOR2_X2 U379 ( .A(n488), .B(n487), .ZN(n764) );
  XNOR2_X2 U380 ( .A(n452), .B(n451), .ZN(n488) );
  XNOR2_X2 U381 ( .A(n489), .B(G469), .ZN(n593) );
  NAND2_X2 U382 ( .A1(n578), .A2(n670), .ZN(n441) );
  XNOR2_X2 U383 ( .A(n438), .B(n437), .ZN(n578) );
  NAND2_X1 U384 ( .A1(G234), .A2(G237), .ZN(n443) );
  XNOR2_X1 U385 ( .A(KEYINPUT5), .B(G137), .ZN(n492) );
  XNOR2_X1 U386 ( .A(G122), .B(KEYINPUT7), .ZN(n454) );
  OR2_X1 U387 ( .A1(G902), .A2(G237), .ZN(n371) );
  XNOR2_X1 U388 ( .A(KEYINPUT16), .B(G122), .ZN(n432) );
  INV_X1 U389 ( .A(G134), .ZN(n451) );
  INV_X1 U390 ( .A(G902), .ZN(n514) );
  INV_X2 U391 ( .A(G953), .ZN(n393) );
  AND2_X1 U392 ( .A1(n410), .A2(n671), .ZN(n350) );
  XNOR2_X1 U393 ( .A(n530), .B(n529), .ZN(n563) );
  NAND2_X2 U394 ( .A1(n642), .A2(n641), .ZN(n381) );
  NOR2_X2 U395 ( .A1(n550), .A2(n483), .ZN(n484) );
  XNOR2_X2 U396 ( .A(n600), .B(n442), .ZN(n595) );
  NOR2_X2 U397 ( .A1(G953), .A2(G237), .ZN(n491) );
  AND2_X1 U398 ( .A1(n768), .A2(n636), .ZN(n635) );
  XNOR2_X1 U399 ( .A(n528), .B(n527), .ZN(n657) );
  XNOR2_X1 U400 ( .A(n537), .B(n536), .ZN(n652) );
  OR2_X1 U401 ( .A1(n364), .A2(n538), .ZN(n736) );
  INV_X1 U402 ( .A(KEYINPUT38), .ZN(n361) );
  XOR2_X1 U403 ( .A(G137), .B(G140), .Z(n511) );
  NAND2_X1 U404 ( .A1(n353), .A2(n351), .ZN(n392) );
  NAND2_X1 U405 ( .A1(n352), .A2(KEYINPUT116), .ZN(n351) );
  AND2_X1 U406 ( .A1(n357), .A2(n354), .ZN(n353) );
  NOR2_X1 U407 ( .A1(n665), .A2(n664), .ZN(n669) );
  AND2_X1 U408 ( .A1(n355), .A2(n393), .ZN(n354) );
  NAND2_X1 U409 ( .A1(n356), .A2(KEYINPUT116), .ZN(n355) );
  INV_X1 U410 ( .A(n704), .ZN(n356) );
  NAND2_X1 U411 ( .A1(n705), .A2(n657), .ZN(n530) );
  XNOR2_X1 U412 ( .A(n360), .B(KEYINPUT42), .ZN(n778) );
  AND2_X1 U413 ( .A1(n403), .A2(n350), .ZN(n615) );
  XNOR2_X1 U414 ( .A(n613), .B(n361), .ZN(n671) );
  XNOR2_X1 U415 ( .A(n728), .B(n729), .ZN(n730) );
  NOR2_X1 U416 ( .A1(G902), .A2(n644), .ZN(n461) );
  XNOR2_X1 U417 ( .A(n460), .B(n459), .ZN(n644) );
  NOR2_X1 U418 ( .A1(n447), .A2(n576), .ZN(n448) );
  XNOR2_X1 U419 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U420 ( .A(n764), .B(G146), .ZN(n500) );
  XOR2_X2 U421 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n444) );
  XNOR2_X2 U422 ( .A(KEYINPUT18), .B(KEYINPUT91), .ZN(n423) );
  XNOR2_X2 U423 ( .A(G143), .B(G128), .ZN(n365) );
  XNOR2_X2 U424 ( .A(KEYINPUT66), .B(G101), .ZN(n494) );
  XNOR2_X1 U425 ( .A(KEYINPUT90), .B(KEYINPUT15), .ZN(n435) );
  XNOR2_X1 U426 ( .A(KEYINPUT23), .B(KEYINPUT96), .ZN(n505) );
  NAND2_X1 U427 ( .A1(n359), .A2(n358), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n413), .B(n412), .ZN(n359) );
  INV_X1 U429 ( .A(n359), .ZN(n352) );
  AND2_X1 U430 ( .A1(n704), .A2(n394), .ZN(n358) );
  NOR2_X1 U431 ( .A1(n622), .A2(n621), .ZN(n402) );
  NOR2_X1 U432 ( .A1(n700), .A2(n618), .ZN(n360) );
  NOR2_X1 U433 ( .A1(n676), .A2(n673), .ZN(n617) );
  XNOR2_X1 U434 ( .A(n381), .B(KEYINPUT64), .ZN(n362) );
  OR2_X2 U435 ( .A1(n364), .A2(n690), .ZN(n537) );
  BUF_X1 U436 ( .A(n699), .Z(n363) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n364) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n550) );
  XNOR2_X2 U439 ( .A(n441), .B(n440), .ZN(n600) );
  XNOR2_X1 U440 ( .A(n549), .B(n548), .ZN(n699) );
  NAND2_X1 U441 ( .A1(n425), .A2(n424), .ZN(n368) );
  NAND2_X1 U442 ( .A1(n366), .A2(n367), .ZN(n369) );
  NAND2_X1 U443 ( .A1(n369), .A2(n368), .ZN(n428) );
  INV_X1 U444 ( .A(n425), .ZN(n366) );
  INV_X1 U445 ( .A(n424), .ZN(n367) );
  XNOR2_X1 U446 ( .A(KEYINPUT4), .B(G131), .ZN(n487) );
  INV_X1 U447 ( .A(n651), .ZN(n400) );
  XNOR2_X1 U448 ( .A(G113), .B(KEYINPUT68), .ZN(n430) );
  NAND2_X1 U449 ( .A1(n587), .A2(KEYINPUT73), .ZN(n408) );
  XOR2_X1 U450 ( .A(G478), .B(n461), .Z(n553) );
  XNOR2_X1 U451 ( .A(G104), .B(G110), .ZN(n426) );
  XNOR2_X1 U452 ( .A(n511), .B(n390), .ZN(n389) );
  INV_X1 U453 ( .A(KEYINPUT94), .ZN(n390) );
  XOR2_X1 U454 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n477) );
  NAND2_X1 U455 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U456 ( .A(KEYINPUT84), .ZN(n398) );
  XOR2_X1 U457 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n465) );
  XNOR2_X1 U458 ( .A(G104), .B(G113), .ZN(n462) );
  XOR2_X1 U459 ( .A(G131), .B(G143), .Z(n463) );
  XNOR2_X1 U460 ( .A(n411), .B(n370), .ZN(n410) );
  NAND2_X1 U461 ( .A1(n407), .A2(n404), .ZN(n403) );
  NAND2_X1 U462 ( .A1(n406), .A2(n405), .ZN(n404) );
  AND2_X1 U463 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X1 U464 ( .A(KEYINPUT0), .ZN(n378) );
  XNOR2_X1 U465 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U466 ( .A(n500), .B(n387), .ZN(n722) );
  XNOR2_X1 U467 ( .A(n486), .B(n388), .ZN(n387) );
  XNOR2_X1 U468 ( .A(n389), .B(n485), .ZN(n388) );
  INV_X1 U469 ( .A(KEYINPUT53), .ZN(n391) );
  INV_X1 U470 ( .A(G953), .ZN(n449) );
  XNOR2_X1 U471 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n370) );
  AND2_X1 U472 ( .A1(n559), .A2(KEYINPUT86), .ZN(n372) );
  AND2_X1 U473 ( .A1(n768), .A2(n667), .ZN(n373) );
  NOR2_X1 U474 ( .A1(n591), .A2(n683), .ZN(n374) );
  XNOR2_X1 U475 ( .A(n381), .B(KEYINPUT64), .ZN(n643) );
  BUF_X1 U476 ( .A(n726), .Z(n375) );
  AND2_X2 U477 ( .A1(n362), .A2(n414), .ZN(n376) );
  AND2_X2 U478 ( .A1(n643), .A2(n414), .ZN(n726) );
  XNOR2_X1 U479 ( .A(n399), .B(n398), .ZN(n630) );
  BUF_X1 U480 ( .A(n593), .Z(n377) );
  NOR2_X2 U481 ( .A1(n595), .A2(n448), .ZN(n379) );
  BUF_X1 U482 ( .A(n657), .Z(n380) );
  NAND2_X1 U483 ( .A1(n417), .A2(n373), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n382), .B(KEYINPUT85), .ZN(n570) );
  NAND2_X1 U485 ( .A1(n561), .A2(n562), .ZN(n382) );
  NAND2_X1 U486 ( .A1(n666), .A2(KEYINPUT80), .ZN(n418) );
  NAND2_X1 U487 ( .A1(n668), .A2(n768), .ZN(n665) );
  NAND2_X1 U488 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U489 ( .A1(n726), .A2(G478), .ZN(n645) );
  NAND2_X1 U490 ( .A1(n384), .A2(n383), .ZN(n561) );
  NAND2_X1 U491 ( .A1(n386), .A2(n372), .ZN(n383) );
  NAND2_X1 U492 ( .A1(n385), .A2(n560), .ZN(n384) );
  NAND2_X1 U493 ( .A1(n386), .A2(n559), .ZN(n385) );
  XNOR2_X1 U494 ( .A(n543), .B(KEYINPUT103), .ZN(n386) );
  XNOR2_X2 U495 ( .A(n756), .B(n494), .ZN(n486) );
  XNOR2_X2 U496 ( .A(n427), .B(G107), .ZN(n756) );
  XNOR2_X1 U497 ( .A(n392), .B(n391), .ZN(G75) );
  INV_X1 U498 ( .A(KEYINPUT116), .ZN(n394) );
  XNOR2_X1 U499 ( .A(n396), .B(n510), .ZN(n395) );
  XNOR2_X1 U500 ( .A(n397), .B(n509), .ZN(n396) );
  INV_X1 U501 ( .A(n508), .ZN(n397) );
  NAND2_X1 U502 ( .A1(n401), .A2(n400), .ZN(n399) );
  XNOR2_X1 U503 ( .A(n402), .B(KEYINPUT48), .ZN(n401) );
  NAND2_X1 U504 ( .A1(n591), .A2(n670), .ZN(n411) );
  NAND2_X1 U505 ( .A1(n403), .A2(n410), .ZN(n614) );
  NOR2_X1 U506 ( .A1(n587), .A2(KEYINPUT73), .ZN(n405) );
  INV_X1 U507 ( .A(n577), .ZN(n406) );
  NAND2_X1 U508 ( .A1(n577), .A2(KEYINPUT73), .ZN(n409) );
  INV_X1 U509 ( .A(KEYINPUT81), .ZN(n412) );
  INV_X1 U510 ( .A(n669), .ZN(n414) );
  NAND2_X1 U511 ( .A1(n418), .A2(n416), .ZN(n415) );
  INV_X1 U512 ( .A(n751), .ZN(n417) );
  XNOR2_X1 U513 ( .A(n615), .B(KEYINPUT39), .ZN(n627) );
  XNOR2_X1 U514 ( .A(n531), .B(n490), .ZN(n519) );
  NOR2_X2 U515 ( .A1(n589), .A2(n534), .ZN(n681) );
  INV_X1 U516 ( .A(KEYINPUT46), .ZN(n619) );
  NAND2_X1 U517 ( .A1(n656), .A2(KEYINPUT44), .ZN(n559) );
  INV_X1 U518 ( .A(KEYINPUT88), .ZN(n440) );
  BUF_X1 U519 ( .A(n668), .Z(n751) );
  INV_X1 U520 ( .A(KEYINPUT104), .ZN(n490) );
  BUF_X1 U521 ( .A(n652), .Z(n654) );
  INV_X1 U522 ( .A(KEYINPUT119), .ZN(n647) );
  NAND2_X1 U523 ( .A1(n519), .A2(n374), .ZN(n705) );
  XNOR2_X2 U524 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n420) );
  NAND2_X1 U525 ( .A1(n449), .A2(G224), .ZN(n419) );
  XNOR2_X1 U526 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U527 ( .A(G146), .B(G125), .ZN(n468) );
  INV_X1 U528 ( .A(n468), .ZN(n421) );
  XNOR2_X1 U529 ( .A(n422), .B(n421), .ZN(n425) );
  XNOR2_X2 U530 ( .A(G143), .B(G128), .ZN(n452) );
  XNOR2_X1 U531 ( .A(n365), .B(n423), .ZN(n424) );
  INV_X1 U532 ( .A(n426), .ZN(n427) );
  XNOR2_X1 U533 ( .A(n428), .B(n486), .ZN(n434) );
  XNOR2_X1 U534 ( .A(G119), .B(G116), .ZN(n429) );
  XNOR2_X1 U535 ( .A(n429), .B(KEYINPUT3), .ZN(n431) );
  XNOR2_X1 U536 ( .A(n431), .B(n430), .ZN(n498) );
  XNOR2_X1 U537 ( .A(n432), .B(KEYINPUT70), .ZN(n433) );
  XNOR2_X1 U538 ( .A(n498), .B(n433), .ZN(n757) );
  XNOR2_X1 U539 ( .A(n434), .B(n757), .ZN(n727) );
  NAND2_X1 U540 ( .A1(n727), .A2(n632), .ZN(n438) );
  XNOR2_X1 U541 ( .A(KEYINPUT72), .B(n371), .ZN(n439) );
  AND2_X1 U542 ( .A1(n439), .A2(G210), .ZN(n436) );
  NAND2_X1 U543 ( .A1(n439), .A2(G214), .ZN(n670) );
  XNOR2_X1 U544 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n444), .B(n443), .ZN(n446) );
  NAND2_X1 U546 ( .A1(n446), .A2(G902), .ZN(n445) );
  XNOR2_X1 U547 ( .A(n445), .B(KEYINPUT93), .ZN(n572) );
  NOR2_X1 U548 ( .A1(G898), .A2(n393), .ZN(n761) );
  AND2_X1 U549 ( .A1(n572), .A2(n761), .ZN(n447) );
  NAND2_X1 U550 ( .A1(n446), .A2(G952), .ZN(n698) );
  NOR2_X1 U551 ( .A1(n698), .A2(G953), .ZN(n576) );
  NAND2_X1 U552 ( .A1(G234), .A2(n393), .ZN(n450) );
  XOR2_X1 U553 ( .A(KEYINPUT8), .B(n450), .Z(n502) );
  NAND2_X1 U554 ( .A1(n502), .A2(G217), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n488), .B(n453), .ZN(n460) );
  XOR2_X1 U556 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n455) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U558 ( .A(n456), .B(KEYINPUT100), .Z(n458) );
  XNOR2_X1 U559 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U560 ( .A(n463), .B(n462), .ZN(n467) );
  XNOR2_X1 U561 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U562 ( .A(n467), .B(n466), .Z(n471) );
  XNOR2_X1 U563 ( .A(n468), .B(KEYINPUT10), .ZN(n513) );
  NAND2_X1 U564 ( .A1(n491), .A2(G214), .ZN(n469) );
  XNOR2_X1 U565 ( .A(n513), .B(n469), .ZN(n470) );
  XNOR2_X1 U566 ( .A(n471), .B(n470), .ZN(n714) );
  NOR2_X1 U567 ( .A1(G902), .A2(n714), .ZN(n473) );
  XNOR2_X1 U568 ( .A(KEYINPUT13), .B(G475), .ZN(n472) );
  XNOR2_X1 U569 ( .A(n473), .B(n472), .ZN(n552) );
  NOR2_X1 U570 ( .A1(n553), .A2(n552), .ZN(n475) );
  INV_X1 U571 ( .A(KEYINPUT102), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n475), .B(n474), .ZN(n673) );
  INV_X1 U573 ( .A(n673), .ZN(n482) );
  NAND2_X1 U574 ( .A1(G234), .A2(n632), .ZN(n476) );
  XNOR2_X1 U575 ( .A(n477), .B(n476), .ZN(n515) );
  NAND2_X1 U576 ( .A1(G221), .A2(n515), .ZN(n479) );
  INV_X1 U577 ( .A(KEYINPUT21), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n479), .B(n478), .ZN(n684) );
  INV_X1 U579 ( .A(KEYINPUT98), .ZN(n480) );
  XNOR2_X1 U580 ( .A(n684), .B(n480), .ZN(n534) );
  INV_X1 U581 ( .A(n534), .ZN(n481) );
  NAND2_X1 U582 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U583 ( .A(n484), .B(KEYINPUT22), .ZN(n520) );
  NAND2_X1 U584 ( .A1(G227), .A2(n393), .ZN(n485) );
  NAND2_X1 U585 ( .A1(n722), .A2(n514), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n593), .B(KEYINPUT1), .ZN(n535) );
  INV_X1 U587 ( .A(n535), .ZN(n521) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n491), .A2(G210), .ZN(n493) );
  XNOR2_X1 U590 ( .A(n493), .B(n492), .ZN(n496) );
  INV_X1 U591 ( .A(n494), .ZN(n495) );
  XNOR2_X1 U592 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U593 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U594 ( .A(n500), .B(n499), .ZN(n707) );
  OR2_X1 U595 ( .A1(n707), .A2(G902), .ZN(n501) );
  XNOR2_X2 U596 ( .A(n501), .B(G472), .ZN(n591) );
  NAND2_X1 U597 ( .A1(G221), .A2(n502), .ZN(n510) );
  XOR2_X1 U598 ( .A(KEYINPUT24), .B(G128), .Z(n504) );
  XNOR2_X1 U599 ( .A(G110), .B(G119), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n504), .B(n503), .ZN(n509) );
  INV_X1 U601 ( .A(n505), .ZN(n507) );
  XNOR2_X1 U602 ( .A(KEYINPUT95), .B(KEYINPUT75), .ZN(n506) );
  XNOR2_X1 U603 ( .A(n507), .B(n506), .ZN(n508) );
  INV_X1 U604 ( .A(n511), .ZN(n512) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n765) );
  NAND2_X1 U606 ( .A1(n659), .A2(n514), .ZN(n518) );
  NAND2_X1 U607 ( .A1(n515), .A2(G217), .ZN(n516) );
  XNOR2_X1 U608 ( .A(n516), .B(KEYINPUT25), .ZN(n517) );
  XNOR2_X2 U609 ( .A(n518), .B(n517), .ZN(n589) );
  INV_X1 U610 ( .A(n589), .ZN(n683) );
  BUF_X1 U611 ( .A(n520), .Z(n525) );
  INV_X1 U612 ( .A(n521), .ZN(n680) );
  INV_X1 U613 ( .A(KEYINPUT89), .ZN(n522) );
  XNOR2_X1 U614 ( .A(n680), .B(n522), .ZN(n607) );
  XNOR2_X1 U615 ( .A(n591), .B(KEYINPUT6), .ZN(n602) );
  AND2_X1 U616 ( .A1(n602), .A2(n589), .ZN(n523) );
  AND2_X1 U617 ( .A1(n607), .A2(n523), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n525), .A2(n524), .ZN(n528) );
  INV_X1 U619 ( .A(KEYINPUT77), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n526), .B(KEYINPUT32), .ZN(n527) );
  INV_X1 U621 ( .A(KEYINPUT87), .ZN(n529) );
  NAND2_X1 U622 ( .A1(n563), .A2(KEYINPUT44), .ZN(n562) );
  INV_X1 U623 ( .A(n531), .ZN(n533) );
  AND2_X1 U624 ( .A1(n602), .A2(n683), .ZN(n532) );
  NAND2_X1 U625 ( .A1(n533), .A2(n532), .ZN(n662) );
  AND2_X2 U626 ( .A1(n535), .A2(n681), .ZN(n544) );
  NAND2_X1 U627 ( .A1(n544), .A2(n591), .ZN(n690) );
  INV_X1 U628 ( .A(KEYINPUT31), .ZN(n536) );
  NAND2_X1 U629 ( .A1(n681), .A2(n377), .ZN(n577) );
  OR2_X1 U630 ( .A1(n577), .A2(n591), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n652), .A2(n736), .ZN(n541) );
  INV_X1 U632 ( .A(n553), .ZN(n540) );
  NOR2_X1 U633 ( .A1(n552), .A2(n540), .ZN(n539) );
  XNOR2_X1 U634 ( .A(KEYINPUT101), .B(n539), .ZN(n740) );
  NAND2_X1 U635 ( .A1(n552), .A2(n540), .ZN(n744) );
  AND2_X1 U636 ( .A1(n740), .A2(n744), .ZN(n675) );
  XNOR2_X1 U637 ( .A(n675), .B(KEYINPUT79), .ZN(n584) );
  NAND2_X1 U638 ( .A1(n541), .A2(n584), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n662), .A2(n542), .ZN(n543) );
  XNOR2_X1 U640 ( .A(n544), .B(KEYINPUT105), .ZN(n545) );
  INV_X1 U641 ( .A(n545), .ZN(n547) );
  INV_X1 U642 ( .A(n602), .ZN(n546) );
  XNOR2_X1 U643 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n548) );
  NOR2_X1 U644 ( .A1(n364), .A2(n699), .ZN(n551) );
  XNOR2_X1 U645 ( .A(n551), .B(KEYINPUT34), .ZN(n555) );
  AND2_X1 U646 ( .A1(n553), .A2(n552), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT76), .ZN(n554) );
  NAND2_X1 U648 ( .A1(n555), .A2(n554), .ZN(n558) );
  INV_X1 U649 ( .A(KEYINPUT83), .ZN(n556) );
  XNOR2_X1 U650 ( .A(n556), .B(KEYINPUT35), .ZN(n557) );
  XNOR2_X2 U651 ( .A(n558), .B(n557), .ZN(n656) );
  INV_X1 U652 ( .A(KEYINPUT86), .ZN(n560) );
  BUF_X1 U653 ( .A(n563), .Z(n564) );
  INV_X1 U654 ( .A(n564), .ZN(n568) );
  INV_X1 U655 ( .A(n656), .ZN(n566) );
  INV_X1 U656 ( .A(KEYINPUT44), .ZN(n565) );
  AND2_X1 U657 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U659 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X2 U660 ( .A(n571), .B(KEYINPUT45), .ZN(n668) );
  NAND2_X1 U661 ( .A1(n675), .A2(KEYINPUT47), .ZN(n582) );
  NAND2_X1 U662 ( .A1(G953), .A2(n572), .ZN(n573) );
  NOR2_X1 U663 ( .A1(G900), .A2(n573), .ZN(n574) );
  XNOR2_X1 U664 ( .A(n574), .B(KEYINPUT106), .ZN(n575) );
  NOR2_X1 U665 ( .A1(n576), .A2(n575), .ZN(n587) );
  BUF_X1 U666 ( .A(n578), .Z(n613) );
  NAND2_X1 U667 ( .A1(n579), .A2(n613), .ZN(n580) );
  NOR2_X1 U668 ( .A1(n614), .A2(n580), .ZN(n650) );
  INV_X1 U669 ( .A(n650), .ZN(n581) );
  NAND2_X1 U670 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U671 ( .A(n583), .B(KEYINPUT78), .Z(n599) );
  INV_X1 U672 ( .A(n584), .ZN(n585) );
  NOR2_X1 U673 ( .A1(n585), .A2(KEYINPUT47), .ZN(n597) );
  INV_X1 U674 ( .A(n684), .ZN(n586) );
  NOR2_X1 U675 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U676 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U677 ( .A(KEYINPUT67), .B(n590), .Z(n601) );
  INV_X1 U678 ( .A(n591), .ZN(n688) );
  NOR2_X1 U679 ( .A1(n601), .A2(n688), .ZN(n592) );
  XNOR2_X1 U680 ( .A(n592), .B(KEYINPUT28), .ZN(n594) );
  NAND2_X1 U681 ( .A1(n594), .A2(n377), .ZN(n618) );
  BUF_X1 U682 ( .A(n595), .Z(n596) );
  NOR2_X1 U683 ( .A1(n618), .A2(n596), .ZN(n746) );
  NAND2_X1 U684 ( .A1(n597), .A2(n746), .ZN(n598) );
  AND2_X1 U685 ( .A1(n599), .A2(n598), .ZN(n612) );
  BUF_X1 U686 ( .A(n600), .Z(n604) );
  OR2_X1 U687 ( .A1(n601), .A2(n744), .ZN(n603) );
  NOR2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n623) );
  NAND2_X1 U689 ( .A1(n604), .A2(n623), .ZN(n606) );
  XOR2_X1 U690 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n605) );
  XNOR2_X1 U691 ( .A(n606), .B(n605), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n608), .A2(n607), .ZN(n750) );
  INV_X1 U693 ( .A(n746), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n609), .A2(KEYINPUT47), .ZN(n610) );
  AND2_X1 U695 ( .A1(n750), .A2(n610), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n622) );
  NOR2_X1 U697 ( .A1(n744), .A2(n627), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT40), .ZN(n780) );
  NAND2_X1 U699 ( .A1(n671), .A2(n670), .ZN(n676) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT41), .ZN(n700) );
  NOR2_X1 U701 ( .A1(n780), .A2(n778), .ZN(n620) );
  XNOR2_X1 U702 ( .A(n620), .B(n619), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n623), .A2(n670), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n680), .A2(n624), .ZN(n625) );
  XNOR2_X1 U705 ( .A(n625), .B(KEYINPUT43), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n626), .A2(n613), .ZN(n651) );
  OR2_X1 U707 ( .A1(n627), .A2(n740), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(KEYINPUT109), .ZN(n779) );
  INV_X1 U709 ( .A(n779), .ZN(n629) );
  AND2_X2 U710 ( .A1(n630), .A2(n629), .ZN(n768) );
  INV_X1 U711 ( .A(KEYINPUT2), .ZN(n664) );
  NOR2_X1 U712 ( .A1(n664), .A2(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n637) );
  INV_X1 U714 ( .A(n637), .ZN(n634) );
  INV_X1 U715 ( .A(n632), .ZN(n633) );
  OR2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n668), .A2(n635), .ZN(n642) );
  INV_X1 U718 ( .A(n636), .ZN(n640) );
  NAND2_X1 U719 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n638) );
  AND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  OR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U722 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X2 U723 ( .A1(n646), .A2(n732), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n648), .B(n647), .ZN(G63) );
  XNOR2_X1 U725 ( .A(G143), .B(KEYINPUT112), .ZN(n649) );
  XOR2_X1 U726 ( .A(n650), .B(n649), .Z(G45) );
  XOR2_X1 U727 ( .A(G140), .B(n651), .Z(G42) );
  NOR2_X1 U728 ( .A1(n654), .A2(n744), .ZN(n653) );
  XOR2_X1 U729 ( .A(G113), .B(n653), .Z(G15) );
  NOR2_X1 U730 ( .A1(n654), .A2(n740), .ZN(n655) );
  XOR2_X1 U731 ( .A(G116), .B(n655), .Z(G18) );
  XOR2_X1 U732 ( .A(G122), .B(n656), .Z(G24) );
  XNOR2_X1 U733 ( .A(n380), .B(G119), .ZN(G21) );
  AND2_X2 U734 ( .A1(n726), .A2(G217), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(n659), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n660), .A2(n732), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n661), .B(KEYINPUT120), .ZN(G66) );
  BUF_X1 U738 ( .A(n662), .Z(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(G101), .ZN(G3) );
  NAND2_X1 U740 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U741 ( .A1(KEYINPUT2), .A2(KEYINPUT80), .ZN(n667) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT114), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n679), .A2(n363), .ZN(n695) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT50), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U751 ( .A(n685), .B(KEYINPUT49), .Z(n686) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n691) );
  AND2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U755 ( .A(KEYINPUT51), .B(n692), .Z(n693) );
  NOR2_X1 U756 ( .A1(n700), .A2(n693), .ZN(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U758 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n700), .A2(n363), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U762 ( .A(KEYINPUT115), .B(n703), .Z(n704) );
  XNOR2_X1 U763 ( .A(n705), .B(G110), .ZN(G12) );
  NAND2_X1 U764 ( .A1(n376), .A2(G472), .ZN(n709) );
  XNOR2_X1 U765 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X2 U767 ( .A1(n710), .A2(n732), .ZN(n712) );
  XNOR2_X1 U768 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n712), .B(n711), .ZN(G57) );
  NAND2_X1 U770 ( .A1(n376), .A2(G475), .ZN(n716) );
  XNOR2_X1 U771 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X2 U773 ( .A1(n717), .A2(n732), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n718), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U775 ( .A1(n375), .A2(G469), .ZN(n724) );
  XOR2_X1 U776 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n720) );
  XNOR2_X1 U777 ( .A(KEYINPUT118), .B(KEYINPUT117), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U779 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U781 ( .A1(n725), .A2(n732), .ZN(G54) );
  NAND2_X1 U782 ( .A1(n376), .A2(G210), .ZN(n731) );
  BUF_X1 U783 ( .A(n727), .Z(n728) );
  XNOR2_X1 U784 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n729) );
  XNOR2_X1 U785 ( .A(n731), .B(n730), .ZN(n733) );
  NOR2_X2 U786 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n734), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U788 ( .A1(n736), .A2(n744), .ZN(n735) );
  XOR2_X1 U789 ( .A(G104), .B(n735), .Z(G6) );
  NOR2_X1 U790 ( .A1(n736), .A2(n740), .ZN(n738) );
  XNOR2_X1 U791 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n737) );
  XNOR2_X1 U792 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U793 ( .A(G107), .B(n739), .ZN(G9) );
  XOR2_X1 U794 ( .A(G128), .B(KEYINPUT29), .Z(n743) );
  INV_X1 U795 ( .A(n740), .ZN(n741) );
  NAND2_X1 U796 ( .A1(n746), .A2(n741), .ZN(n742) );
  XNOR2_X1 U797 ( .A(n743), .B(n742), .ZN(G30) );
  XOR2_X1 U798 ( .A(G146), .B(KEYINPUT113), .Z(n748) );
  INV_X1 U799 ( .A(n744), .ZN(n745) );
  NAND2_X1 U800 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U801 ( .A(n748), .B(n747), .ZN(G48) );
  XOR2_X1 U802 ( .A(G125), .B(KEYINPUT37), .Z(n749) );
  XNOR2_X1 U803 ( .A(n750), .B(n749), .ZN(G27) );
  NAND2_X1 U804 ( .A1(n751), .A2(n393), .ZN(n755) );
  NAND2_X1 U805 ( .A1(G953), .A2(G224), .ZN(n752) );
  XNOR2_X1 U806 ( .A(KEYINPUT61), .B(n752), .ZN(n753) );
  NAND2_X1 U807 ( .A1(n753), .A2(G898), .ZN(n754) );
  NAND2_X1 U808 ( .A1(n755), .A2(n754), .ZN(n763) );
  XNOR2_X1 U809 ( .A(n756), .B(KEYINPUT121), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U811 ( .A(n759), .B(G101), .ZN(n760) );
  NOR2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(G69) );
  XNOR2_X1 U814 ( .A(n764), .B(KEYINPUT122), .ZN(n766) );
  XNOR2_X1 U815 ( .A(n766), .B(n765), .ZN(n771) );
  XNOR2_X1 U816 ( .A(KEYINPUT123), .B(n771), .ZN(n767) );
  XNOR2_X1 U817 ( .A(n768), .B(n767), .ZN(n769) );
  NAND2_X1 U818 ( .A1(n393), .A2(n769), .ZN(n770) );
  XNOR2_X1 U819 ( .A(n770), .B(KEYINPUT124), .ZN(n775) );
  XNOR2_X1 U820 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U822 ( .A1(G953), .A2(n773), .ZN(n774) );
  NAND2_X1 U823 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U824 ( .A(KEYINPUT125), .B(n776), .Z(G72) );
  XOR2_X1 U825 ( .A(G137), .B(KEYINPUT126), .Z(n777) );
  XNOR2_X1 U826 ( .A(n778), .B(n777), .ZN(G39) );
  XOR2_X1 U827 ( .A(G134), .B(n779), .Z(G36) );
  XOR2_X1 U828 ( .A(n780), .B(G131), .Z(G33) );
endmodule

