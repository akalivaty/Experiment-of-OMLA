//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g0013(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n202), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT68), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n206), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n210), .B(new_n221), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n216), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G116), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n255), .A2(new_n257), .A3(new_n216), .A4(G87), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT22), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(KEYINPUT76), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT76), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n263), .A3(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G87), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n259), .A2(new_n265), .A3(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n255), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT85), .B1(new_n216), .B2(G107), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT23), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT23), .ZN(new_n270));
  OAI211_X1 g0070(.A(KEYINPUT85), .B(new_n270), .C1(new_n216), .C2(G107), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n260), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT24), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n214), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT66), .B1(G1), .B2(G13), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n260), .A2(new_n267), .A3(KEYINPUT24), .A4(new_n272), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT87), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G13), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT86), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT25), .ZN(new_n287));
  AOI21_X1  g0087(.A(G107), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n285), .B(new_n288), .C1(new_n286), .C2(new_n287), .ZN(new_n289));
  OAI211_X1 g0089(.A(KEYINPUT86), .B(KEYINPUT25), .C1(new_n284), .C2(G107), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G107), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n279), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n282), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n276), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n213), .B2(new_n214), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(G107), .A3(new_n292), .A4(new_n284), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n299), .A2(KEYINPUT87), .A3(new_n290), .A4(new_n289), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n281), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G294), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT70), .B(G1698), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n304), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n264), .A2(new_n255), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G41), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n213), .A2(new_n214), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(G1), .A3(G13), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n283), .A2(G45), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT5), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(G41), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(KEYINPUT80), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT80), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT5), .ZN(new_n318));
  AOI21_X1  g0118(.A(G41), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT81), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI211_X1 g0121(.A(KEYINPUT81), .B(G41), .C1(new_n316), .C2(new_n318), .ZN(new_n322));
  OAI211_X1 g0122(.A(G264), .B(new_n312), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n316), .A2(new_n318), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT81), .B1(new_n324), .B2(G41), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n320), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n312), .A2(G274), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n315), .A4(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n311), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n311), .A2(new_n323), .A3(new_n332), .A4(new_n328), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n302), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT88), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n302), .A2(new_n331), .A3(KEYINPUT88), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(G200), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n311), .A2(new_n323), .A3(G190), .A4(new_n328), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n338), .A2(new_n301), .A3(new_n281), .A4(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n251), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(G20), .B2(G77), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(G20), .A2(G33), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n298), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n298), .B1(G1), .B2(new_n216), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n284), .A2(G77), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n283), .B1(G41), .B2(G45), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(new_n312), .A3(G274), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n312), .A2(new_n356), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n359), .B1(G244), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n304), .A2(G232), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT3), .B(G33), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G238), .A2(G1698), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n255), .A2(new_n257), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n294), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(KEYINPUT71), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n310), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT71), .B1(new_n366), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n362), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n355), .B1(new_n372), .B2(new_n330), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n372), .A2(G179), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n373), .B2(new_n374), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n355), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n372), .B2(G200), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n372), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g0185(.A(new_n385), .B(KEYINPUT73), .Z(new_n386));
  NAND2_X1  g0186(.A1(new_n203), .A2(G20), .ZN(new_n387));
  INV_X1    g0187(.A(G150), .ZN(new_n388));
  INV_X1    g0188(.A(new_n348), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n387), .B1(new_n388), .B2(new_n389), .C1(new_n251), .C2(new_n346), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(new_n279), .B1(new_n244), .B2(new_n285), .ZN(new_n391));
  INV_X1    g0191(.A(new_n351), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G50), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n304), .A2(G222), .ZN(new_n395));
  INV_X1    g0195(.A(G223), .ZN(new_n396));
  INV_X1    g0196(.A(G1698), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n364), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n310), .B1(G77), .B2(new_n364), .C1(new_n395), .C2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n359), .B1(G226), .B2(new_n361), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n330), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n332), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n394), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n401), .A2(new_n383), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(G200), .B2(new_n401), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT9), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n391), .A2(new_n408), .A3(new_n393), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n391), .B2(new_n393), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT10), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n407), .B(new_n413), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n405), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n304), .A2(G226), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G232), .A2(G1698), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n367), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G97), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n310), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n359), .B1(G238), .B2(new_n361), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n421), .B2(new_n422), .ZN(new_n425));
  OAI21_X1  g0225(.A(G169), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT14), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n421), .A2(new_n422), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(KEYINPUT14), .A3(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n431), .B(KEYINPUT74), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n425), .A2(new_n332), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G68), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G20), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n440), .B1(new_n251), .B2(new_n352), .C1(new_n389), .C2(new_n244), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n279), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT75), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT11), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n442), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n283), .A2(KEYINPUT12), .A3(G13), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n285), .A2(KEYINPUT12), .B1(new_n440), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n351), .A2(KEYINPUT12), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G68), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n445), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n438), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n432), .A2(G200), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n424), .B(KEYINPUT74), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n430), .A2(G190), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n453), .B(new_n456), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n415), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n347), .A2(new_n284), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n392), .B2(new_n347), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n255), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G33), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT7), .B1(new_n466), .B2(G20), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(new_n264), .B2(new_n255), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT7), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n470), .A3(G68), .ZN(new_n471));
  AND2_X1   g0271(.A1(G58), .A2(G68), .ZN(new_n472));
  OAI21_X1  g0272(.A(G20), .B1(new_n472), .B2(new_n202), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n348), .A2(G159), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(KEYINPUT77), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT77), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT16), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n298), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n469), .A2(G20), .ZN(new_n481));
  AOI21_X1  g0281(.A(G33), .B1(new_n261), .B2(new_n263), .ZN(new_n482));
  INV_X1    g0282(.A(new_n257), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n469), .B1(new_n364), .B2(G20), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n439), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n473), .A2(new_n474), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT77), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n475), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n478), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n463), .B1(new_n480), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n361), .A2(G232), .B1(new_n327), .B2(new_n357), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n397), .A2(KEYINPUT70), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT70), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G1698), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n496), .A3(G223), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G226), .A2(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n466), .A2(new_n499), .B1(G33), .B2(G87), .ZN(new_n500));
  OAI211_X1 g0300(.A(G179), .B(new_n493), .C1(new_n500), .C2(new_n309), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n358), .B1(new_n360), .B2(new_n236), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n304), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n503), .A2(new_n306), .B1(new_n254), .B2(new_n265), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(new_n310), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n501), .B1(new_n505), .B2(new_n330), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT18), .B1(new_n492), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n471), .A2(new_n479), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n491), .A3(new_n279), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n462), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT18), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(new_n506), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT17), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n383), .A2(KEYINPUT78), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n383), .A2(KEYINPUT78), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n517), .B(new_n493), .C1(new_n500), .C2(new_n309), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n505), .B2(G200), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n514), .B1(new_n492), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g0320(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n521));
  AND4_X1   g0321(.A1(new_n510), .A2(new_n462), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n508), .B(new_n513), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n386), .A2(new_n460), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G303), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n364), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n494), .A2(new_n496), .A3(G257), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G264), .A2(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n528), .B1(new_n466), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT83), .B1(new_n532), .B2(new_n309), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n367), .A2(G303), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n304), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n306), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(new_n310), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G270), .B(new_n312), .C1(new_n321), .C2(new_n322), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n540), .A2(new_n328), .ZN(new_n541));
  INV_X1    g0341(.A(new_n517), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT20), .ZN(new_n544));
  AOI21_X1  g0344(.A(G20), .B1(G33), .B2(G283), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n254), .A2(G97), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT84), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n545), .B2(new_n546), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n252), .A2(G20), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n279), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n544), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n550), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n548), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n215), .A2(new_n276), .B1(G20), .B2(new_n252), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n284), .A2(G116), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n279), .A2(new_n293), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(G116), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n540), .A2(new_n328), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n533), .B2(new_n538), .ZN(new_n566));
  INV_X1    g0366(.A(G200), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n543), .B(new_n564), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(G179), .A3(new_n563), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n539), .A2(new_n541), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n330), .B1(new_n559), .B2(new_n562), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n570), .B2(new_n571), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n568), .B(new_n569), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G257), .B(new_n312), .C1(new_n321), .C2(new_n322), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n328), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n264), .A2(G244), .A3(new_n255), .A4(new_n304), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G283), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT4), .A4(G244), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G250), .A2(G1698), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n364), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n310), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n579), .A2(new_n332), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n580), .A2(new_n581), .B1(G33), .B2(G283), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n309), .B1(new_n591), .B2(new_n587), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n330), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT6), .ZN(new_n594));
  INV_X1    g0394(.A(G97), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(new_n294), .ZN(new_n596));
  NOR2_X1   g0396(.A1(G97), .A2(G107), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n294), .A2(KEYINPUT6), .A3(G97), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n600), .A2(new_n216), .B1(new_n352), .B2(new_n389), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n294), .B1(new_n484), .B2(new_n485), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n279), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n284), .A2(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n561), .B2(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n590), .A2(new_n593), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n313), .A2(G274), .ZN(new_n608));
  INV_X1    g0408(.A(G250), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n313), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n312), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n254), .A2(new_n252), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n494), .A2(new_n496), .A3(G238), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G244), .A2(G1698), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n466), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(G179), .B(new_n611), .C1(new_n616), .C2(new_n309), .ZN(new_n617));
  INV_X1    g0417(.A(new_n611), .ZN(new_n618));
  INV_X1    g0418(.A(new_n612), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n304), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n306), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n621), .B2(new_n310), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n617), .B1(new_n622), .B2(new_n330), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT82), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n617), .B(KEYINPUT82), .C1(new_n622), .C2(new_n330), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n264), .A2(new_n216), .A3(G68), .A4(new_n255), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT19), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n419), .B2(new_n216), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n265), .A2(new_n595), .A3(new_n294), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n216), .A2(G33), .A3(G97), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n629), .A2(new_n630), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n298), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n343), .A2(new_n284), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n561), .A2(new_n343), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n625), .A2(new_n626), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n579), .A2(G190), .A3(new_n589), .ZN(new_n641));
  INV_X1    g0441(.A(new_n605), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n598), .A2(new_n599), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(G20), .B1(G77), .B2(new_n348), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n484), .A2(new_n485), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n294), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n642), .B1(new_n646), .B2(new_n279), .ZN(new_n647));
  OAI21_X1  g0447(.A(G200), .B1(new_n592), .B2(new_n578), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n641), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n279), .A2(new_n293), .A3(new_n265), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n633), .A2(new_n635), .A3(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(G190), .B(new_n611), .C1(new_n616), .C2(new_n309), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n651), .B(new_n652), .C1(new_n567), .C2(new_n622), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n607), .A2(new_n640), .A3(new_n649), .A4(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n341), .A2(new_n526), .A3(new_n576), .A4(new_n654), .ZN(G372));
  NAND2_X1  g0455(.A1(new_n412), .A2(new_n414), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n520), .A2(new_n522), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n379), .A2(new_n459), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n455), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n508), .A2(new_n513), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n404), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n590), .A2(new_n593), .A3(new_n606), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n623), .A2(KEYINPUT89), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n617), .B(new_n665), .C1(new_n622), .C2(new_n330), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n639), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n663), .A2(new_n667), .A3(new_n668), .A4(new_n653), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n667), .ZN(new_n670));
  INV_X1    g0470(.A(new_n653), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n638), .B1(new_n623), .B2(new_n624), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n626), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n668), .B1(new_n673), .B2(new_n663), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n334), .B(new_n569), .C1(new_n573), .C2(new_n574), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n607), .A2(new_n649), .A3(new_n340), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n638), .B1(new_n623), .B2(KEYINPUT89), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n678), .B2(new_n666), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n662), .B1(new_n525), .B2(new_n682), .ZN(G369));
  OAI21_X1  g0483(.A(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n283), .A2(new_n216), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(G213), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT90), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n564), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n575), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n689), .B(KEYINPUT90), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n302), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n341), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n334), .A2(new_n691), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT92), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n684), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n698), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n702), .A2(KEYINPUT92), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT92), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n700), .B2(new_n701), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n706), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n334), .A2(new_n698), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n704), .A2(new_n710), .A3(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n207), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  OR3_X1    g0514(.A1(new_n713), .A2(new_n714), .A3(G41), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n713), .B2(G41), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n630), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n219), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n698), .B1(new_n675), .B2(new_n680), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n679), .A2(new_n340), .A3(new_n607), .A4(new_n649), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n336), .A2(new_n337), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n705), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n667), .A2(new_n653), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT26), .B1(new_n726), .B2(new_n607), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n673), .A2(new_n668), .A3(new_n663), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n667), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n691), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  MUX2_X1   g0530(.A(new_n722), .B(new_n730), .S(KEYINPUT29), .Z(new_n731));
  NAND3_X1  g0531(.A1(new_n589), .A2(new_n328), .A3(new_n577), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n622), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n570), .A2(new_n732), .A3(new_n329), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n592), .A2(new_n578), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n311), .A2(new_n323), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n617), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n566), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n566), .A2(new_n738), .A3(new_n736), .A4(KEYINPUT30), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n611), .B1(new_n616), .B2(new_n309), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n329), .A2(new_n332), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT94), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n570), .A4(new_n732), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n735), .A2(new_n741), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n698), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n741), .A2(new_n742), .A3(new_n734), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n691), .A2(new_n749), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n576), .A2(new_n341), .A3(new_n654), .A4(new_n691), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n696), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n731), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n721), .B1(new_n755), .B2(G1), .ZN(G364));
  OR2_X1    g0556(.A1(new_n697), .A2(KEYINPUT95), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n697), .A2(KEYINPUT95), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n717), .ZN(new_n760));
  INV_X1    g0560(.A(G13), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n283), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n695), .B2(new_n696), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT96), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n695), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n765), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n216), .A2(new_n332), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n567), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G68), .A2(new_n777), .B1(new_n779), .B2(G77), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n517), .A2(new_n776), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G58), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n517), .A2(new_n778), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n780), .B1(new_n244), .B2(new_n782), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n216), .A2(G179), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n383), .A3(new_n567), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n787), .A2(new_n383), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n294), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n367), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n265), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n383), .A2(G179), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n216), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n796), .B1(G97), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n791), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n784), .A2(G322), .B1(new_n779), .B2(G311), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  INV_X1    g0603(.A(new_n777), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT33), .B(G317), .Z(new_n805));
  OAI221_X1 g0605(.A(new_n802), .B1(new_n803), .B2(new_n792), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n781), .A2(G326), .B1(new_n799), .B2(G294), .ZN(new_n807));
  INV_X1    g0607(.A(new_n788), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n364), .B1(new_n808), .B2(G329), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(new_n527), .C2(new_n795), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n786), .A2(new_n801), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n215), .B1(G20), .B2(new_n330), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n774), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n772), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n364), .A2(new_n207), .ZN(new_n816));
  INV_X1    g0616(.A(G355), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(G116), .B2(new_n207), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n246), .A2(G45), .ZN(new_n819));
  INV_X1    g0619(.A(G45), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n713), .B(new_n466), .C1(new_n820), .C2(new_n220), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n773), .B(new_n813), .C1(new_n815), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n769), .A2(new_n823), .ZN(G396));
  NOR3_X1   g0624(.A1(new_n691), .A2(new_n355), .A3(KEYINPUT99), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT99), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n381), .B2(new_n698), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n384), .B(new_n828), .C1(new_n376), .C2(new_n378), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n373), .A2(new_n374), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n691), .A2(new_n355), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n830), .A2(new_n375), .A3(new_n377), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n722), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n663), .A2(new_n640), .A3(new_n653), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT26), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(new_n667), .A3(new_n669), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n833), .B(new_n691), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n754), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n834), .A2(new_n754), .A3(new_n839), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n774), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n840), .B1(new_n842), .B2(KEYINPUT100), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(KEYINPUT100), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n812), .A2(new_n770), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n765), .B1(G77), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT97), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n781), .A2(G303), .B1(new_n779), .B2(G116), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n803), .B2(new_n804), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT98), .Z(new_n851));
  INV_X1    g0651(.A(new_n795), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n784), .A2(G294), .B1(G107), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n799), .A2(G97), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n364), .B1(new_n808), .B2(G311), .ZN(new_n855));
  INV_X1    g0655(.A(new_n792), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(G87), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n781), .A2(G137), .B1(new_n779), .B2(G159), .ZN(new_n860));
  INV_X1    g0660(.A(G143), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n861), .B2(new_n785), .C1(new_n388), .C2(new_n804), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(G68), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n864), .B1(new_n244), .B2(new_n795), .C1(new_n783), .C2(new_n798), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n306), .B(new_n865), .C1(G132), .C2(new_n808), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n859), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n812), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n848), .B1(new_n867), .B2(new_n868), .C1(new_n833), .C2(new_n771), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n844), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  NOR3_X1   g0671(.A1(new_n219), .A2(new_n352), .A3(new_n472), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(KEYINPUT102), .B1(G68), .B2(new_n201), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(KEYINPUT102), .B2(new_n873), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(G1), .A3(new_n761), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT103), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT36), .ZN(new_n878));
  OAI211_X1 g0678(.A(G116), .B(new_n217), .C1(new_n643), .C2(KEYINPUT35), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n879), .A2(KEYINPUT101), .B1(KEYINPUT35), .B2(new_n643), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(KEYINPUT101), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n877), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n878), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n454), .A2(new_n698), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n428), .A2(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n459), .B(new_n884), .C1(new_n885), .C2(new_n453), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n438), .A2(new_n454), .A3(new_n698), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n380), .A2(new_n698), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n839), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT104), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n510), .A2(new_n462), .A3(new_n519), .ZN(new_n894));
  OAI21_X1  g0694(.A(G68), .B1(new_n468), .B2(new_n469), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n466), .A2(KEYINPUT7), .A3(G20), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n478), .B1(new_n897), .B2(new_n490), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n463), .B1(new_n898), .B2(new_n480), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n894), .B1(new_n899), .B2(new_n507), .ZN(new_n900));
  INV_X1    g0700(.A(new_n688), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n511), .A2(new_n506), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n511), .A2(new_n688), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n894), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n523), .A2(new_n902), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n892), .A2(new_n893), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n890), .B1(new_n722), .B2(new_n833), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n913), .A2(KEYINPUT104), .A3(new_n889), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n660), .A2(new_n901), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT39), .B1(new_n910), .B2(new_n911), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n894), .B1(new_n492), .B2(new_n507), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n492), .A2(new_n901), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n907), .A2(new_n922), .B1(new_n523), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n918), .B(new_n919), .C1(KEYINPUT38), .C2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n438), .A2(new_n454), .A3(new_n691), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n916), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n526), .A2(new_n731), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n662), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n748), .A2(new_n749), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n753), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n526), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT105), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n922), .A2(new_n907), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n523), .A2(new_n921), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n910), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n918), .B(KEYINPUT105), .C1(KEYINPUT38), .C2(new_n923), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n886), .A2(new_n887), .B1(new_n829), .B2(new_n832), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n934), .A2(KEYINPUT40), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n934), .B(new_n943), .C1(new_n910), .C2(new_n911), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n935), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n935), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(G330), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n931), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n283), .B2(new_n762), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n931), .A2(new_n952), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n883), .B1(new_n954), .B2(new_n955), .ZN(G367));
  OAI211_X1 g0756(.A(new_n607), .B(new_n649), .C1(new_n647), .C2(new_n691), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n663), .A2(new_n698), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n703), .A2(new_n706), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT106), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT42), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n960), .B2(KEYINPUT42), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n724), .A2(new_n957), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n698), .B1(new_n965), .B2(new_n607), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n960), .B2(KEYINPUT42), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n691), .A2(new_n651), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n667), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n679), .B2(new_n970), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n968), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n959), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n704), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n964), .A2(new_n973), .A3(new_n972), .A4(new_n967), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n979), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n717), .B(KEYINPUT41), .ZN(new_n984));
  INV_X1    g0784(.A(new_n704), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n710), .A2(new_n711), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT107), .B1(new_n986), .B2(new_n978), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT107), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n710), .A2(new_n988), .A3(new_n711), .A4(new_n959), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n991), .A3(new_n978), .ZN(new_n992));
  INV_X1    g0792(.A(new_n986), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT44), .B1(new_n993), .B2(new_n959), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT45), .B1(new_n987), .B2(new_n989), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n985), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n994), .A2(new_n992), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n987), .A2(new_n989), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n998), .A2(new_n1001), .A3(new_n704), .A4(new_n990), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n703), .B(new_n706), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n697), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n757), .A3(new_n758), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n755), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n997), .A2(new_n1002), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n984), .B1(new_n1009), .B2(new_n755), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n983), .B1(new_n1010), .B2(new_n764), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n814), .B1(new_n207), .B2(new_n342), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n466), .A2(new_n713), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n240), .B2(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n782), .A2(new_n861), .B1(new_n439), .B2(new_n798), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G159), .B2(new_n777), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n364), .B1(new_n792), .B2(new_n352), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT109), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n784), .A2(G150), .B1(G137), .B2(new_n808), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n201), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n779), .A2(new_n1020), .B1(new_n852), .B2(G58), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(G294), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n779), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n804), .A2(new_n1023), .B1(new_n1024), .B2(new_n803), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT46), .B1(new_n852), .B2(G116), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n852), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G303), .A2(new_n784), .B1(new_n781), .B2(G311), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n294), .C2(new_n798), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n306), .B1(new_n595), .B2(new_n792), .C1(new_n1031), .C2(new_n788), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT108), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1022), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n774), .B(new_n1014), .C1(new_n1036), .C2(new_n812), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n772), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n975), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1011), .A2(new_n1039), .ZN(G387));
  NAND3_X1  g0840(.A1(new_n1005), .A2(new_n764), .A3(new_n1006), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n816), .A2(new_n718), .B1(G107), .B2(new_n207), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n237), .A2(G45), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n718), .A2(KEYINPUT111), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n820), .B1(new_n439), .B2(new_n352), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n718), .B2(KEYINPUT111), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(G50), .B2(new_n346), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n347), .A2(new_n1047), .A3(new_n244), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1044), .A2(new_n1046), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1051), .A2(new_n1013), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1042), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n765), .B1(new_n1053), .B2(new_n815), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1024), .A2(new_n439), .B1(new_n795), .B2(new_n352), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n347), .B2(new_n777), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n306), .B1(G150), .B2(new_n808), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n781), .A2(G159), .B1(G97), .B2(new_n856), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n784), .A2(G50), .B1(new_n799), .B2(new_n343), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n466), .B1(G326), .B2(new_n808), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n781), .A2(G322), .B1(new_n777), .B2(G311), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n527), .B2(new_n1024), .C1(new_n1031), .C2(new_n785), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n799), .A2(G283), .B1(new_n852), .B2(G294), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT49), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT113), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1061), .B1(new_n252), .B2(new_n792), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1069), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1060), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1054), .B1(new_n1074), .B2(new_n812), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n703), .B2(new_n1038), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1007), .A2(new_n760), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n755), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1041), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  NAND3_X1  g0879(.A1(new_n997), .A2(new_n1002), .A3(new_n764), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n814), .B1(new_n595), .B2(new_n207), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n249), .B2(new_n1013), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G311), .A2(new_n784), .B1(new_n781), .B2(G317), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT52), .Z(new_n1084));
  AOI211_X1 g0884(.A(new_n364), .B(new_n793), .C1(G322), .C2(new_n808), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G303), .A2(new_n777), .B1(new_n779), .B2(G294), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n799), .A2(G116), .B1(new_n852), .B2(G283), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G150), .A2(new_n781), .B1(new_n784), .B2(G159), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n804), .A2(new_n201), .B1(new_n1024), .B2(new_n346), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n798), .A2(new_n352), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n788), .A2(new_n861), .B1(new_n795), .B2(new_n439), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT114), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1093), .A2(new_n466), .A3(new_n857), .A4(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n774), .B(new_n1082), .C1(new_n1097), .C2(new_n812), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n959), .B2(new_n1038), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1080), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1009), .A2(new_n760), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n997), .A2(new_n1002), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1007), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  OAI211_X1 g0905(.A(new_n691), .B(new_n833), .C1(new_n725), .C2(new_n729), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n891), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT115), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n886), .A2(new_n887), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n942), .A3(new_n926), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n926), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n917), .B(new_n924), .C1(new_n892), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n754), .A2(new_n833), .A3(new_n888), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n926), .B1(new_n913), .B2(new_n889), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1114), .B1(new_n940), .B2(new_n941), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1118), .A2(new_n925), .B1(new_n1119), .B2(new_n1112), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT31), .B1(new_n747), .B2(new_n698), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n696), .B1(new_n1123), .B2(new_n753), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n943), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1117), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(new_n763), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n765), .B1(new_n347), .B2(new_n846), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n777), .A2(G137), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n367), .B(new_n1129), .C1(G125), .C2(new_n808), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n784), .A2(G132), .B1(new_n799), .B2(G159), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n781), .A2(G128), .B1(new_n1020), .B2(new_n856), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  NAND2_X1  g0933(.A1(new_n779), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n852), .A2(G150), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n364), .B(new_n796), .C1(G294), .C2(new_n808), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1092), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G116), .A2(new_n784), .B1(new_n781), .B2(G283), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1138), .A2(new_n864), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G107), .A2(new_n777), .B1(new_n779), .B2(G97), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT117), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1135), .A2(new_n1137), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1128), .B1(new_n1144), .B2(new_n812), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n925), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n771), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1127), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n833), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n934), .A2(G330), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1107), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n1116), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT116), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n754), .A2(new_n833), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1156), .A2(new_n889), .B1(new_n1124), .B2(new_n943), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1157), .B2(new_n913), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n913), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1125), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n888), .B1(new_n754), .B2(new_n833), .ZN(new_n1161));
  OAI211_X1 g0961(.A(KEYINPUT116), .B(new_n1159), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1154), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n526), .A2(new_n1124), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n929), .A2(new_n1165), .A3(new_n662), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1167), .A2(new_n1126), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n717), .B1(new_n1167), .B2(new_n1126), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1148), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G378));
  AOI21_X1  g0971(.A(new_n696), .B1(new_n946), .B2(new_n947), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT121), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n945), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n945), .B2(new_n1172), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT120), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n415), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n415), .A2(new_n1176), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n415), .A2(new_n1176), .ZN(new_n1182));
  AOI211_X1 g0982(.A(KEYINPUT120), .B(new_n405), .C1(new_n412), .C2(new_n414), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n394), .A2(new_n688), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1181), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1174), .A2(new_n1175), .A3(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n945), .A2(new_n1172), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1191), .A2(new_n1192), .A3(KEYINPUT121), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1190), .A2(new_n1193), .A3(new_n928), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n915), .A2(new_n927), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(KEYINPUT121), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n945), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n1191), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1174), .B1(new_n1175), .B2(new_n1189), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1194), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n764), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1189), .A2(new_n770), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n784), .A2(G107), .B1(new_n777), .B2(G97), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n342), .B2(new_n1024), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n781), .A2(G116), .B1(G77), .B2(new_n852), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n466), .A2(G41), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n799), .A2(G68), .B1(new_n808), .B2(G283), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n792), .A2(new_n783), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT118), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1205), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1207), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n244), .C1(G33), .C2(G41), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G125), .A2(new_n781), .B1(new_n784), .B2(G128), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n799), .A2(G150), .B1(new_n852), .B2(new_n1133), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G132), .A2(new_n777), .B1(new_n779), .B2(G137), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n856), .A2(G159), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n808), .C2(G124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1218), .B1(new_n1223), .B2(new_n1227), .C1(new_n1214), .C2(new_n1212), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n812), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n845), .A2(new_n201), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1203), .A2(new_n765), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1202), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n928), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1198), .A2(new_n1199), .A3(new_n1195), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1166), .B1(new_n1163), .B2(new_n1126), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1233), .A2(KEYINPUT57), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n760), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1237), .A2(KEYINPUT122), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT122), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1236), .A2(new_n1241), .A3(new_n760), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1232), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G375));
  INV_X1    g1044(.A(new_n984), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n929), .A2(new_n1165), .A3(new_n662), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1163), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1167), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G132), .A2(new_n781), .B1(new_n784), .B2(G137), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n777), .A2(new_n1133), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT124), .Z(new_n1252));
  AOI22_X1  g1052(.A1(G50), .A2(new_n799), .B1(new_n779), .B2(G150), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n789), .B2(new_n795), .ZN(new_n1254));
  INV_X1    g1054(.A(G128), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n466), .B1(new_n1255), .B2(new_n788), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1254), .A2(new_n1211), .A3(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n782), .A2(new_n1023), .B1(new_n804), .B2(new_n252), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n364), .B1(new_n856), .B2(G77), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n342), .B2(new_n798), .C1(new_n785), .C2(new_n803), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G107), .C2(new_n779), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n788), .A2(new_n527), .B1(new_n795), .B2(new_n595), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT123), .Z(new_n1263));
  AOI22_X1  g1063(.A1(new_n1252), .A2(new_n1257), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n765), .B1(G68), .B2(new_n846), .C1(new_n1264), .C2(new_n868), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1149), .B2(new_n770), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1164), .B2(new_n764), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1248), .A2(new_n1267), .ZN(G381));
  AND3_X1   g1068(.A1(new_n1011), .A2(new_n1104), .A3(new_n1039), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G396), .A2(G393), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n870), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1271), .A2(G378), .A3(G381), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1272), .A3(new_n1243), .ZN(G407));
  INV_X1    g1073(.A(G343), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(G213), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1243), .A2(new_n1170), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G407), .A2(G213), .A3(new_n1277), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1278), .B(KEYINPUT125), .Z(G409));
  AOI211_X1 g1079(.A(new_n1170), .B(new_n1232), .C1(new_n1240), .C2(new_n1242), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT126), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1194), .B2(new_n1200), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1233), .A2(KEYINPUT126), .A3(new_n1234), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1282), .A2(new_n764), .A3(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1231), .B1(new_n1239), .B2(new_n984), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1170), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1275), .B1(new_n1280), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1247), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n1246), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1290), .A2(new_n1167), .A3(new_n760), .A4(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G384), .A3(new_n1267), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G384), .B1(new_n1292), .B2(new_n1267), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G2897), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1275), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1295), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1293), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(G2897), .A3(new_n1276), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT61), .B1(new_n1288), .B2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1275), .B(new_n1296), .C1(new_n1280), .C2(new_n1287), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1104), .B1(new_n1011), .B2(new_n1039), .ZN(new_n1307));
  AND2_X1   g1107(.A1(G396), .A2(G393), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1308), .A2(new_n1270), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1269), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1309), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G387), .A2(G390), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1011), .A2(new_n1104), .A3(new_n1039), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1237), .A2(KEYINPUT122), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1239), .A2(new_n1238), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1242), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1232), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(G378), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1276), .B1(new_n1320), .B2(new_n1286), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1296), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1303), .A2(new_n1306), .A3(new_n1315), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1304), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1321), .A2(KEYINPUT62), .A3(new_n1296), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1326), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT127), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1309), .B1(new_n1269), .B2(new_n1307), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1312), .A2(new_n1313), .A3(new_n1311), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1331), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1323), .B1(new_n1330), .B2(new_n1336), .ZN(G405));
  NOR2_X1   g1137(.A1(new_n1243), .A2(G378), .ZN(new_n1338));
  OR3_X1    g1138(.A1(new_n1338), .A2(new_n1280), .A3(new_n1296), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1296), .B1(new_n1338), .B2(new_n1280), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1315), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1315), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(G402));
endmodule


