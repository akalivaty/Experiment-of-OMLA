//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1311, new_n1312, new_n1313, new_n1314, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI221_X1 g0009(.A(new_n206), .B1(new_n202), .B2(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n205), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n205), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT64), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n212), .A2(new_n214), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(new_n217), .A2(KEYINPUT1), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n219), .A2(new_n223), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n213), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  OR2_X1    g0052(.A1(new_n252), .A2(G264), .ZN(new_n253));
  INV_X1    g0053(.A(G257), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n252), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n251), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT66), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT66), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n249), .A2(new_n260), .A3(new_n250), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G303), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n256), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT85), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(KEYINPUT85), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n273), .B(G45), .C1(new_n266), .C2(KEYINPUT5), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  AND2_X1   g0076(.A1(G1), .A2(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n272), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n264), .A2(new_n265), .B1(new_n271), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n278), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n284));
  AOI21_X1  g0084(.A(G41), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(G270), .B(new_n282), .C1(new_n285), .C2(new_n274), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT88), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n265), .B1(new_n275), .B2(new_n269), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT88), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(G270), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n281), .A2(G190), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n273), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT72), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n297), .A2(new_n273), .A3(G13), .A4(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(new_n224), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n224), .ZN(new_n303));
  AOI211_X1 g0103(.A(KEYINPUT72), .B(new_n303), .C1(new_n296), .C2(new_n298), .ZN(new_n304));
  OAI211_X1 g0104(.A(G116), .B(new_n293), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G283), .ZN(new_n306));
  INV_X1    g0106(.A(G97), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n306), .B(new_n225), .C1(G33), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G116), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n303), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT20), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n312), .ZN(new_n314));
  INV_X1    g0114(.A(new_n299), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n313), .A2(new_n314), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n305), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n280), .A2(new_n271), .ZN(new_n318));
  INV_X1    g0118(.A(new_n256), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n263), .B1(new_n259), .B2(new_n261), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n265), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n291), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n292), .B(new_n317), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n305), .A2(new_n316), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(G179), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n305), .B2(new_n316), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT21), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n291), .A2(new_n318), .A3(new_n321), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n328), .B2(new_n330), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n324), .B(new_n326), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n252), .A2(G222), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G223), .A2(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n262), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n265), .C1(G77), .C2(new_n262), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n265), .A2(new_n276), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G45), .ZN(new_n341));
  AOI21_X1  g0141(.A(G1), .B1(new_n266), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n265), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(G226), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n323), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n338), .A2(G190), .A3(new_n344), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n201), .A2(new_n225), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT67), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT8), .B(G58), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n248), .A2(G20), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G20), .A2(G33), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n353), .A2(new_n354), .B1(G150), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n301), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT9), .ZN(new_n359));
  INV_X1    g0159(.A(new_n295), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n303), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n225), .A2(G1), .ZN(new_n362));
  INV_X1    g0162(.A(G50), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n361), .A2(new_n364), .B1(new_n363), .B2(new_n360), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n365), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT9), .B1(new_n357), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT73), .B(KEYINPUT10), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n369), .A2(new_n346), .A3(new_n347), .A4(new_n370), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n346), .A3(new_n347), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT10), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n371), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n358), .A2(new_n365), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT68), .A2(G179), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT68), .A2(G179), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n338), .A2(new_n381), .A3(new_n344), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(G169), .B1(new_n338), .B2(new_n344), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n343), .A2(G244), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n279), .A2(new_n342), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT69), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n259), .A2(new_n261), .ZN(new_n390));
  INV_X1    g0190(.A(G107), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G238), .A2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n213), .B2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n392), .B(new_n265), .C1(new_n390), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT69), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n386), .A2(new_n396), .A3(new_n387), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n381), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n327), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n302), .A2(new_n304), .B1(G1), .B2(new_n225), .ZN(new_n402));
  NOR2_X1   g0202(.A1(G13), .A2(G33), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n205), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n202), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT70), .ZN(new_n407));
  INV_X1    g0207(.A(new_n355), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n352), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n407), .B2(new_n408), .ZN(new_n410));
  INV_X1    g0210(.A(new_n354), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n303), .B1(new_n202), .B2(new_n315), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n400), .B(new_n401), .C1(new_n406), .C2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G190), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n398), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n406), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n398), .A2(G200), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n414), .A4(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n377), .A2(new_n385), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT75), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G232), .A2(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(G226), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n427), .B2(G1698), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n259), .A2(new_n261), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n248), .A2(new_n307), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n265), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n282), .A2(new_n339), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n387), .B1(new_n435), .B2(new_n215), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n282), .B1(new_n429), .B2(new_n431), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT13), .B1(new_n439), .B2(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G169), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n425), .B1(new_n442), .B2(KEYINPUT76), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n327), .B1(new_n438), .B2(new_n440), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n441), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n443), .A2(new_n446), .B1(G179), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n441), .A2(new_n425), .A3(G169), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n411), .A2(new_n202), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n408), .A2(new_n363), .B1(new_n225), .B2(G68), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n303), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT11), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n455), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n360), .A2(KEYINPUT12), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n315), .A2(KEYINPUT12), .A3(new_n214), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n214), .B1(new_n402), .B2(KEYINPUT12), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n447), .A2(G190), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n461), .B(new_n460), .C1(G200), .C2(new_n441), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n451), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT75), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n377), .A2(new_n466), .A3(new_n385), .A4(new_n422), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n352), .A2(new_n362), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n468), .A2(new_n361), .B1(new_n360), .B2(new_n352), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT7), .B1(new_n390), .B2(new_n225), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT7), .ZN(new_n471));
  NOR4_X1   g0271(.A1(new_n257), .A2(new_n258), .A3(new_n471), .A4(G20), .ZN(new_n472));
  OAI21_X1  g0272(.A(G68), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G58), .A2(G68), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT78), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G58), .A3(G68), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n477), .A3(new_n227), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G159), .B2(new_n355), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT16), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n257), .A2(new_n258), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT7), .B1(new_n481), .B2(new_n225), .ZN(new_n482));
  OAI21_X1  g0282(.A(G68), .B1(new_n482), .B2(new_n472), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(KEYINPUT16), .A3(new_n479), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n303), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n469), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G223), .A2(G1698), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n427), .B2(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n251), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n265), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n282), .A2(G232), .A3(new_n339), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n387), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n399), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n488), .A2(new_n251), .B1(G33), .B2(G87), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT79), .B1(new_n497), .B2(new_n282), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n497), .A2(new_n282), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n327), .B1(new_n500), .B2(new_n495), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n486), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT18), .ZN(new_n505));
  INV_X1    g0305(.A(new_n479), .ZN(new_n506));
  INV_X1    g0306(.A(new_n472), .ZN(new_n507));
  AOI21_X1  g0307(.A(G20), .B1(new_n259), .B2(new_n261), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(KEYINPUT7), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(G68), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n303), .B(new_n484), .C1(new_n510), .C2(KEYINPUT16), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n502), .B1(new_n511), .B2(new_n469), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT18), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n387), .A2(new_n494), .A3(new_n417), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n493), .A2(new_n498), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n323), .B1(new_n500), .B2(new_n495), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n469), .B(new_n519), .C1(new_n480), .C2(new_n485), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT17), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT17), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n511), .A2(new_n522), .A3(new_n469), .A4(new_n519), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n521), .A2(KEYINPUT80), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n515), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n424), .A2(new_n465), .A3(new_n467), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n254), .A2(G1698), .ZN(new_n531));
  OAI221_X1 g0331(.A(new_n531), .B1(G250), .B2(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G294), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n282), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G264), .B(new_n282), .C1(new_n285), .C2(new_n274), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT90), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n275), .A2(new_n269), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(KEYINPUT90), .A3(G264), .A4(new_n282), .ZN(new_n539));
  AOI221_X4 g0339(.A(new_n534), .B1(new_n280), .B2(new_n271), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G179), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n539), .ZN(new_n543));
  INV_X1    g0343(.A(new_n534), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n318), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n327), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n225), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT22), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT89), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT89), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n550), .A3(KEYINPUT22), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n208), .A2(KEYINPUT22), .A3(G20), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n549), .A2(new_n551), .B1(new_n262), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT23), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n225), .B2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n391), .A2(KEYINPUT23), .A3(G20), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n555), .A2(new_n556), .B1(new_n354), .B2(G116), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT24), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n551), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n550), .B1(new_n547), .B2(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(new_n552), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n560), .A2(new_n561), .B1(new_n390), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n557), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n301), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n360), .A2(KEYINPUT25), .A3(new_n391), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT25), .B1(new_n360), .B2(new_n391), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n301), .A2(new_n295), .A3(new_n293), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n568), .A2(new_n569), .B1(new_n570), .B2(new_n391), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n542), .B(new_n546), .C1(new_n566), .C2(new_n571), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n553), .A2(KEYINPUT24), .A3(new_n558), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n564), .B1(new_n563), .B2(new_n557), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n303), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n543), .A2(new_n417), .A3(new_n318), .A4(new_n544), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n540), .B2(G200), .ZN(new_n577));
  INV_X1    g0377(.A(new_n571), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n570), .A2(new_n307), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT82), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n295), .B2(G97), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n360), .A2(KEYINPUT82), .A3(new_n307), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  AND2_X1   g0386(.A1(G97), .A2(G107), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g0390(.A1(KEYINPUT6), .A2(G97), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(G107), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n391), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(G97), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G20), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n355), .A2(G77), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(G107), .B2(new_n509), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n585), .B1(new_n598), .B2(new_n301), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT83), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n252), .A2(G244), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n249), .B2(new_n250), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n602), .B2(KEYINPUT4), .ZN(new_n603));
  OAI211_X1 g0403(.A(G244), .B(new_n252), .C1(new_n257), .C2(new_n258), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT4), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(KEYINPUT83), .A3(new_n605), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n601), .A2(new_n605), .B1(new_n209), .B2(new_n252), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n259), .A3(new_n261), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n603), .A2(new_n306), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n265), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n280), .A2(new_n271), .B1(new_n288), .B2(G257), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n327), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n381), .A3(new_n611), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n599), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n602), .A2(new_n600), .A3(KEYINPUT4), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT83), .B1(new_n604), .B2(new_n605), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n608), .A2(new_n306), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n282), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n288), .A2(G257), .ZN(new_n621));
  INV_X1    g0421(.A(new_n271), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n272), .A2(new_n275), .A3(new_n279), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(G200), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n594), .A2(G20), .B1(G77), .B2(new_n355), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n390), .A2(new_n225), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n472), .B1(new_n627), .B2(new_n471), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n628), .B2(new_n391), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n303), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n610), .A2(G190), .A3(new_n611), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n625), .A2(new_n630), .A3(new_n585), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n273), .A2(new_n276), .A3(G45), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n209), .B1(new_n341), .B2(G1), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n282), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n248), .A2(new_n309), .ZN(new_n636));
  NAND2_X1  g0436(.A1(G244), .A2(G1698), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n215), .B2(G1698), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n636), .B1(new_n251), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n635), .B1(new_n639), .B2(new_n282), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n399), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n327), .B2(new_n640), .ZN(new_n642));
  NOR3_X1   g0442(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT86), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(KEYINPUT19), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT19), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(KEYINPUT86), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n430), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n643), .B1(new_n648), .B2(new_n225), .ZN(new_n649));
  XNOR2_X1  g0449(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n225), .A2(G33), .A3(G97), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n225), .B(G68), .C1(new_n257), .C2(new_n258), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n303), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n315), .A2(new_n412), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n570), .A2(new_n412), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n642), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n215), .A2(G1698), .ZN(new_n661));
  AND2_X1   g0461(.A1(G244), .A2(G1698), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n257), .B2(new_n258), .ZN(new_n663));
  INV_X1    g0463(.A(new_n636), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n282), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n635), .ZN(new_n666));
  OAI21_X1  g0466(.A(G200), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n570), .A2(new_n208), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n655), .A2(new_n667), .A3(new_n656), .A4(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n640), .B2(G200), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(KEYINPUT87), .A3(new_n656), .A4(new_n655), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n640), .A2(new_n417), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n615), .A2(new_n632), .A3(new_n660), .A4(new_n677), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n334), .A2(new_n530), .A3(new_n580), .A4(new_n678), .ZN(G372));
  INV_X1    g0479(.A(new_n385), .ZN(new_n680));
  INV_X1    g0480(.A(new_n377), .ZN(new_n681));
  AOI211_X1 g0481(.A(KEYINPUT18), .B(new_n502), .C1(new_n511), .C2(new_n469), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n513), .B1(new_n486), .B2(new_n503), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n416), .B1(new_n464), .B2(new_n463), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n451), .B2(new_n462), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n521), .A2(KEYINPUT80), .A3(new_n523), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT80), .B1(new_n521), .B2(new_n523), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n684), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n681), .B1(new_n690), .B2(KEYINPUT94), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT94), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n692), .B(new_n684), .C1(new_n686), .C2(new_n689), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n680), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n615), .A2(new_n632), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  INV_X1    g0496(.A(new_n670), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n697), .A2(new_n676), .B1(new_n642), .B2(new_n659), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n579), .A4(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n615), .A2(new_n632), .A3(new_n698), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT91), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n317), .A2(new_n330), .A3(new_n541), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n328), .A2(new_n330), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT21), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n572), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n699), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n610), .A2(new_n381), .A3(new_n611), .ZN(new_n711));
  AOI21_X1  g0511(.A(G169), .B1(new_n610), .B2(new_n611), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n677), .A3(new_n599), .A4(new_n660), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT26), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n659), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n640), .A2(new_n327), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n399), .B2(new_n640), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n717), .A2(new_n719), .B1(new_n670), .B2(new_n675), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n715), .B1(new_n615), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT92), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n717), .A2(new_n719), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n674), .A2(new_n676), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n672), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n599), .A2(new_n614), .A3(new_n613), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(KEYINPUT93), .A3(KEYINPUT26), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n728), .B(new_n715), .C1(new_n615), .C2(new_n720), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n716), .A2(new_n722), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n709), .A2(new_n730), .A3(new_n660), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n530), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n694), .A2(new_n732), .ZN(G369));
  OAI21_X1  g0533(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n273), .A2(new_n225), .A3(G13), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT95), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT27), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(G213), .ZN(new_n740));
  INV_X1    g0540(.A(G343), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n317), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n333), .B2(new_n744), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n742), .B1(new_n566), .B2(new_n571), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n580), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n572), .B2(new_n743), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n572), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n743), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n707), .A2(new_n742), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n580), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(G399));
  INV_X1    g0557(.A(new_n220), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G41), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n643), .A2(new_n309), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n759), .A2(new_n273), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n229), .B2(new_n759), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT28), .Z(new_n763));
  INV_X1    g0563(.A(KEYINPUT29), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n731), .A2(new_n764), .A3(new_n743), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n579), .A2(new_n615), .A3(new_n632), .A4(new_n698), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n707), .B2(new_n572), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT26), .B1(new_n615), .B2(new_n720), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n768), .B(new_n660), .C1(new_n714), .C2(KEYINPUT26), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n743), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT29), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT30), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n281), .A2(new_n291), .A3(new_n610), .A4(new_n611), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n640), .A2(new_n541), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n543), .A2(new_n775), .A3(new_n544), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n776), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n624), .B1(new_n265), .B2(new_n609), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n778), .A2(new_n322), .A3(new_n779), .A4(KEYINPUT30), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n640), .A2(new_n381), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n612), .A2(new_n330), .A3(new_n545), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n777), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n783), .A2(KEYINPUT31), .A3(new_n742), .ZN(new_n784));
  AOI21_X1  g0584(.A(KEYINPUT31), .B1(new_n783), .B2(new_n742), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n334), .A2(new_n580), .A3(new_n678), .A4(new_n743), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G330), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n772), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT96), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT96), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n772), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n763), .B1(new_n794), .B2(G1), .ZN(G364));
  INV_X1    g0595(.A(new_n759), .ZN(new_n796));
  INV_X1    g0596(.A(G13), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G45), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(G1), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n758), .A2(new_n251), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G45), .B2(new_n228), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n242), .B2(G45), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n262), .A2(G355), .A3(new_n220), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G116), .B2(new_n220), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n403), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n224), .B1(G20), .B2(new_n327), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n801), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n381), .A2(new_n225), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n417), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(G190), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT33), .B(G317), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G326), .A2(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n225), .A2(G190), .A3(G200), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n381), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n225), .A2(G179), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n823), .A2(new_n417), .A3(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n822), .A2(G311), .B1(new_n825), .B2(G283), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n823), .A2(G190), .A3(G200), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n390), .B1(new_n263), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n417), .A2(G200), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n814), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n828), .B1(new_n831), .B2(G322), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n821), .A2(G179), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n829), .A2(new_n541), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n833), .A2(G329), .B1(new_n835), .B2(G294), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n819), .A2(new_n826), .A3(new_n832), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(G159), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT32), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G58), .B2(new_n831), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n816), .A2(G50), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n390), .B1(new_n822), .B2(G77), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n827), .A2(new_n208), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G107), .B2(new_n825), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n835), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n307), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n817), .B2(G68), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n837), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n813), .B1(new_n850), .B2(new_n810), .ZN(new_n851));
  INV_X1    g0651(.A(new_n809), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n746), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n747), .A2(new_n800), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n746), .A2(G330), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(G396));
  INV_X1    g0656(.A(KEYINPUT100), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n422), .A2(new_n743), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n731), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n857), .B1(new_n731), .B2(new_n858), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n731), .A2(new_n743), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n742), .B1(new_n415), .B2(new_n406), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n421), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n416), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n416), .A2(new_n742), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n859), .A2(new_n860), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n801), .B1(new_n868), .B2(new_n789), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n789), .B2(new_n868), .ZN(new_n870));
  INV_X1    g0670(.A(new_n810), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n262), .B(new_n847), .C1(new_n831), .C2(G294), .ZN(new_n872));
  INV_X1    g0672(.A(new_n833), .ZN(new_n873));
  INV_X1    g0673(.A(G311), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n873), .A2(new_n874), .B1(new_n827), .B2(new_n391), .ZN(new_n875));
  INV_X1    g0675(.A(new_n822), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n876), .A2(new_n309), .B1(new_n208), .B2(new_n824), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G283), .A2(new_n817), .B1(new_n816), .B2(G303), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n872), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n481), .B1(new_n833), .B2(G132), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n363), .A2(new_n827), .B1(new_n824), .B2(new_n214), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G58), .B2(new_n835), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n831), .A2(G143), .B1(G159), .B2(new_n822), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n816), .A2(G137), .ZN(new_n885));
  INV_X1    g0685(.A(G150), .ZN(new_n886));
  INV_X1    g0686(.A(new_n817), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT34), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n881), .B(new_n883), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n880), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT99), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n871), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n810), .A2(new_n403), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n800), .B1(new_n202), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n895), .B(new_n897), .C1(new_n867), .C2(new_n808), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n870), .A2(new_n898), .ZN(G384));
  NOR2_X1   g0699(.A1(new_n798), .A2(new_n273), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  INV_X1    g0701(.A(new_n865), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n731), .A2(new_n858), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT100), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n731), .A2(new_n857), .A3(new_n858), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n462), .A2(new_n742), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n448), .B2(new_n450), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n465), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n901), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n865), .B1(new_n859), .B2(new_n860), .ZN(new_n911));
  INV_X1    g0711(.A(new_n446), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT14), .B1(new_n444), .B2(new_n445), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n912), .A2(new_n913), .B1(new_n541), .B2(new_n441), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n449), .A2(KEYINPUT77), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT77), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n444), .B2(new_n425), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n462), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n464), .A2(new_n463), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n907), .ZN(new_n921));
  INV_X1    g0721(.A(new_n908), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n911), .A2(KEYINPUT101), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n520), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n512), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT37), .ZN(new_n927));
  INV_X1    g0727(.A(new_n740), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT102), .B1(new_n486), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n486), .A2(KEYINPUT102), .A3(new_n928), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n926), .B(new_n927), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT16), .B1(new_n483), .B2(new_n479), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n469), .B1(new_n485), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n503), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n928), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n520), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT37), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n528), .B2(new_n935), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT38), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(new_n942));
  INV_X1    g0742(.A(new_n935), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(KEYINPUT38), .A3(new_n938), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n910), .A2(new_n924), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT39), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n930), .A2(new_n929), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n504), .A2(new_n520), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT37), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n684), .A2(new_n524), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n951), .A2(new_n931), .B1(new_n952), .B2(new_n949), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n945), .B1(new_n953), .B2(KEYINPUT38), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n948), .B1(KEYINPUT39), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n919), .A2(new_n742), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n955), .A2(new_n956), .B1(new_n515), .B2(new_n740), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n947), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n691), .A2(new_n693), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n385), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n529), .B1(new_n771), .B2(new_n765), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n958), .B(new_n962), .Z(new_n963));
  INV_X1    g0763(.A(G330), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n866), .B1(new_n786), .B2(new_n787), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(new_n923), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT40), .B1(new_n946), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n965), .A2(new_n923), .A3(KEYINPUT40), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n954), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n529), .B1(new_n787), .B2(new_n786), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n900), .B1(new_n963), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n963), .B2(new_n972), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n975), .A2(G116), .A3(new_n226), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT36), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n229), .A2(G77), .A3(new_n477), .A4(new_n475), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(G50), .B2(new_n214), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(G1), .A3(new_n797), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(G367));
  NAND3_X1  g0782(.A1(new_n655), .A2(new_n656), .A3(new_n669), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n742), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT103), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n720), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n723), .B2(new_n985), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n809), .ZN(new_n988));
  INV_X1    g0788(.A(new_n412), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n812), .B1(new_n758), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n238), .A2(new_n802), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n800), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT107), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n827), .B2(new_n309), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n817), .A2(G294), .B1(KEYINPUT46), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n816), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(KEYINPUT46), .B2(new_n994), .C1(new_n874), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n833), .A2(G317), .ZN(new_n998));
  INV_X1    g0798(.A(G283), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n998), .B1(new_n846), .B2(new_n391), .C1(new_n876), .C2(new_n999), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n481), .B1(new_n307), .B2(new_n824), .C1(new_n830), .C2(new_n263), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT108), .Z(new_n1003));
  OAI22_X1  g0803(.A1(new_n212), .A2(new_n827), .B1(new_n824), .B2(new_n202), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n846), .A2(new_n214), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(G50), .C2(new_n822), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n831), .A2(G150), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n390), .B1(new_n833), .B2(G137), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G143), .A2(new_n816), .B1(new_n817), .B2(G159), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1003), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT47), .Z(new_n1012));
  OAI211_X1 g0812(.A(new_n988), .B(new_n992), .C1(new_n1012), .C2(new_n871), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n799), .A2(G1), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n756), .B1(new_n751), .B2(new_n755), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(new_n747), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n791), .B2(new_n793), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n599), .A2(new_n742), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n695), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n713), .A2(new_n599), .A3(new_n742), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT104), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(KEYINPUT105), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n756), .A2(new_n754), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1025), .A2(KEYINPUT105), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT45), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n1031), .A2(new_n1034), .A3(new_n752), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n752), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1017), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT106), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT106), .B1(new_n1017), .B2(new_n1037), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n794), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n759), .B(KEYINPUT41), .Z(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1014), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1032), .A2(new_n756), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT42), .Z(new_n1047));
  NAND2_X1  g0847(.A1(new_n1024), .A2(new_n753), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n742), .B1(new_n1048), .B2(new_n615), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT43), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1047), .A2(new_n1049), .B1(new_n1050), .B2(new_n987), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n987), .A2(new_n1050), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1051), .B(new_n1052), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n752), .A2(new_n1032), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1013), .B1(new_n1045), .B2(new_n1056), .ZN(G387));
  INV_X1    g0857(.A(new_n1017), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n791), .A2(new_n793), .A3(new_n1016), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n759), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n817), .A2(new_n353), .B1(G68), .B2(new_n822), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT111), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n251), .B1(new_n824), .B2(new_n307), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n835), .A2(new_n989), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n202), .B2(new_n827), .C1(new_n873), .C2(new_n886), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G50), .C2(new_n831), .ZN(new_n1066));
  INV_X1    g0866(.A(G159), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1062), .B(new_n1066), .C1(new_n1067), .C2(new_n996), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G311), .A2(new_n817), .B1(new_n816), .B2(G322), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT112), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(KEYINPUT112), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n831), .A2(G317), .B1(G303), .B2(new_n822), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(G294), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n846), .A2(new_n999), .B1(new_n827), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n251), .B1(new_n833), .B2(G326), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n309), .C2(new_n824), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT49), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1068), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n810), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n802), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n352), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT50), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n353), .B2(new_n363), .ZN(new_n1088));
  AOI211_X1 g0888(.A(G45), .B(new_n760), .C1(G68), .C2(G77), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1086), .B(new_n1088), .C1(new_n1090), .C2(KEYINPUT109), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1090), .A2(KEYINPUT109), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1085), .B(new_n1093), .C1(G45), .C2(new_n235), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n262), .A2(new_n220), .A3(new_n760), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(G107), .B2(new_n220), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1094), .A2(KEYINPUT110), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n812), .ZN(new_n1098));
  OAI21_X1  g0898(.A(KEYINPUT110), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n800), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1084), .B(new_n1100), .C1(new_n751), .C2(new_n852), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1014), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1060), .B(new_n1101), .C1(new_n1102), .C2(new_n1016), .ZN(G393));
  INV_X1    g0903(.A(new_n812), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n307), .B2(new_n220), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n245), .A2(new_n1085), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n801), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n833), .A2(G143), .B1(new_n835), .B2(G77), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n214), .B2(new_n827), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n481), .B(new_n1109), .C1(G87), .C2(new_n825), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n817), .A2(G50), .B1(new_n353), .B2(new_n822), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1111), .A2(KEYINPUT113), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(KEYINPUT113), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n816), .A2(G150), .B1(new_n831), .B2(G159), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n816), .A2(G317), .B1(new_n831), .B2(G311), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n817), .A2(G303), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n262), .B1(G107), .B2(new_n825), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n833), .A2(G322), .B1(new_n835), .B2(G116), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n827), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n822), .A2(G294), .B1(new_n1122), .B2(G283), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1114), .A2(new_n1116), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1107), .B1(new_n1125), .B2(new_n810), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1024), .B2(new_n852), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1037), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n1102), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1038), .B(new_n1039), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n796), .B1(new_n1058), .B2(new_n1128), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G390));
  AOI221_X4 g0933(.A(new_n940), .B1(new_n931), .B2(new_n937), .C1(new_n942), .C2(new_n943), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n951), .A2(new_n931), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n952), .A2(new_n949), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT38), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1138), .A2(new_n956), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT114), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n909), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n923), .A2(KEYINPUT114), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n743), .B(new_n864), .C1(new_n767), .C2(new_n769), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n865), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1139), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n956), .B1(new_n911), .B2(new_n923), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n955), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n964), .B(new_n866), .C1(new_n786), .C2(new_n787), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n923), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1147), .C1(new_n1148), .C2(new_n955), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT115), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n529), .A2(new_n789), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n694), .B(new_n1157), .C1(new_n529), .C2(new_n772), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n788), .A2(G330), .A3(new_n867), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n909), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1151), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1145), .B1(new_n1150), .B2(new_n923), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1141), .A2(new_n1159), .A3(new_n1142), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n911), .A2(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1156), .B1(new_n1158), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT115), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1155), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1153), .A2(new_n1154), .A3(new_n1166), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n759), .A3(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n955), .A2(new_n808), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n896), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n801), .B1(new_n353), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G107), .A2(new_n817), .B1(new_n816), .B2(G283), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n262), .B(new_n843), .C1(new_n831), .C2(G116), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G68), .A2(new_n825), .B1(new_n835), .B2(G77), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n822), .A2(G97), .B1(new_n833), .B2(G294), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n833), .A2(G125), .B1(new_n825), .B2(G50), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n1067), .B2(new_n846), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G137), .B2(new_n817), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n886), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT53), .B1(new_n827), .B2(new_n886), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT54), .B(G143), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n390), .B1(new_n822), .B2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n816), .A2(G128), .B1(new_n831), .B2(G132), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT116), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1178), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1173), .B1(new_n1190), .B2(new_n810), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1171), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1155), .B2(new_n1102), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT117), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(KEYINPUT117), .B(new_n1192), .C1(new_n1155), .C2(new_n1102), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1170), .A2(new_n1195), .A3(new_n1196), .ZN(G378));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n377), .A2(new_n385), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1200), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n377), .A2(new_n385), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n378), .A2(new_n928), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1201), .A2(new_n378), .A3(new_n928), .A4(new_n1203), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n965), .A2(new_n923), .A3(KEYINPUT40), .ZN(new_n1209));
  OAI21_X1  g1009(.A(G330), .B1(new_n1138), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1210), .B2(new_n967), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT40), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT38), .B1(new_n944), .B2(new_n938), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1134), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n965), .A2(new_n923), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1212), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n964), .B1(new_n968), .B2(new_n954), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n958), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n947), .A2(new_n1220), .A3(new_n957), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1198), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n529), .A2(new_n789), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n960), .A2(new_n961), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1169), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1211), .A2(KEYINPUT119), .A3(new_n1219), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT119), .B1(new_n1211), .B2(new_n1219), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n958), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1223), .A2(new_n1232), .B1(new_n1169), .B2(new_n1226), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1228), .B(new_n759), .C1(new_n1233), .C2(KEYINPUT57), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1223), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1218), .A2(new_n403), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n801), .B1(G50), .B2(new_n1172), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1122), .A2(new_n1185), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT118), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n817), .A2(G132), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n822), .A2(G137), .B1(new_n835), .B2(G150), .ZN(new_n1241));
  INV_X1    g1041(.A(G128), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1240), .B(new_n1241), .C1(new_n1242), .C2(new_n830), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1239), .B(new_n1243), .C1(G125), .C2(new_n816), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT59), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n248), .B(new_n266), .C1(new_n824), .C2(new_n1067), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G124), .B2(new_n833), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n251), .A2(G41), .ZN(new_n1251));
  AOI211_X1 g1051(.A(G50), .B(new_n1251), .C1(new_n248), .C2(new_n266), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1251), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1253), .B(new_n1005), .C1(G107), .C2(new_n831), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n822), .A2(new_n989), .B1(new_n1122), .B2(G77), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n824), .A2(new_n212), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G283), .B2(new_n833), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G97), .A2(new_n817), .B1(new_n816), .B2(G116), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT58), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1252), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1250), .B(new_n1261), .C1(new_n1260), .C2(new_n1259), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1237), .B1(new_n1262), .B2(new_n810), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1235), .A2(new_n1014), .B1(new_n1236), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1234), .A2(new_n1264), .ZN(G375));
  NAND2_X1  g1065(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1167), .A2(new_n1044), .A3(new_n1165), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1161), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n906), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1014), .B(KEYINPUT120), .Z(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1143), .A2(new_n403), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT121), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n801), .B1(G68), .B2(new_n1172), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n816), .A2(G132), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT123), .Z(new_n1277));
  AOI22_X1  g1077(.A1(new_n817), .A2(new_n1185), .B1(new_n831), .B2(G137), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT124), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G159), .A2(new_n1122), .B1(new_n835), .B2(G50), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1281), .B1(new_n876), .B2(new_n886), .C1(new_n1242), .C2(new_n873), .ZN(new_n1282));
  OR3_X1    g1082(.A1(new_n1282), .A2(new_n481), .A3(new_n1256), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1064), .B1(new_n830), .B2(new_n999), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT122), .Z(new_n1285));
  OAI21_X1  g1085(.A(new_n390), .B1(new_n202), .B2(new_n824), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n873), .A2(new_n263), .B1(new_n827), .B2(new_n307), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1286), .B(new_n1287), .C1(G107), .C2(new_n822), .ZN(new_n1288));
  OAI221_X1 g1088(.A(new_n1288), .B1(new_n309), .B2(new_n887), .C1(new_n1076), .C2(new_n996), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1280), .A2(new_n1283), .B1(new_n1285), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1275), .B1(new_n1290), .B2(new_n810), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1272), .B1(new_n1274), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1267), .A2(new_n1294), .ZN(G381));
  OAI211_X1 g1095(.A(new_n1013), .B(new_n1132), .C1(new_n1045), .C2(new_n1056), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1193), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1170), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G384), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1267), .A2(new_n1294), .A3(new_n1300), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(new_n1299), .A2(new_n1301), .A3(G396), .A4(G393), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1235), .A2(new_n1014), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1236), .A2(new_n1263), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1235), .A2(new_n1227), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1198), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n796), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1305), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1297), .A2(new_n1302), .A3(new_n1309), .ZN(G407));
  INV_X1    g1110(.A(new_n1299), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n741), .A2(G213), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1309), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(G407), .A2(G213), .A3(new_n1314), .ZN(G409));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT60), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1226), .B2(new_n1270), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1226), .A2(new_n1270), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1158), .A2(new_n1164), .A3(KEYINPUT60), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n759), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1316), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1322), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1266), .B1(new_n1166), .B2(new_n1317), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(KEYINPUT126), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(G384), .B1(new_n1327), .B2(new_n1294), .ZN(new_n1328));
  AOI211_X1 g1128(.A(new_n1300), .B(new_n1293), .C1(new_n1323), .C2(new_n1326), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1234), .A2(G378), .A3(new_n1264), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n947), .A2(new_n1220), .A3(new_n957), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1220), .B1(new_n947), .B2(new_n957), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1271), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1304), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1235), .A2(new_n1227), .A3(new_n1044), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT125), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1335), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1235), .A2(new_n1227), .A3(KEYINPUT125), .A4(new_n1044), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1299), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1312), .B(new_n1330), .C1(new_n1331), .C2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(KEYINPUT62), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1313), .A2(G2897), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1328), .A2(new_n1329), .A3(new_n1345), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1320), .A2(new_n1322), .A3(new_n1316), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT126), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1294), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1300), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1327), .A2(G384), .A3(new_n1294), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1344), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1346), .A2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1227), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT119), .ZN(new_n1355));
  NOR3_X1   g1155(.A1(new_n1210), .A2(new_n967), .A3(new_n1208), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1355), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  AOI22_X1  g1158(.A1(new_n1358), .A2(new_n1229), .B1(new_n947), .B2(new_n957), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1044), .B1(new_n1359), .B2(new_n1332), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1337), .B1(new_n1354), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1335), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1361), .A2(new_n1339), .A3(new_n1362), .ZN(new_n1363));
  AOI22_X1  g1163(.A1(new_n1309), .A2(G378), .B1(new_n1363), .B2(new_n1311), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1353), .B1(new_n1364), .B2(new_n1313), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1311), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1234), .A2(G378), .A3(new_n1264), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT62), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1368), .A2(new_n1369), .A3(new_n1312), .A4(new_n1330), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1342), .A2(new_n1343), .A3(new_n1365), .A4(new_n1370), .ZN(new_n1371));
  XOR2_X1   g1171(.A(G393), .B(G396), .Z(new_n1372));
  AOI21_X1  g1172(.A(new_n1043), .B1(new_n1130), .B2(new_n794), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1055), .B1(new_n1373), .B2(new_n1014), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1132), .B1(new_n1374), .B2(new_n1013), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1296), .A2(KEYINPUT127), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1372), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(G387), .A2(G390), .ZN(new_n1378));
  INV_X1    g1178(.A(new_n1372), .ZN(new_n1379));
  NAND4_X1  g1179(.A1(new_n1378), .A2(new_n1379), .A3(KEYINPUT127), .A4(new_n1296), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1377), .A2(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1371), .A2(new_n1381), .ZN(new_n1382));
  AND2_X1   g1182(.A1(new_n1377), .A2(new_n1380), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1368), .A2(new_n1312), .ZN(new_n1384));
  AOI21_X1  g1184(.A(KEYINPUT61), .B1(new_n1384), .B2(new_n1353), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT63), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1341), .A2(new_n1386), .ZN(new_n1387));
  NAND4_X1  g1187(.A1(new_n1368), .A2(KEYINPUT63), .A3(new_n1312), .A4(new_n1330), .ZN(new_n1388));
  NAND4_X1  g1188(.A1(new_n1383), .A2(new_n1385), .A3(new_n1387), .A4(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1382), .A2(new_n1389), .ZN(G405));
  NAND2_X1  g1190(.A1(G375), .A2(new_n1311), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1391), .A2(new_n1367), .ZN(new_n1392));
  OR2_X1    g1192(.A1(new_n1392), .A2(new_n1330), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1392), .A2(new_n1330), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1393), .A2(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1395), .A2(new_n1381), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1383), .A2(new_n1394), .A3(new_n1393), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1396), .A2(new_n1397), .ZN(G402));
endmodule


