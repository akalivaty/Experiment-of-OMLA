//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  AND4_X1   g007(.A1(KEYINPUT25), .A2(new_n205), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT24), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(G183gat), .A3(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n215));
  OR3_X1    g014(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT67), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT65), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT23), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n221), .A2(new_n208), .A3(new_n224), .A4(new_n207), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n211), .A2(new_n213), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n220), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n217), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n219), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n227), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n237), .A2(KEYINPUT69), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n237), .A2(KEYINPUT69), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n222), .A2(KEYINPUT70), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT70), .B1(new_n222), .B2(new_n240), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n238), .B(new_n239), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT28), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n233), .A2(KEYINPUT68), .A3(new_n244), .A4(new_n227), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n236), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n232), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT29), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT78), .B(G218gat), .Z(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT77), .B(G211gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT22), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G197gat), .B(G204gat), .Z(new_n258));
  OAI211_X1 g057(.A(KEYINPUT79), .B(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(KEYINPUT79), .ZN(new_n260));
  INV_X1    g059(.A(new_n258), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT77), .B(G211gat), .Z(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT78), .B(G218gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n260), .B(new_n261), .C1(new_n264), .C2(KEYINPUT22), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n252), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n259), .A2(new_n265), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT80), .B(KEYINPUT29), .Z(new_n269));
  AOI21_X1  g068(.A(new_n248), .B1(new_n247), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n249), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G64gat), .ZN(new_n273));
  INV_X1    g072(.A(G92gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n267), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(KEYINPUT81), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n275), .B1(new_n267), .B2(new_n271), .ZN(new_n283));
  INV_X1    g082(.A(new_n276), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n286), .A2(KEYINPUT35), .ZN(new_n287));
  XNOR2_X1  g086(.A(G141gat), .B(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291));
  OR2_X1    g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(KEYINPUT82), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G155gat), .B(G162gat), .Z(new_n296));
  INV_X1    g095(.A(new_n288), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n291), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n298), .B2(new_n299), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n295), .A2(new_n296), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n302), .A2(KEYINPUT83), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT83), .B1(new_n302), .B2(new_n303), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n295), .A2(new_n296), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G127gat), .B(G134gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(G120gat), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n318), .C1(G113gat), .C2(new_n317), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n312), .A2(new_n313), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n311), .B1(KEYINPUT1), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n309), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n322), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n302), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT4), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n331), .A3(new_n302), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n307), .A2(new_n308), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n325), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n338), .B1(new_n341), .B2(new_n335), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n306), .A2(new_n326), .B1(new_n330), .B2(new_n332), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n337), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n346));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G57gat), .ZN(new_n349));
  INV_X1    g148(.A(G85gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT90), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(new_n351), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n346), .B1(new_n345), .B2(new_n351), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT88), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n344), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n351), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n362), .A2(new_n354), .A3(new_n363), .A4(new_n346), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n353), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n236), .A2(new_n243), .A3(new_n245), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n209), .A2(new_n217), .A3(new_n230), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n230), .B1(new_n209), .B2(new_n217), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n367), .B1(new_n370), .B2(new_n229), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT74), .B1(new_n371), .B2(new_n328), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n247), .A2(new_n373), .A3(new_n325), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n232), .A2(new_n328), .A3(new_n246), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n232), .A2(new_n328), .A3(KEYINPUT73), .A4(new_n246), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n372), .A2(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT32), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  XOR2_X1   g182(.A(G15gat), .B(G43gat), .Z(new_n384));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n386), .ZN(new_n388));
  OAI221_X1 g187(.A(KEYINPUT32), .B1(new_n382), .B2(new_n388), .C1(new_n379), .C2(new_n380), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n374), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n377), .A2(new_n378), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n380), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n397));
  INV_X1    g196(.A(new_n269), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n302), .B2(new_n303), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n399), .B2(new_n266), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n309), .A2(new_n269), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(new_n268), .A3(KEYINPUT85), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n259), .B2(new_n265), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n339), .B1(new_n403), .B2(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n400), .A2(new_n402), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n405), .B(KEYINPUT84), .Z(new_n408));
  NOR2_X1   g207(.A1(new_n399), .A2(new_n266), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n254), .B(new_n261), .C1(new_n264), .C2(KEYINPUT22), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n269), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n302), .B1(new_n412), .B2(new_n303), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n408), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT86), .B1(new_n415), .B2(G22gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT31), .ZN(new_n418));
  INV_X1    g217(.A(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n407), .B2(new_n414), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n407), .A2(new_n422), .A3(new_n414), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n416), .A2(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n423), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n422), .A3(new_n414), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(KEYINPUT86), .A3(new_n427), .A4(new_n420), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n394), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n393), .B(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n387), .A3(new_n389), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n396), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n287), .A2(new_n366), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(KEYINPUT91), .ZN(new_n435));
  INV_X1    g234(.A(new_n356), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n352), .B1(new_n436), .B2(new_n354), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n286), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT91), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n396), .A2(new_n429), .A3(new_n439), .A4(new_n432), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(KEYINPUT92), .A3(KEYINPUT35), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n434), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n267), .A2(new_n447), .A3(new_n271), .ZN(new_n448));
  INV_X1    g247(.A(new_n275), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT38), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n252), .A2(new_n268), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n266), .B1(new_n249), .B2(new_n270), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(KEYINPUT37), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n448), .A2(new_n455), .A3(new_n452), .A4(new_n449), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT89), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n267), .A2(new_n271), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n449), .A3(new_n448), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n284), .B1(new_n462), .B2(KEYINPUT38), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n365), .A2(new_n353), .A3(new_n459), .A4(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n283), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n277), .B2(new_n276), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n280), .B2(new_n281), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n329), .A2(new_n334), .A3(new_n340), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT39), .B(new_n468), .C1(new_n343), .C2(new_n334), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n327), .A2(new_n333), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n335), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n472), .A3(new_n351), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT40), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n469), .A2(new_n472), .A3(KEYINPUT40), .A4(new_n351), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n362), .A3(new_n476), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n467), .A2(KEYINPUT87), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n479));
  INV_X1    g278(.A(new_n477), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n286), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n464), .B(new_n429), .C1(new_n478), .C2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n429), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n286), .B2(new_n437), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n396), .A2(new_n432), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT36), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT36), .B1(new_n396), .B2(new_n432), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(KEYINPUT76), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(KEYINPUT76), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n482), .B(new_n484), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n202), .B1(new_n446), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n434), .ZN(new_n494));
  INV_X1    g293(.A(new_n445), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT92), .B1(new_n441), .B2(KEYINPUT35), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT93), .A3(new_n491), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT98), .ZN(new_n500));
  INV_X1    g299(.A(G43gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n419), .ZN(new_n502));
  NAND2_X1  g301(.A1(G43gat), .A2(G50gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OR3_X1    g307(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT94), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n506), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n502), .A2(new_n516), .A3(new_n503), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n505), .A2(new_n515), .A3(new_n512), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(KEYINPUT17), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  INV_X1    g319(.A(new_n518), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(new_n513), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n523), .A2(G1gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT16), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT95), .B(G8gat), .Z(new_n529));
  NAND4_X1  g328(.A1(new_n524), .A2(new_n525), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(G1gat), .B2(new_n523), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n531), .A2(KEYINPUT96), .B1(new_n532), .B2(G8gat), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n519), .A2(new_n522), .A3(new_n530), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(KEYINPUT96), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(G8gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n514), .A2(new_n518), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n541), .A2(KEYINPUT97), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT97), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n540), .B(KEYINPUT13), .Z(new_n545));
  NOR2_X1   g344(.A1(new_n537), .A2(new_n538), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n533), .A2(new_n530), .B1(new_n514), .B2(new_n518), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n534), .A2(new_n539), .A3(KEYINPUT18), .A4(new_n540), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n543), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G113gat), .B(G141gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT11), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G169gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G197gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n553), .B(new_n203), .ZN(new_n556));
  INV_X1    g355(.A(G197gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n555), .A2(new_n558), .A3(KEYINPUT12), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT12), .B1(new_n555), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n500), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n541), .A2(new_n542), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n548), .A2(new_n549), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(KEYINPUT98), .B(new_n563), .C1(new_n568), .C2(new_n543), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n561), .A2(new_n567), .A3(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  INV_X1    g372(.A(G71gat), .ZN(new_n574));
  INV_X1    g373(.A(G78gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n578), .B(new_n579), .C1(KEYINPUT99), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(KEYINPUT99), .ZN(new_n582));
  XNOR2_X1  g381(.A(G71gat), .B(G78gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n580), .A2(new_n573), .ZN(new_n585));
  OAI22_X1  g384(.A1(new_n581), .A2(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n530), .B(new_n533), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n226), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT101), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n586), .A2(new_n587), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(G211gat), .Z(new_n598));
  OR2_X1    g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n598), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  INV_X1    g403(.A(KEYINPUT103), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n274), .ZN(new_n606));
  NAND2_X1  g405(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n350), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT104), .ZN(new_n609));
  INV_X1    g408(.A(G99gat), .ZN(new_n610));
  INV_X1    g409(.A(G106gat), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT8), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n608), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n616), .B(new_n604), .C1(new_n613), .C2(new_n614), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(KEYINPUT105), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT105), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n615), .A2(new_n621), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n538), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n519), .A2(new_n522), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n624), .B(new_n625), .C1(new_n623), .C2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n627), .A2(new_n628), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n630), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n630), .B2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n601), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G176gat), .ZN(new_n641));
  INV_X1    g440(.A(G204gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT107), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n620), .A2(new_n586), .A3(new_n622), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT106), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n620), .A2(new_n649), .A3(new_n586), .A4(new_n622), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  INV_X1    g451(.A(new_n618), .ZN(new_n653));
  INV_X1    g452(.A(new_n619), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n653), .A2(new_n654), .A3(new_n586), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n586), .A2(new_n652), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n622), .B2(new_n620), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n646), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n655), .B1(new_n648), .B2(new_n650), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n645), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n644), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n644), .ZN(new_n665));
  AOI211_X1 g464(.A(KEYINPUT10), .B(new_n655), .C1(new_n648), .C2(new_n650), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n645), .B1(new_n666), .B2(new_n659), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n639), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT108), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n499), .A2(new_n572), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n352), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n355), .B2(new_n356), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n526), .ZN(G1324gat));
  INV_X1    g476(.A(new_n673), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n286), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n678), .A2(KEYINPUT42), .A3(new_n286), .A4(new_n679), .ZN(new_n683));
  OAI21_X1  g482(.A(G8gat), .B1(new_n673), .B2(new_n467), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(G1325gat));
  NOR2_X1   g484(.A1(new_n489), .A2(new_n490), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n673), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n485), .A2(G15gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n673), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n688), .B(KEYINPUT109), .C1(new_n673), .C2(new_n690), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n673), .A2(new_n429), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT110), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n696), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n638), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n493), .A2(new_n498), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n484), .A2(KEYINPUT111), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n484), .A2(KEYINPUT111), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n482), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n686), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n638), .B1(new_n446), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n701), .ZN(new_n709));
  INV_X1    g508(.A(new_n601), .ZN(new_n710));
  INV_X1    g509(.A(new_n572), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(new_n669), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n703), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT112), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n703), .A2(new_n709), .A3(new_n715), .A4(new_n712), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n437), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G29gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n710), .A2(new_n669), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n638), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G29gat), .A3(new_n675), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n499), .A2(new_n572), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT45), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n714), .A2(new_n286), .A3(new_n716), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G36gat), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n720), .A2(G36gat), .A3(new_n467), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n499), .A2(new_n572), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT113), .B(KEYINPUT46), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(G1329gat));
  OAI21_X1  g530(.A(G43gat), .B1(new_n713), .B2(new_n687), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n499), .A2(new_n572), .A3(new_n638), .A4(new_n719), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n486), .A2(new_n501), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n732), .B(KEYINPUT47), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n714), .A2(new_n686), .A3(new_n716), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n738), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g538(.A(G50gat), .B1(new_n713), .B2(new_n429), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n483), .A2(new_n419), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n740), .B(KEYINPUT48), .C1(new_n733), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n733), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n714), .A2(new_n483), .A3(new_n716), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G50gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n745), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n446), .A2(new_n707), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n639), .A2(new_n711), .A3(new_n669), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n437), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g550(.A1(new_n747), .A2(new_n467), .A3(new_n748), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  AND2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n752), .B2(new_n753), .ZN(G1333gat));
  NOR2_X1   g555(.A1(new_n687), .A2(new_n574), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(KEYINPUT114), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(KEYINPUT114), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n485), .B(KEYINPUT115), .Z(new_n761));
  AND2_X1   g560(.A1(new_n749), .A2(new_n761), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n759), .A2(new_n760), .B1(G71gat), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n483), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n710), .A2(new_n572), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n638), .B(new_n767), .C1(new_n446), .C2(new_n707), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n350), .A3(new_n437), .A4(new_n669), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n710), .A2(new_n670), .A3(new_n572), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n703), .A2(new_n709), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n437), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(new_n350), .ZN(G1336gat));
  NAND4_X1  g574(.A1(new_n770), .A2(new_n274), .A3(new_n286), .A4(new_n669), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n703), .A2(new_n709), .A3(new_n286), .A4(new_n772), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n606), .A2(new_n607), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n768), .A2(new_n782), .A3(new_n769), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n467), .A2(new_n670), .A3(G92gat), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n783), .B(new_n784), .C1(new_n770), .C2(new_n782), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n780), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n786), .B2(new_n777), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n486), .A3(new_n669), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n687), .A2(new_n610), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n788), .A2(new_n610), .B1(new_n773), .B2(new_n789), .ZN(G1338gat));
  NOR3_X1   g589(.A1(new_n670), .A2(G106gat), .A3(new_n429), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n783), .B(new_n791), .C1(new_n770), .C2(new_n782), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n703), .A2(new_n709), .A3(new_n483), .A4(new_n772), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT53), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT53), .B1(new_n770), .B2(new_n791), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1339gat));
  AOI21_X1  g598(.A(new_n659), .B1(new_n662), .B2(new_n652), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n646), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT117), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n657), .A2(new_n803), .A3(new_n646), .A4(new_n660), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n667), .A4(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n643), .B1(new_n661), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT118), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n570), .A2(new_n571), .B1(new_n667), .B2(new_n665), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n667), .A2(new_n804), .A3(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n803), .B1(new_n800), .B2(new_n646), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n807), .B(KEYINPUT55), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n809), .A2(new_n814), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n555), .A2(new_n558), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n546), .A2(new_n547), .A3(new_n545), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n540), .B1(new_n534), .B2(new_n539), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n571), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n669), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n638), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n813), .A2(new_n638), .A3(new_n668), .A4(new_n825), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n809), .A3(new_n819), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n601), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n639), .A2(new_n711), .A3(new_n670), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n483), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n286), .A2(new_n675), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n486), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n836), .A2(new_n315), .A3(new_n711), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n675), .B1(new_n832), .B2(new_n833), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n435), .A2(new_n440), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n467), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n572), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n837), .B1(new_n842), .B2(new_n315), .ZN(G1340gat));
  NOR3_X1   g642(.A1(new_n836), .A2(new_n317), .A3(new_n670), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n669), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n317), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n841), .A2(new_n847), .A3(new_n710), .ZN(new_n848));
  OAI21_X1  g647(.A(G127gat), .B1(new_n836), .B2(new_n601), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n700), .A2(new_n286), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n840), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n836), .B2(new_n700), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(G1343gat));
  NAND2_X1  g656(.A1(new_n687), .A2(new_n835), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n429), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n833), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n817), .A2(new_n813), .A3(new_n810), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n638), .B1(new_n864), .B2(new_n826), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n830), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT119), .B(new_n638), .C1(new_n864), .C2(new_n826), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n601), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n863), .B1(new_n869), .B2(KEYINPUT120), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n601), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n862), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n832), .A2(new_n833), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT57), .B1(new_n874), .B2(new_n483), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n859), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G141gat), .B1(new_n876), .B2(new_n711), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n686), .A2(new_n429), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n838), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n711), .A2(G141gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n467), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT122), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n877), .A2(new_n886), .A3(new_n883), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1344gat));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n483), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n831), .A2(new_n865), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n710), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n672), .A2(new_n711), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n860), .B(new_n483), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n669), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G148gat), .B1(new_n897), .B2(new_n858), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT59), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n669), .B(new_n859), .C1(new_n873), .C2(new_n875), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901));
  INV_X1    g700(.A(G148gat), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(KEYINPUT59), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n879), .A2(new_n467), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n902), .A3(new_n669), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1345gat));
  NOR3_X1   g708(.A1(new_n876), .A2(new_n298), .A3(new_n601), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n710), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  AOI21_X1  g711(.A(G155gat), .B1(new_n911), .B2(KEYINPUT124), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1346gat));
  OAI211_X1 g713(.A(new_n638), .B(new_n859), .C1(new_n873), .C2(new_n875), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n299), .B1(new_n915), .B2(KEYINPUT125), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(KEYINPUT125), .B2(new_n915), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n879), .A2(new_n299), .A3(new_n852), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1347gat));
  AOI21_X1  g718(.A(new_n437), .B1(new_n832), .B2(new_n833), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n839), .A2(new_n286), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n203), .A3(new_n572), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n467), .A2(new_n437), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n834), .A2(new_n761), .A3(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n711), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n927), .B2(new_n670), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n923), .A2(new_n204), .A3(new_n669), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1349gat));
  AOI21_X1  g733(.A(new_n226), .B1(new_n926), .B2(new_n710), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n710), .A2(new_n233), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n923), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n227), .A3(new_n638), .ZN(new_n940));
  OAI21_X1  g739(.A(G190gat), .B1(new_n927), .B2(new_n700), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n878), .A2(new_n286), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n920), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n557), .B1(new_n947), .B2(new_n711), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n892), .A2(new_n687), .A3(new_n896), .A4(new_n925), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n572), .A2(G197gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n947), .A2(G204gat), .A3(new_n670), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n687), .A2(new_n925), .ZN(new_n955));
  OAI21_X1  g754(.A(G204gat), .B1(new_n897), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  NAND4_X1  g756(.A1(new_n920), .A2(new_n946), .A3(new_n262), .A4(new_n710), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n949), .A2(new_n601), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n960));
  OAI211_X1 g759(.A(KEYINPUT63), .B(G211gat), .C1(new_n949), .C2(new_n601), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n960), .B2(new_n962), .ZN(G1354gat));
  NAND2_X1  g762(.A1(new_n638), .A2(new_n255), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n700), .ZN(new_n965));
  OAI22_X1  g764(.A1(new_n949), .A2(new_n964), .B1(G218gat), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(G1355gat));
endmodule


