//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G197gat), .B(G204gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT75), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n209), .B2(KEYINPUT22), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n212));
  OAI21_X1  g011(.A(G211gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(KEYINPUT75), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n204), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n203), .B1(new_n216), .B2(KEYINPUT76), .ZN(new_n217));
  INV_X1    g016(.A(new_n204), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n213), .A2(KEYINPUT75), .A3(new_n214), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT75), .B1(new_n213), .B2(new_n214), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT76), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n202), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT27), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT68), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT69), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OR3_X1    g036(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n237), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n231), .A2(KEYINPUT69), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT28), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT69), .B1(new_n231), .B2(KEYINPUT68), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n235), .B(new_n245), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n230), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(new_n237), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n255), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n238), .A2(KEYINPUT23), .A3(new_n240), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n243), .A2(KEYINPUT23), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT25), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267));
  OR2_X1    g066(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(KEYINPUT23), .A3(new_n262), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n236), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(new_n253), .A3(new_n250), .ZN(new_n273));
  AND4_X1   g072(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(new_n264), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n249), .A2(new_n266), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT78), .B1(new_n281), .B2(new_n277), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n264), .B(new_n259), .C1(new_n252), .C2(new_n257), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n274), .B1(new_n283), .B2(KEYINPUT25), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT29), .B1(new_n284), .B2(new_n249), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT78), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n285), .A2(new_n286), .A3(new_n278), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n225), .B(new_n279), .C1(new_n282), .C2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n278), .B1(new_n276), .B2(new_n280), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n277), .B1(new_n284), .B2(new_n249), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n224), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n279), .B1(new_n278), .B2(new_n285), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n289), .B1(new_n294), .B2(new_n224), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n288), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n224), .B1(new_n290), .B2(new_n291), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT77), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n292), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n304), .A2(KEYINPUT30), .A3(new_n288), .A4(new_n299), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n281), .A2(KEYINPUT78), .A3(new_n277), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n286), .B1(new_n285), .B2(new_n278), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n291), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n303), .A2(new_n292), .B1(new_n309), .B2(new_n225), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT30), .B1(new_n310), .B2(new_n299), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT87), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT34), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(KEYINPUT1), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G113gat), .B(G120gat), .Z(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n315), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n284), .A2(new_n323), .A3(new_n249), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n314), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n322), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n276), .A2(KEYINPUT70), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G227gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n313), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  AOI211_X1 g132(.A(KEYINPUT34), .B(new_n331), .C1(new_n325), .C2(new_n327), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n325), .A2(new_n331), .A3(new_n327), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G15gat), .B(G43gat), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT71), .ZN(new_n341));
  XOR2_X1   g140(.A(G71gat), .B(G99gat), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT72), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n341), .B(new_n343), .Z(new_n344));
  NAND3_X1  g143(.A1(new_n337), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n344), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n336), .B(KEYINPUT32), .C1(new_n338), .C2(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n335), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n333), .ZN(new_n349));
  INV_X1    g148(.A(new_n334), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n345), .A2(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n304), .A2(new_n288), .A3(new_n299), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n301), .A4(new_n305), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  NAND2_X1  g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(KEYINPUT2), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n359), .A3(KEYINPUT2), .ZN(new_n363));
  INV_X1    g162(.A(G155gat), .ZN(new_n364));
  INV_X1    g163(.A(G162gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n360), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT80), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n369), .A3(new_n360), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n362), .A2(new_n363), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n358), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n360), .A2(KEYINPUT2), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n372), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n371), .A2(new_n322), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n368), .A2(new_n370), .ZN(new_n376));
  INV_X1    g175(.A(new_n361), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n377), .A3(new_n363), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n358), .B1(new_n360), .B2(new_n366), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n373), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n379), .A2(new_n381), .B1(new_n321), .B2(new_n318), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT5), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n376), .A2(new_n378), .B1(new_n380), .B2(new_n373), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(new_n371), .B2(new_n374), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n322), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n379), .A2(new_n381), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n322), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n326), .A2(new_n386), .A3(KEYINPUT4), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n390), .A2(new_n393), .A3(new_n384), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n393), .A2(new_n394), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(KEYINPUT5), .A3(new_n384), .A4(new_n390), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT0), .ZN(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405));
  INV_X1    g204(.A(new_n403), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT6), .A4(new_n406), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT35), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n312), .A2(new_n352), .A3(new_n357), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n217), .A2(new_n223), .A3(new_n280), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n217), .A2(new_n223), .A3(new_n414), .A4(new_n280), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n387), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n392), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n217), .A2(new_n223), .B1(new_n388), .B2(new_n280), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n221), .A2(new_n202), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n216), .A2(new_n203), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n280), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n386), .B1(new_n426), .B2(new_n387), .ZN(new_n427));
  INV_X1    g226(.A(G228gat), .ZN(new_n428));
  OAI22_X1  g227(.A1(new_n427), .A2(new_n418), .B1(new_n428), .B2(new_n330), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n422), .A2(KEYINPUT84), .A3(new_n423), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT3), .B1(new_n412), .B2(KEYINPUT83), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n386), .B1(new_n431), .B2(new_n415), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n423), .B(new_n429), .C1(new_n432), .C2(new_n420), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n420), .B1(new_n416), .B2(new_n392), .ZN(new_n436));
  INV_X1    g235(.A(new_n429), .ZN(new_n437));
  OAI21_X1  g236(.A(G22gat), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(G78gat), .B(G106gat), .Z(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT31), .B(G50gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n439), .A2(KEYINPUT85), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n422), .A2(new_n429), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n442), .B1(new_n448), .B2(G22gat), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n433), .A2(new_n450), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n411), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n439), .A2(KEYINPUT85), .A3(new_n442), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT85), .B1(new_n439), .B2(new_n442), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n408), .A2(new_n409), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n355), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n301), .B2(new_n305), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n301), .A2(new_n305), .A3(new_n460), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT82), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n306), .A2(KEYINPUT79), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n409), .A2(new_n408), .B1(new_n353), .B2(new_n354), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n345), .A2(new_n347), .ZN(new_n470));
  INV_X1    g269(.A(new_n335), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n335), .A2(new_n345), .A3(new_n347), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT73), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(KEYINPUT73), .B2(new_n472), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n457), .A2(new_n464), .A3(new_n469), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n454), .B1(new_n476), .B2(KEYINPUT35), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n453), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n445), .B2(new_n446), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT82), .B1(new_n462), .B2(new_n463), .ZN(new_n481));
  AND4_X1   g280(.A1(KEYINPUT82), .A2(new_n465), .A3(new_n463), .A4(new_n466), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n288), .B(new_n485), .C1(new_n293), .C2(new_n295), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT90), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT90), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n304), .A2(new_n488), .A3(new_n288), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n309), .A2(new_n224), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n294), .B2(new_n225), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT38), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n300), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n458), .B1(new_n310), .B2(new_n299), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n492), .B1(new_n304), .B2(new_n288), .ZN(new_n497));
  AOI211_X1 g296(.A(new_n299), .B(new_n497), .C1(new_n487), .C2(new_n489), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT38), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n495), .B(new_n496), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n312), .A2(new_n357), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n383), .A2(new_n384), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(KEYINPUT88), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n397), .A2(new_n390), .ZN(new_n505));
  OAI221_X1 g304(.A(new_n504), .B1(KEYINPUT88), .B2(new_n503), .C1(new_n505), .C2(new_n384), .ZN(new_n506));
  OR3_X1    g305(.A1(new_n505), .A2(KEYINPUT39), .A3(new_n384), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n403), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n407), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n501), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n457), .A2(new_n500), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n475), .A2(KEYINPUT36), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n483), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n478), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT103), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(new_n364), .ZN(new_n523));
  XNOR2_X1  g322(.A(G183gat), .B(G211gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G57gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(G64gat), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT100), .B(G57gat), .Z(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(G64gat), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT101), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI22_X1  g338(.A1(new_n530), .A2(new_n536), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G127gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(G1gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n546), .B1(new_n548), .B2(G1gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT95), .B1(new_n546), .B2(G1gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n547), .B(new_n549), .C1(KEYINPUT95), .C2(G8gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n541), .B2(new_n540), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n545), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n545), .A2(new_n556), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n526), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n545), .A2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n556), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n525), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT15), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n565), .B2(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OR3_X1    g372(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OR4_X1    g375(.A1(new_n575), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n576), .A2(new_n577), .B1(G29gat), .B2(G36gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n565), .A2(KEYINPUT15), .ZN(new_n580));
  NAND2_X1  g379(.A1(G29gat), .A2(G36gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n574), .A2(new_n572), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT7), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n588), .B1(new_n587), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G232gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n330), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n585), .A2(new_n596), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n583), .B1(new_n571), .B2(new_n578), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT17), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n595), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n599), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n606), .A2(new_n607), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n611), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n612), .B2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n521), .B1(new_n564), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(KEYINPUT103), .A3(new_n563), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT106), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  INV_X1    g428(.A(new_n540), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n587), .A2(new_n592), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n588), .A2(KEYINPUT105), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n595), .A2(new_n540), .A3(KEYINPUT104), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT104), .B1(new_n595), .B2(new_n540), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n629), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n596), .A2(new_n630), .A3(KEYINPUT10), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n628), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(new_n636), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n630), .B2(new_n633), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n627), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n626), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n637), .A2(new_n638), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n627), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n645), .B(new_n625), .C1(new_n627), .C2(new_n641), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n620), .A2(new_n622), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n585), .A2(new_n650), .A3(new_n554), .A4(new_n553), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT96), .B1(new_n555), .B2(new_n600), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n555), .A2(new_n600), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n656));
  NAND2_X1  g455(.A1(G229gat), .A2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n601), .B(new_n555), .C1(new_n600), .C2(new_n603), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n653), .A2(KEYINPUT18), .A3(new_n661), .A4(new_n657), .ZN(new_n662));
  XNOR2_X1  g461(.A(G113gat), .B(G141gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G169gat), .B(G197gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT12), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n657), .A3(new_n661), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT18), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n653), .A2(KEYINPUT97), .A3(new_n661), .A4(new_n657), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n669), .B1(new_n675), .B2(KEYINPUT99), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT99), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n672), .A2(new_n677), .A3(new_n673), .A4(new_n674), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n675), .A2(new_n660), .A3(new_n662), .ZN(new_n679));
  INV_X1    g478(.A(new_n668), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n676), .A2(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n649), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n520), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n458), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n501), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT16), .B(G8gat), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(G8gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(G1325gat));
  INV_X1    g493(.A(new_n683), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n518), .A2(KEYINPUT107), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n516), .A2(new_n697), .A3(new_n517), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G15gat), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n352), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(G15gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n695), .B2(new_n703), .ZN(G1326gat));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n480), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT43), .B(G22gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NOR3_X1   g506(.A1(new_n681), .A2(new_n563), .A3(new_n647), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n520), .A2(new_n619), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n458), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  AND3_X1   g510(.A1(new_n483), .A2(new_n515), .A3(new_n518), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n619), .B1(new_n712), .B2(new_n477), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT44), .B(new_n619), .C1(new_n712), .C2(new_n477), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n708), .B(KEYINPUT108), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n458), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n711), .A2(new_n720), .ZN(G1328gat));
  AND2_X1   g520(.A1(new_n312), .A2(new_n357), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n709), .A2(G36gat), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n719), .B2(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1329gat));
  OAI21_X1  g526(.A(G43gat), .B1(new_n719), .B2(new_n518), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n709), .A2(G43gat), .A3(new_n702), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n699), .A3(new_n716), .A4(new_n718), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n733), .A2(new_n734), .A3(G43gat), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n733), .B2(G43gat), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n735), .A2(new_n736), .A3(new_n729), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n732), .B1(new_n737), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g537(.A(G50gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n709), .B2(new_n457), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n480), .A2(G50gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n719), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT48), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n744), .B(new_n740), .C1(new_n719), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1331gat));
  AND4_X1   g545(.A1(new_n681), .A2(new_n620), .A3(new_n622), .A4(new_n647), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n520), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n458), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(new_n529), .ZN(G1332gat));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n722), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  AND2_X1   g554(.A1(new_n520), .A2(new_n747), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n352), .B(KEYINPUT111), .Z(new_n757));
  AOI21_X1  g556(.A(G71gat), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(G71gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n748), .A2(new_n700), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g561(.A1(new_n756), .A2(new_n480), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n684), .A2(new_n590), .A3(new_n647), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n675), .A2(KEYINPUT99), .ZN(new_n768));
  INV_X1    g567(.A(new_n669), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n678), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n679), .A2(new_n680), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n563), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n619), .B(new_n773), .C1(new_n712), .C2(new_n477), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n767), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n767), .B1(new_n774), .B2(new_n775), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n766), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n772), .A2(new_n563), .A3(new_n648), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n715), .A2(new_n684), .A3(new_n716), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G85gat), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n765), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n774), .B(new_n775), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n779), .B1(new_n787), .B2(new_n767), .ZN(new_n788));
  OAI211_X1 g587(.A(KEYINPUT113), .B(new_n784), .C1(new_n788), .C2(new_n766), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1336gat));
  NOR3_X1   g589(.A1(new_n722), .A2(G92gat), .A3(new_n648), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n715), .A2(new_n501), .A3(new_n716), .A4(new_n782), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n787), .A2(new_n791), .B1(new_n794), .B2(G92gat), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n793), .A2(new_n797), .B1(new_n796), .B2(new_n798), .ZN(G1337gat));
  NAND3_X1  g598(.A1(new_n717), .A2(new_n699), .A3(new_n782), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G99gat), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n702), .A2(G99gat), .A3(new_n648), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n788), .B2(new_n802), .ZN(G1338gat));
  OR3_X1    g602(.A1(new_n457), .A2(G106gat), .A3(new_n648), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n715), .A2(new_n480), .A3(new_n716), .A4(new_n782), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n804), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n787), .A2(new_n810), .B1(new_n806), .B2(G106gat), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n805), .A2(new_n809), .B1(new_n808), .B2(new_n811), .ZN(G1339gat));
  AND4_X1   g611(.A1(new_n681), .A2(new_n620), .A3(new_n622), .A4(new_n648), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  AOI211_X1 g613(.A(KEYINPUT54), .B(new_n628), .C1(new_n637), .C2(new_n638), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n625), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  INV_X1    g616(.A(new_n628), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n644), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(KEYINPUT114), .A3(new_n626), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n644), .B2(new_n627), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n637), .A2(new_n628), .A3(new_n638), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n816), .A2(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT115), .B1(new_n823), .B2(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n822), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n815), .A2(new_n814), .A3(new_n625), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT114), .B1(new_n819), .B2(new_n626), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n667), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n655), .A2(new_n659), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n657), .B1(new_n653), .B2(new_n661), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n676), .A2(new_n678), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT55), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n646), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n832), .A2(new_n619), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n646), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n681), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(new_n832), .B1(new_n647), .B2(new_n840), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(new_n619), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n813), .B1(new_n847), .B2(new_n564), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n501), .A2(new_n458), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n457), .A2(new_n475), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n772), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n848), .A2(new_n480), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n352), .A3(new_n849), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT117), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n772), .A2(G113gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(G1340gat));
  AOI21_X1  g660(.A(G120gat), .B1(new_n854), .B2(new_n647), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n647), .A2(G120gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n859), .B2(new_n863), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n858), .B2(new_n564), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n853), .A2(G127gat), .A3(new_n564), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1342gat));
  OAI21_X1  g666(.A(G134gat), .B1(new_n858), .B2(new_n621), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n621), .A2(G134gat), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OR3_X1    g669(.A1(new_n853), .A2(KEYINPUT118), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT118), .B1(new_n853), .B2(new_n870), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n871), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(G1343gat));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n850), .B1(new_n517), .B2(new_n516), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT119), .B1(new_n823), .B2(KEYINPUT55), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n828), .A2(new_n880), .A3(new_n830), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n842), .A2(new_n772), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n840), .A2(new_n647), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n621), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n843), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n564), .ZN(new_n887));
  INV_X1    g686(.A(new_n813), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n457), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n878), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n848), .A2(KEYINPUT57), .A3(new_n457), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n891), .A2(new_n681), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(G141gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n877), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n699), .A2(new_n457), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n851), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n894), .A3(new_n772), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n899), .A3(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  OAI221_X1 g700(.A(new_n898), .B1(new_n877), .B2(new_n901), .C1(new_n893), .C2(new_n894), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n904), .B(G148gat), .C1(new_n897), .C2(new_n647), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n891), .A2(new_n648), .A3(new_n892), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT57), .B1(new_n848), .B2(new_n457), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n563), .B1(new_n885), .B2(new_n843), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n890), .B(new_n480), .C1(new_n908), .C2(new_n813), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n647), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n878), .A2(KEYINPUT59), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n906), .A2(KEYINPUT59), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n905), .B1(new_n913), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n364), .A3(new_n563), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n891), .A2(new_n564), .A3(new_n892), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n364), .ZN(G1346gat));
  AOI21_X1  g716(.A(G162gat), .B1(new_n897), .B2(new_n619), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n891), .A2(new_n892), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n621), .A2(new_n365), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1347gat));
  NOR3_X1   g720(.A1(new_n722), .A2(KEYINPUT121), .A3(new_n684), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n501), .B2(new_n458), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n757), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n856), .A2(new_n772), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT123), .B1(new_n929), .B2(G169gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n848), .A2(new_n684), .A3(new_n722), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n852), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n772), .A2(new_n268), .A3(new_n269), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n930), .A2(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT124), .ZN(G1348gat));
  AND4_X1   g735(.A1(new_n647), .A2(new_n856), .A3(new_n927), .A4(new_n928), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n647), .A2(new_n262), .ZN(new_n938));
  OAI22_X1  g737(.A1(new_n937), .A2(new_n262), .B1(new_n933), .B2(new_n938), .ZN(G1349gat));
  AND4_X1   g738(.A1(new_n563), .A2(new_n856), .A3(new_n927), .A4(new_n928), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n563), .A2(new_n227), .A3(new_n229), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n940), .A2(new_n226), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g742(.A1(new_n856), .A2(new_n619), .A3(new_n927), .A4(new_n928), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G190gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n948), .A3(G190gat), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n947), .B1(new_n946), .B2(new_n949), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n619), .A2(new_n230), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n950), .A2(new_n951), .B1(new_n933), .B2(new_n952), .ZN(G1351gat));
  NOR2_X1   g752(.A1(new_n922), .A2(new_n924), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n699), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n910), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(G197gat), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(new_n681), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n932), .A2(new_n896), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n772), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n958), .A2(new_n961), .ZN(G1352gat));
  INV_X1    g761(.A(new_n955), .ZN(new_n963));
  OAI21_X1  g762(.A(G204gat), .B1(new_n911), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n648), .A2(G204gat), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n959), .A2(KEYINPUT62), .A3(new_n965), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(G1353gat));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n907), .A2(new_n909), .A3(new_n563), .A4(new_n955), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G211gat), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n970), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n910), .A2(KEYINPUT126), .A3(new_n563), .A4(new_n955), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n206), .B1(new_n970), .B2(new_n971), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT63), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(KEYINPUT127), .A3(new_n978), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n959), .A2(G211gat), .A3(new_n564), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n976), .B2(new_n977), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n979), .A2(new_n983), .ZN(G1354gat));
  AOI211_X1 g783(.A(new_n621), .B(new_n956), .C1(new_n207), .C2(new_n208), .ZN(new_n985));
  AOI21_X1  g784(.A(G218gat), .B1(new_n960), .B2(new_n619), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


