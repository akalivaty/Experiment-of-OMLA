//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  OR2_X1    g0006(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n209));
  AND3_X1   g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT66), .Z(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n203), .A2(new_n205), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n216), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n208), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n212), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n223), .B1(KEYINPUT1), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n221), .A2(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n202), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n248), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT75), .ZN(new_n255));
  INV_X1    g0055(.A(G169), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT69), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT69), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  OAI211_X1 g0062(.A(G232), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  OAI211_X1 g0064(.A(G226), .B(new_n264), .C1(new_n261), .C2(new_n262), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  OAI21_X1  g0072(.A(G274), .B1(new_n272), .B2(new_n217), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  AND2_X1   g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n268), .ZN(new_n280));
  INV_X1    g0080(.A(new_n276), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT68), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n269), .A2(new_n276), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n277), .A2(new_n282), .B1(new_n225), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT13), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT13), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n271), .A2(new_n288), .A3(new_n285), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n256), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT14), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT74), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g0092(.A(KEYINPUT13), .B(new_n284), .C1(new_n267), .C2(new_n270), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(new_n271), .B2(new_n285), .ZN(new_n294));
  OAI21_X1  g0094(.A(G169), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT74), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT14), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n291), .B(G169), .C1(new_n293), .C2(new_n294), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n287), .A2(G179), .A3(new_n289), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n292), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n218), .A2(G33), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n208), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n217), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT11), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n304), .A2(KEYINPUT11), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT73), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n306), .B1(new_n275), .B2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G68), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT12), .B1(new_n315), .B2(G68), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n315), .A2(KEYINPUT12), .A3(G68), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n311), .B2(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n300), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n293), .A2(new_n294), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n323), .B2(G190), .ZN(new_n324));
  OAI21_X1  g0124(.A(G200), .B1(new_n293), .B2(new_n294), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n255), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g0128(.A(KEYINPUT75), .B(new_n326), .C1(new_n300), .C2(new_n321), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n258), .A2(new_n260), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT69), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(G222), .A3(new_n264), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(G223), .A3(G1698), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n261), .A2(new_n262), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G77), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT70), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n269), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT70), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n274), .B1(new_n273), .B2(new_n276), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n281), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G226), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n283), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(G179), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n218), .B1(new_n207), .B2(new_n209), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n301), .A2(G150), .ZN(new_n353));
  OR2_X1    g0153(.A1(KEYINPUT71), .A2(G58), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT71), .A2(G58), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT8), .ZN(new_n357));
  OR2_X1    g0157(.A1(KEYINPUT8), .A2(G58), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n353), .B1(new_n359), .B2(new_n303), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n306), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n315), .A2(G50), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n313), .B2(G50), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n348), .B1(new_n341), .B2(new_n342), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(G169), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n351), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT9), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n361), .A2(KEYINPUT9), .A3(new_n363), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n365), .C2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n365), .A2(G190), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT10), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n369), .A2(new_n370), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n350), .A2(G200), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT10), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n365), .A2(G190), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n367), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n346), .B1(new_n226), .B2(new_n283), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n334), .A2(G232), .A3(new_n264), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n334), .A2(G238), .A3(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n337), .A2(G107), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n381), .B1(new_n385), .B2(new_n270), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G190), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n313), .A2(G77), .ZN(new_n388));
  INV_X1    g0188(.A(new_n315), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n208), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g0191(.A(KEYINPUT8), .B(G58), .Z(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n301), .B1(G20), .B2(G77), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT72), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(new_n303), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n391), .B1(new_n399), .B2(new_n306), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n387), .B(new_n400), .C1(new_n371), .C2(new_n386), .ZN(new_n401));
  INV_X1    g0201(.A(G179), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n386), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n400), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(G169), .C2(new_n386), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT79), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n277), .A2(new_n282), .B1(new_n238), .B2(new_n283), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n347), .B2(G1698), .ZN(new_n410));
  OR2_X1    g0210(.A1(KEYINPUT76), .A2(G33), .ZN(new_n411));
  NAND2_X1  g0211(.A1(KEYINPUT76), .A2(G33), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(KEYINPUT3), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n413), .A3(new_n258), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n269), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n407), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n269), .A2(G232), .A3(new_n276), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n344), .B2(new_n345), .ZN(new_n419));
  INV_X1    g0219(.A(new_n258), .ZN(new_n420));
  AND2_X1   g0220(.A1(KEYINPUT76), .A2(G33), .ZN(new_n421));
  NOR2_X1   g0221(.A1(KEYINPUT76), .A2(G33), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n420), .B1(new_n423), .B2(KEYINPUT3), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n410), .B1(G33), .B2(G87), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n419), .B(KEYINPUT79), .C1(new_n425), .C2(new_n269), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n256), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n419), .B(new_n402), .C1(new_n425), .C2(new_n269), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT78), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n416), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n432), .A2(KEYINPUT78), .A3(new_n402), .A4(new_n419), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n359), .A2(new_n313), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n315), .B2(new_n359), .ZN(new_n437));
  INV_X1    g0237(.A(new_n306), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n202), .B1(new_n354), .B2(new_n355), .ZN(new_n439));
  OAI21_X1  g0239(.A(G20), .B1(new_n439), .B2(new_n220), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n301), .A2(G159), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(G20), .B1(new_n413), .B2(new_n258), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT7), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n202), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT7), .B1(new_n424), .B2(G20), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n438), .B1(new_n447), .B2(KEYINPUT16), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT16), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n332), .A2(new_n218), .A3(new_n333), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n444), .ZN(new_n451));
  OR3_X1    g0251(.A1(new_n257), .A2(KEYINPUT77), .A3(G33), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n260), .A2(KEYINPUT77), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n453), .C1(new_n423), .C2(KEYINPUT3), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n444), .A2(G20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n202), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n449), .B1(new_n457), .B2(new_n442), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n437), .B1(new_n448), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT18), .B1(new_n435), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT17), .ZN(new_n461));
  INV_X1    g0261(.A(new_n437), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT7), .B1(new_n337), .B2(new_n218), .ZN(new_n463));
  INV_X1    g0263(.A(new_n455), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n452), .A2(new_n453), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n411), .A2(new_n412), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n257), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(G68), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n355), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT71), .A2(G58), .ZN(new_n471));
  OAI21_X1  g0271(.A(G68), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(new_n205), .A3(new_n203), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(G20), .B1(G159), .B2(new_n301), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT16), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n421), .A2(new_n422), .A3(new_n257), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n444), .B(new_n218), .C1(new_n476), .C2(new_n420), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G68), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n443), .A2(new_n444), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n474), .B(KEYINPUT16), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n306), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n462), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n408), .A2(new_n416), .A3(G190), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n427), .B2(new_n371), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n461), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n256), .A2(new_n427), .B1(new_n431), .B2(new_n433), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT18), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n427), .A2(new_n371), .ZN(new_n489));
  INV_X1    g0289(.A(new_n483), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n459), .A3(KEYINPUT17), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n460), .A2(new_n485), .A3(new_n488), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n380), .A2(new_n406), .A3(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n328), .A2(new_n329), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n226), .A2(G1698), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT82), .B1(new_n424), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n413), .A2(KEYINPUT82), .A3(new_n258), .A4(new_n497), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G250), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n500), .A2(new_n226), .A3(G1698), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n261), .B2(new_n262), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n270), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT5), .B(G41), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n280), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n270), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(G257), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n256), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n508), .A2(new_n402), .A3(new_n515), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  XOR2_X1   g0320(.A(G97), .B(G107), .Z(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(KEYINPUT6), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(G20), .B1(G77), .B2(new_n301), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n450), .A2(new_n444), .B1(new_n454), .B2(new_n455), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n519), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n306), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT80), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n389), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT80), .B1(new_n315), .B2(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n275), .A2(G33), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n315), .A2(new_n531), .A3(new_n217), .A4(new_n305), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n529), .B(new_n530), .C1(new_n528), .C2(new_n532), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n533), .B(KEYINPUT81), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n517), .A2(new_n518), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n534), .B1(new_n306), .B2(new_n525), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n508), .A2(G190), .A3(new_n515), .ZN(new_n539));
  INV_X1    g0339(.A(new_n515), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n334), .A2(new_n504), .B1(G33), .B2(G283), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n503), .C1(new_n498), .C2(new_n501), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n542), .B2(new_n270), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n538), .B(new_n539), .C1(new_n371), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g0345(.A1(G250), .A2(G1698), .ZN(new_n546));
  INV_X1    g0346(.A(G257), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G1698), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n413), .A2(new_n258), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n466), .A2(G294), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n269), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n511), .A2(new_n510), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n552), .A2(G264), .A3(new_n269), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G190), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n512), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n551), .A2(new_n553), .A3(new_n513), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(G200), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n413), .A2(new_n218), .A3(G87), .A4(new_n258), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(G87), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n562), .A2(KEYINPUT22), .A3(G20), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n261), .B2(new_n262), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n466), .A2(new_n218), .A3(G116), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n218), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n519), .A2(KEYINPUT23), .A3(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n559), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g0373(.A(KEYINPUT24), .B(new_n571), .C1(new_n561), .C2(new_n564), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n306), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT89), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT25), .B1(new_n389), .B2(new_n519), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n389), .A2(KEYINPUT25), .A3(new_n519), .ZN(new_n579));
  INV_X1    g0379(.A(new_n532), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(G107), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n558), .A2(new_n575), .A3(new_n576), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n558), .A2(new_n575), .A3(new_n581), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT89), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n545), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G303), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n261), .A2(new_n262), .A3(new_n586), .ZN(new_n587));
  MUX2_X1   g0387(.A(G257), .B(G264), .S(G1698), .Z(new_n588));
  AND3_X1   g0388(.A1(new_n588), .A2(new_n413), .A3(new_n258), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n270), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n552), .A2(G270), .A3(new_n269), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n591), .A2(new_n512), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(KEYINPUT87), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n332), .A2(G303), .A3(new_n333), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(new_n413), .A3(new_n258), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n269), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n591), .A2(new_n512), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n593), .A2(new_n599), .A3(G200), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n506), .B(new_n218), .C1(G33), .C2(new_n528), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G20), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n306), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n315), .A2(G116), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n580), .B2(G116), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n600), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n593), .A2(new_n599), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(new_n555), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n600), .A2(KEYINPUT88), .A3(new_n609), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OR3_X1    g0416(.A1(new_n509), .A2(KEYINPUT83), .A3(G1), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT83), .B1(new_n509), .B2(G1), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(G250), .A3(new_n269), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n280), .A2(new_n510), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(G238), .A2(G1698), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n226), .B2(G1698), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n413), .A3(new_n258), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n466), .A2(G116), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n622), .B1(new_n627), .B2(new_n269), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n256), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT85), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n398), .B2(new_n532), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n413), .A2(new_n218), .A3(G68), .A4(new_n258), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT19), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n218), .B1(new_n266), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n562), .A2(new_n528), .A3(new_n519), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n218), .A2(G33), .A3(G97), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n634), .A2(new_n635), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n306), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n398), .A2(new_n389), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n396), .A2(new_n580), .A3(KEYINPUT85), .A4(new_n397), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n631), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n269), .B1(new_n625), .B2(new_n626), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n621), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT84), .B1(new_n644), .B2(new_n402), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT84), .ZN(new_n646));
  NOR4_X1   g0446(.A1(new_n643), .A2(new_n621), .A3(new_n646), .A4(G179), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n629), .B(new_n642), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n622), .B(G190), .C1(new_n627), .C2(new_n269), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT86), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n628), .A2(G200), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n644), .A2(KEYINPUT86), .A3(G190), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n580), .A2(G87), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n639), .A2(new_n640), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n651), .A2(new_n652), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n549), .A2(new_n550), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n270), .ZN(new_n659));
  INV_X1    g0459(.A(new_n553), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n659), .A2(new_n402), .A3(new_n660), .A4(new_n512), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n557), .B2(G169), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n575), .B2(new_n581), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n256), .B1(new_n606), .B2(new_n608), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT21), .B1(new_n613), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n593), .A2(new_n599), .A3(new_n665), .A4(KEYINPUT21), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n597), .A2(new_n598), .A3(new_n402), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n609), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n616), .A2(new_n664), .A3(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n496), .A2(new_n585), .A3(new_n672), .ZN(G372));
  NAND2_X1  g0473(.A1(new_n460), .A2(new_n488), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n485), .A2(new_n492), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n405), .B1(new_n324), .B2(new_n325), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n300), .B2(new_n321), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT91), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI211_X1 g0480(.A(KEYINPUT91), .B(new_n677), .C1(new_n300), .C2(new_n321), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n374), .A2(new_n379), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n367), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n496), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n537), .A2(new_n544), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n584), .A2(new_n582), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n629), .B(new_n642), .C1(G179), .C2(new_n628), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n652), .A2(new_n655), .A3(new_n649), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n686), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT90), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT90), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n686), .A2(new_n687), .A3(new_n694), .A4(new_n691), .ZN(new_n695));
  INV_X1    g0495(.A(new_n663), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n671), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  OR3_X1    g0498(.A1(new_n537), .A2(KEYINPUT26), .A3(new_n690), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n537), .B2(new_n657), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n688), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n684), .B1(new_n685), .B2(new_n703), .ZN(G369));
  NAND3_X1  g0504(.A1(new_n275), .A2(new_n218), .A3(G13), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n575), .B2(new_n581), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT92), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n663), .B1(new_n713), .B2(new_n687), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n663), .A2(new_n711), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n609), .A2(new_n711), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n616), .A2(new_n671), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n671), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n711), .B1(new_n666), .B2(new_n670), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n716), .B1(new_n717), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(G399));
  NOR2_X1   g0528(.A1(new_n635), .A2(G116), .ZN(new_n729));
  INV_X1    g0529(.A(G41), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n213), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n731), .A3(G1), .ZN(new_n732));
  INV_X1    g0532(.A(new_n222), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(new_n731), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  OR3_X1    g0535(.A1(new_n537), .A2(new_n657), .A3(KEYINPUT26), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT26), .B1(new_n537), .B2(new_n690), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n736), .A2(new_n688), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n585), .A2(new_n691), .A3(new_n697), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n710), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n710), .B1(new_n698), .B2(new_n702), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n741), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n672), .A2(new_n585), .A3(new_n711), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n668), .A2(new_n554), .A3(new_n644), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n516), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n554), .A2(new_n644), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n543), .A2(KEYINPUT30), .A3(new_n668), .A4(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n557), .A2(new_n644), .A3(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n613), .A2(new_n516), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n749), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n710), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n746), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n745), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n735), .B1(new_n761), .B2(G1), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT94), .Z(G364));
  INV_X1    g0563(.A(new_n722), .ZN(new_n764));
  INV_X1    g0564(.A(G13), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G45), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n768), .A2(G1), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n731), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n764), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n721), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n217), .B1(G20), .B2(new_n256), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n424), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n213), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n253), .A2(new_n509), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n781), .B(new_n782), .C1(new_n509), .C2(new_n222), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n334), .A2(new_n213), .ZN(new_n784));
  INV_X1    g0584(.A(G355), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n785), .B1(G116), .B2(new_n213), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n779), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n772), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n218), .A2(new_n402), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G190), .A3(new_n371), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n790), .A2(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n218), .A2(G179), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n792), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(G329), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n789), .A2(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n555), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n334), .B1(G326), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n555), .A2(G179), .A3(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n218), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n796), .A2(new_n555), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n805), .A2(G294), .B1(new_n807), .B2(G283), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n800), .A2(G190), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT33), .B(G317), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n796), .A2(G190), .A3(G200), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n809), .A2(new_n810), .B1(new_n812), .B2(G303), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n799), .A2(new_n802), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT96), .B(G159), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n797), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT32), .ZN(new_n817));
  INV_X1    g0617(.A(new_n790), .ZN(new_n818));
  INV_X1    g0618(.A(new_n793), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(new_n356), .B1(new_n819), .B2(G77), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n809), .A2(G68), .B1(new_n812), .B2(G87), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n817), .A2(new_n334), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n801), .A2(G50), .B1(new_n807), .B2(G107), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n528), .B2(new_n804), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n814), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT97), .ZN(new_n826));
  INV_X1    g0626(.A(new_n778), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n825), .B2(KEYINPUT97), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n788), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n777), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n721), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n774), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  OAI211_X1 g0633(.A(new_n401), .B(new_n405), .C1(new_n400), .C2(new_n711), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT99), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n404), .B1(new_n386), .B2(G169), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n386), .A2(new_n402), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n835), .B1(new_n838), .B2(new_n710), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n405), .A2(KEYINPUT99), .A3(new_n711), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n834), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT100), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT100), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n834), .B(new_n843), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n742), .B(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n772), .B1(new_n846), .B2(new_n760), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n760), .B2(new_n846), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n780), .B1(G132), .B2(new_n798), .ZN(new_n849));
  INV_X1    g0649(.A(new_n356), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n850), .A2(new_n804), .B1(new_n221), .B2(new_n811), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n806), .A2(new_n202), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n815), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n818), .A2(G143), .B1(new_n819), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G150), .ZN(new_n856));
  INV_X1    g0656(.A(new_n809), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G137), .B2(new_n801), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n849), .B(new_n853), .C1(new_n859), .C2(KEYINPUT34), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(KEYINPUT34), .B2(new_n859), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n334), .B1(G107), .B2(new_n812), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT98), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G116), .A2(new_n819), .B1(new_n798), .B2(G311), .ZN(new_n864));
  INV_X1    g0664(.A(G294), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(new_n790), .ZN(new_n866));
  INV_X1    g0666(.A(G283), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n857), .A2(new_n867), .B1(new_n528), .B2(new_n804), .ZN(new_n868));
  INV_X1    g0668(.A(new_n801), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n869), .A2(new_n586), .B1(new_n806), .B2(new_n562), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n863), .A2(new_n866), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n778), .B1(new_n861), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n772), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n778), .A2(new_n775), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n208), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n872), .B(new_n875), .C1(new_n845), .C2(new_n776), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n848), .A2(new_n876), .ZN(G384));
  NOR2_X1   g0677(.A1(new_n766), .A2(new_n275), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n491), .A2(new_n459), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n447), .A2(KEYINPUT16), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n462), .B1(new_n481), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n486), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n708), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n880), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n482), .A2(new_n486), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n482), .A2(new_n884), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n888), .A2(new_n880), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n885), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n493), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(KEYINPUT102), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n879), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n888), .A2(new_n880), .A3(new_n889), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n891), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n493), .A2(new_n482), .A3(new_n884), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n898), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT104), .B1(new_n901), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n322), .A2(new_n710), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT102), .A4(KEYINPUT38), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n891), .A2(new_n887), .B1(new_n493), .B2(new_n893), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(KEYINPUT38), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT102), .B1(new_n913), .B2(KEYINPUT38), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT39), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n907), .B1(new_n904), .B2(new_n905), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n896), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n879), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT104), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n910), .A2(new_n911), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n405), .A2(new_n710), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n742), .B2(new_n845), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n321), .A2(new_n710), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n290), .A2(KEYINPUT74), .A3(new_n291), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n296), .B1(new_n295), .B2(KEYINPUT14), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n298), .A2(new_n299), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n321), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n327), .B(new_n925), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n321), .B(new_n710), .C1(new_n300), .C2(new_n326), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n895), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n900), .A2(new_n936), .A3(new_n912), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n935), .A2(new_n937), .B1(new_n674), .B2(new_n708), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n496), .B(new_n741), .C1(new_n742), .C2(new_n744), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n684), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(G330), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n931), .A2(new_n932), .B1(new_n842), .B2(new_n844), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n755), .A2(KEYINPUT105), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT105), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n754), .A2(new_n946), .A3(new_n710), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n756), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n746), .A2(new_n948), .A3(new_n758), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n944), .B(new_n949), .C1(new_n914), .C2(new_n915), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(new_n954), .A3(new_n951), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n933), .A2(new_n949), .A3(new_n845), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n918), .A2(new_n951), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n953), .A2(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n496), .A2(new_n949), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n943), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n878), .B1(new_n942), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n942), .B2(new_n961), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n522), .A2(KEYINPUT35), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n964), .A2(G116), .A3(new_n219), .A4(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n733), .A2(new_n208), .A3(new_n439), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n249), .B(KEYINPUT101), .ZN(new_n969));
  OAI211_X1 g0769(.A(G1), .B(new_n765), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n967), .A3(new_n970), .ZN(G367));
  OAI21_X1  g0771(.A(new_n686), .B1(new_n538), .B2(new_n711), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n537), .A2(new_n711), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n723), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n655), .A2(new_n711), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n691), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n688), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n972), .A2(new_n696), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n537), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT107), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n710), .B1(new_n988), .B2(KEYINPUT107), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n717), .A2(new_n726), .A3(new_n974), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n989), .A2(new_n990), .B1(KEYINPUT42), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(KEYINPUT42), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n978), .A2(new_n982), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n984), .A2(new_n985), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n985), .ZN(new_n996));
  INV_X1    g0796(.A(new_n994), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n983), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n731), .B(KEYINPUT41), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n717), .A2(new_n726), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n764), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(KEYINPUT109), .A3(new_n722), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n717), .A2(new_n726), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1004), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n727), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n974), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(KEYINPUT44), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT44), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n727), .B2(new_n974), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n974), .B(new_n715), .C1(new_n714), .C2(new_n725), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT45), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n723), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n724), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1007), .A2(new_n1017), .A3(new_n761), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n999), .B1(new_n1019), .B2(new_n761), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n995), .B(new_n998), .C1(new_n1020), .C2(new_n770), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n781), .A2(new_n244), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n779), .B1(new_n398), .B2(new_n213), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n772), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n812), .A2(G116), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(G317), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n790), .A2(new_n586), .B1(new_n797), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G283), .B2(new_n819), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n807), .A2(G97), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G107), .A2(new_n805), .B1(new_n809), .B2(G294), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n424), .B1(G311), .B2(new_n801), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n337), .B1(G77), .B2(new_n807), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n818), .A2(G150), .B1(new_n798), .B2(G137), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n221), .C2(new_n793), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G143), .A2(new_n801), .B1(new_n809), .B2(new_n854), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n805), .A2(G68), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n850), .C2(new_n811), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1027), .A2(new_n1034), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT47), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1024), .B1(new_n1042), .B2(new_n778), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n981), .B2(new_n830), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1021), .A2(new_n1044), .ZN(G387));
  NAND2_X1  g0845(.A1(new_n1007), .A2(new_n770), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n857), .A2(new_n359), .B1(new_n202), .B2(new_n793), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT113), .Z(new_n1048));
  INV_X1    g0848(.A(new_n398), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n805), .ZN(new_n1050));
  INV_X1    g0850(.A(G159), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1031), .B1(new_n869), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n424), .B1(new_n221), .B2(new_n790), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n811), .A2(new_n208), .B1(new_n797), .B2(new_n856), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT112), .Z(new_n1056));
  NAND4_X1  g0856(.A1(new_n1048), .A2(new_n1050), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n424), .B1(G326), .B2(new_n798), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n804), .A2(new_n867), .B1(new_n811), .B2(new_n865), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n818), .A2(G317), .B1(new_n819), .B2(G303), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n857), .B2(new_n794), .C1(new_n791), .C2(new_n869), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1058), .B1(new_n602), .B2(new_n806), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1057), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT114), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n827), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n241), .A2(G45), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT111), .Z(new_n1073));
  NAND2_X1  g0873(.A1(new_n392), .A2(new_n221), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT50), .Z(new_n1075));
  INV_X1    g0875(.A(new_n729), .ZN(new_n1076));
  AOI211_X1 g0876(.A(G45), .B(new_n1076), .C1(G68), .C2(G77), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n781), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(G107), .B2(new_n213), .C1(new_n729), .C2(new_n784), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n873), .B1(new_n1080), .B2(new_n779), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1071), .B(new_n1081), .C1(new_n717), .C2(new_n830), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1007), .A2(new_n761), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n771), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1007), .A2(new_n761), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1046), .B(new_n1082), .C1(new_n1084), .C2(new_n1085), .ZN(G393));
  NAND3_X1  g0886(.A1(new_n1017), .A2(new_n770), .A3(new_n1018), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n779), .B1(new_n528), .B2(new_n213), .C1(new_n781), .C2(new_n248), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n772), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n869), .A2(new_n1028), .B1(new_n794), .B2(new_n790), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G116), .A2(new_n805), .B1(new_n809), .B2(G303), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1092), .A2(KEYINPUT116), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(KEYINPUT116), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n519), .A2(new_n806), .B1(new_n811), .B2(new_n867), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n793), .A2(new_n865), .B1(new_n797), .B2(new_n791), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n334), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n804), .A2(new_n208), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n392), .B2(new_n819), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n221), .B2(new_n857), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT115), .Z(new_n1102));
  OAI22_X1  g0902(.A1(new_n869), .A2(new_n856), .B1(new_n1051), .B2(new_n790), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT51), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n780), .B1(G143), .B2(new_n798), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n812), .A2(G68), .B1(new_n807), .B2(G87), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1098), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1089), .B1(new_n1108), .B2(new_n778), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n974), .B2(new_n830), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1019), .A2(new_n771), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1007), .A2(new_n761), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1087), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(G390));
  INV_X1    g0913(.A(new_n911), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n924), .B2(new_n934), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n916), .A2(new_n920), .A3(new_n919), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n923), .B1(new_n740), .B2(new_n845), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n934), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n908), .A2(new_n1114), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n759), .A2(new_n845), .A3(G330), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1124), .A2(new_n934), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1118), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n949), .A2(G330), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n944), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n496), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n940), .A2(new_n684), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT117), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n940), .A2(new_n684), .A3(KEYINPUT117), .A4(new_n1131), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1127), .A2(new_n944), .B1(new_n1124), .B2(new_n934), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1119), .B1(new_n1124), .B2(new_n934), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n933), .B1(new_n1127), .B2(new_n845), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1136), .A2(new_n924), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1134), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n731), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT118), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1134), .A2(new_n1139), .A3(new_n1135), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(new_n1126), .C2(new_n1129), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1118), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n910), .A2(new_n921), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1122), .B1(new_n1147), .B2(new_n1115), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1148), .B2(new_n1128), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1141), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n873), .B1(new_n359), .B2(new_n874), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n790), .A2(new_n602), .B1(new_n797), .B2(new_n865), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G97), .B2(new_n819), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n337), .C1(new_n562), .C2(new_n811), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n857), .A2(new_n519), .B1(new_n869), .B2(new_n867), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1155), .A2(new_n852), .A3(new_n1099), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1158), .A2(KEYINPUT119), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(KEYINPUT119), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n811), .A2(new_n856), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n869), .A2(new_n1163), .B1(new_n1051), .B2(new_n804), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G137), .B2(new_n809), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n818), .A2(G132), .B1(new_n819), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(G125), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n797), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n337), .B1(G50), .B2(new_n807), .ZN(new_n1172));
  AND4_X1   g0972(.A1(new_n1162), .A2(new_n1165), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1159), .A2(new_n1160), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1152), .B1(new_n1174), .B2(new_n827), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1147), .B2(new_n775), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1130), .B2(new_n770), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1151), .A2(new_n1177), .ZN(G378));
  INV_X1    g0978(.A(new_n1128), .ZN(new_n1179));
  AOI221_X4 g0979(.A(new_n710), .B1(new_n842), .B2(new_n844), .C1(new_n698), .C2(new_n702), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n933), .B1(new_n1180), .B2(new_n923), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n910), .A2(new_n921), .B1(new_n1181), .B2(new_n1114), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n1182), .B2(new_n1122), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n364), .A2(new_n884), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n380), .B(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n953), .A2(new_n955), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n943), .B1(new_n957), .B2(new_n956), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(KEYINPUT106), .B(KEYINPUT40), .C1(new_n956), .C2(new_n937), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n954), .B1(new_n950), .B2(new_n951), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1194), .B(new_n1192), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n939), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1192), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1203), .A2(new_n922), .A3(new_n938), .A4(new_n1198), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1187), .A2(new_n1205), .A3(KEYINPUT57), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1186), .A2(new_n1184), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n771), .C1(KEYINPUT57), .C2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n770), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1202), .A2(new_n775), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n874), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n772), .B1(G50), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n259), .A2(new_n730), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT120), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n221), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n730), .B2(new_n780), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n850), .A2(new_n806), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n869), .A2(new_n602), .B1(new_n811), .B2(new_n208), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(G97), .C2(new_n809), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1039), .B1(new_n867), .B2(new_n797), .C1(new_n519), .C2(new_n790), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1049), .B2(new_n819), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n730), .A3(new_n1221), .A4(new_n780), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n1223), .B2(KEYINPUT58), .ZN(new_n1224));
  INV_X1    g1024(.A(G137), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n790), .A2(new_n1163), .B1(new_n793), .B2(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n809), .A2(G132), .B1(new_n812), .B2(new_n1167), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1169), .B2(new_n869), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G150), .C2(new_n805), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1214), .B1(G124), .B2(new_n798), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1232), .B1(new_n806), .B2(new_n815), .C1(new_n1229), .C2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1224), .B1(KEYINPUT58), .B2(new_n1223), .C1(new_n1231), .C2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1212), .B1(new_n1235), .B2(new_n778), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1210), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1209), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1208), .A2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n934), .A2(new_n775), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n772), .B1(G68), .B2(new_n1211), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n857), .A2(new_n602), .B1(new_n528), .B2(new_n811), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G294), .B2(new_n801), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n793), .A2(new_n519), .B1(new_n797), .B2(new_n586), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G283), .B2(new_n818), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n334), .B1(G77), .B2(new_n807), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1050), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n780), .A2(new_n1217), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT121), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n790), .A2(new_n1225), .B1(new_n797), .B2(new_n1163), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G150), .B2(new_n819), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G50), .A2(new_n805), .B1(new_n809), .B2(new_n1167), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n801), .A2(G132), .B1(new_n812), .B2(G159), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1248), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1242), .B1(new_n1256), .B2(new_n778), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1139), .A2(new_n770), .B1(new_n1241), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n999), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1143), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1139), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(G381));
  XOR2_X1   g1062(.A(G375), .B(KEYINPUT122), .Z(new_n1263));
  INV_X1    g1063(.A(G390), .ZN(new_n1264));
  INV_X1    g1064(.A(G384), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OR2_X1    g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1266), .A2(G387), .A3(new_n1267), .A4(G381), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1263), .A2(new_n1151), .A3(new_n1177), .A4(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT123), .ZN(G407));
  INV_X1    g1070(.A(G213), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(G343), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G378), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1263), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G407), .A2(new_n1275), .ZN(G409));
  XNOR2_X1  g1076(.A(G393), .B(G396), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1021), .A2(G390), .A3(new_n1044), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G390), .B1(new_n1021), .B2(new_n1044), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(new_n1264), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(new_n832), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1021), .A2(G390), .A3(new_n1044), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1261), .A2(KEYINPUT60), .A3(new_n1143), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n771), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1261), .B1(KEYINPUT60), .B2(new_n1143), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1258), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1265), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G384), .B(new_n1258), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1208), .A2(G378), .A3(new_n1239), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1187), .A2(new_n1205), .A3(new_n1259), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1151), .B(new_n1177), .C1(new_n1238), .C2(new_n1295), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1272), .B(new_n1293), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1293), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1273), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1298), .A2(new_n1303), .A3(KEYINPUT126), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1272), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1272), .A2(G2897), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1293), .B(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1303), .B2(KEYINPUT126), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1286), .B1(new_n1304), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT124), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1297), .B2(KEYINPUT63), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1301), .A2(KEYINPUT124), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1307), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1293), .B(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1285), .B(new_n1317), .C1(new_n1305), .C2(new_n1319), .ZN(new_n1320));
  AND4_X1   g1120(.A1(KEYINPUT63), .A2(new_n1299), .A3(new_n1273), .A4(new_n1300), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1316), .A2(KEYINPUT125), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT125), .B1(new_n1316), .B2(new_n1322), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1311), .B1(new_n1323), .B2(new_n1324), .ZN(G405));
  AOI21_X1  g1125(.A(G378), .B1(new_n1208), .B2(new_n1239), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1326), .A2(new_n1300), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1300), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(KEYINPUT127), .A3(new_n1294), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1294), .A2(KEYINPUT127), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1327), .A2(new_n1331), .A3(new_n1328), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1286), .ZN(G402));
endmodule


