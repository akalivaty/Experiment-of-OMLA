

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587;

  XNOR2_X1 U319 ( .A(n299), .B(n298), .ZN(n303) );
  XNOR2_X1 U320 ( .A(n297), .B(KEYINPUT31), .ZN(n298) );
  XNOR2_X1 U321 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n394) );
  XNOR2_X1 U322 ( .A(n395), .B(n394), .ZN(n569) );
  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n311) );
  XNOR2_X1 U324 ( .A(n577), .B(n311), .ZN(n345) );
  XNOR2_X1 U325 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U326 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U327 ( .A(G85GAT), .ZN(n287) );
  NAND2_X1 U328 ( .A1(G92GAT), .A2(n287), .ZN(n290) );
  INV_X1 U329 ( .A(G92GAT), .ZN(n288) );
  NAND2_X1 U330 ( .A1(n288), .A2(G85GAT), .ZN(n289) );
  NAND2_X1 U331 ( .A1(n290), .A2(n289), .ZN(n292) );
  XNOR2_X1 U332 ( .A(G99GAT), .B(G106GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n323) );
  INV_X1 U334 ( .A(n323), .ZN(n293) );
  NAND2_X1 U335 ( .A1(n293), .A2(KEYINPUT32), .ZN(n296) );
  INV_X1 U336 ( .A(KEYINPUT32), .ZN(n294) );
  NAND2_X1 U337 ( .A1(n323), .A2(n294), .ZN(n295) );
  NAND2_X1 U338 ( .A1(n296), .A2(n295), .ZN(n299) );
  NAND2_X1 U339 ( .A1(G230GAT), .A2(G233GAT), .ZN(n297) );
  INV_X1 U340 ( .A(n303), .ZN(n301) );
  XOR2_X1 U341 ( .A(G57GAT), .B(KEYINPUT13), .Z(n348) );
  XNOR2_X1 U342 ( .A(n348), .B(KEYINPUT33), .ZN(n302) );
  INV_X1 U343 ( .A(n302), .ZN(n300) );
  NAND2_X1 U344 ( .A1(n301), .A2(n300), .ZN(n305) );
  NAND2_X1 U345 ( .A1(n303), .A2(n302), .ZN(n304) );
  NAND2_X1 U346 ( .A1(n305), .A2(n304), .ZN(n306) );
  XOR2_X1 U347 ( .A(G176GAT), .B(G64GAT), .Z(n382) );
  XNOR2_X1 U348 ( .A(n306), .B(n382), .ZN(n310) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  XOR2_X1 U350 ( .A(G78GAT), .B(G148GAT), .Z(n308) );
  XNOR2_X1 U351 ( .A(KEYINPUT70), .B(G204GAT), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n411) );
  XOR2_X1 U353 ( .A(n448), .B(n411), .Z(n309) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n577) );
  XNOR2_X1 U355 ( .A(KEYINPUT108), .B(n345), .ZN(n538) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G43GAT), .Z(n313) );
  XNOR2_X1 U357 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n340) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n314), .B(KEYINPUT74), .ZN(n386) );
  XNOR2_X1 U361 ( .A(n340), .B(n386), .ZN(n327) );
  XOR2_X1 U362 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n316) );
  XNOR2_X1 U363 ( .A(G134GAT), .B(KEYINPUT73), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U365 ( .A(KEYINPUT10), .B(KEYINPUT72), .Z(n318) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U368 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U369 ( .A(G162GAT), .B(KEYINPUT71), .Z(n322) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(G218GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n412) );
  XNOR2_X1 U372 ( .A(n412), .B(n323), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n560) );
  XOR2_X1 U375 ( .A(G8GAT), .B(G15GAT), .Z(n329) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(G197GAT), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U378 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n331) );
  XNOR2_X1 U379 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n344) );
  XOR2_X1 U382 ( .A(G113GAT), .B(G1GAT), .Z(n429) );
  XOR2_X1 U383 ( .A(G141GAT), .B(G22GAT), .Z(n335) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(G50GAT), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U386 ( .A(n429), .B(n336), .Z(n338) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U389 ( .A(n339), .B(KEYINPUT66), .Z(n342) );
  XNOR2_X1 U390 ( .A(n340), .B(KEYINPUT69), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U392 ( .A(n344), .B(n343), .Z(n573) );
  INV_X1 U393 ( .A(n573), .ZN(n563) );
  NAND2_X1 U394 ( .A1(n345), .A2(n563), .ZN(n347) );
  XNOR2_X1 U395 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n365) );
  XOR2_X1 U397 ( .A(G8GAT), .B(KEYINPUT76), .Z(n383) );
  XOR2_X1 U398 ( .A(n348), .B(n383), .Z(n350) );
  XNOR2_X1 U399 ( .A(G78GAT), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n352) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U404 ( .A(n354), .B(n353), .Z(n356) );
  XOR2_X1 U405 ( .A(G22GAT), .B(G155GAT), .Z(n402) );
  XNOR2_X1 U406 ( .A(n402), .B(KEYINPUT14), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n364) );
  XOR2_X1 U408 ( .A(G71GAT), .B(G127GAT), .Z(n358) );
  XNOR2_X1 U409 ( .A(G15GAT), .B(G183GAT), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U411 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n360) );
  XNOR2_X1 U412 ( .A(G1GAT), .B(G64GAT), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U414 ( .A(n362), .B(n361), .Z(n363) );
  XOR2_X1 U415 ( .A(n364), .B(n363), .Z(n566) );
  INV_X1 U416 ( .A(n566), .ZN(n580) );
  NAND2_X1 U417 ( .A1(n365), .A2(n580), .ZN(n366) );
  NOR2_X1 U418 ( .A1(n560), .A2(n366), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n367), .B(KEYINPUT47), .ZN(n373) );
  XOR2_X1 U420 ( .A(KEYINPUT75), .B(n560), .Z(n544) );
  XOR2_X1 U421 ( .A(KEYINPUT36), .B(n544), .Z(n584) );
  NOR2_X1 U422 ( .A1(n584), .A2(n580), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n368), .B(KEYINPUT45), .ZN(n369) );
  NAND2_X1 U424 ( .A1(n369), .A2(n577), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n370), .B(KEYINPUT113), .ZN(n371) );
  NAND2_X1 U426 ( .A1(n371), .A2(n573), .ZN(n372) );
  NAND2_X1 U427 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n374), .B(KEYINPUT48), .ZN(n549) );
  XNOR2_X1 U429 ( .A(KEYINPUT79), .B(KEYINPUT17), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n375), .B(KEYINPUT18), .ZN(n376) );
  XOR2_X1 U431 ( .A(n376), .B(KEYINPUT19), .Z(n378) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G183GAT), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n444) );
  XOR2_X1 U434 ( .A(KEYINPUT94), .B(G92GAT), .Z(n380) );
  XNOR2_X1 U435 ( .A(G218GAT), .B(G204GAT), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n444), .B(n381), .ZN(n393) );
  XOR2_X1 U438 ( .A(n383), .B(n382), .Z(n391) );
  XOR2_X1 U439 ( .A(G211GAT), .B(KEYINPUT21), .Z(n385) );
  XNOR2_X1 U440 ( .A(G197GAT), .B(KEYINPUT83), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n398) );
  XOR2_X1 U442 ( .A(n386), .B(KEYINPUT93), .Z(n388) );
  NAND2_X1 U443 ( .A1(G226GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n398), .B(n389), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n524) );
  NAND2_X1 U448 ( .A1(n549), .A2(n524), .ZN(n395) );
  XOR2_X1 U449 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n397) );
  XNOR2_X1 U450 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n417) );
  XNOR2_X1 U452 ( .A(n417), .B(n398), .ZN(n406) );
  XOR2_X1 U453 ( .A(KEYINPUT82), .B(KEYINPUT23), .Z(n400) );
  XNOR2_X1 U454 ( .A(G106GAT), .B(KEYINPUT24), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U456 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U457 ( .A1(G228GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U460 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n408) );
  XNOR2_X1 U461 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U463 ( .A(n410), .B(n409), .Z(n414) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n414), .B(n413), .ZN(n479) );
  INV_X1 U466 ( .A(n479), .ZN(n415) );
  NOR2_X1 U467 ( .A1(n569), .A2(n415), .ZN(n438) );
  XNOR2_X1 U468 ( .A(G134GAT), .B(G127GAT), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n416), .B(KEYINPUT0), .ZN(n452) );
  XNOR2_X1 U470 ( .A(n452), .B(n417), .ZN(n437) );
  XOR2_X1 U471 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n419) );
  XNOR2_X1 U472 ( .A(G120GAT), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U474 ( .A(G57GAT), .B(KEYINPUT91), .Z(n421) );
  XNOR2_X1 U475 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U477 ( .A(n423), .B(n422), .Z(n435) );
  XOR2_X1 U478 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n425) );
  XNOR2_X1 U479 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n433) );
  XOR2_X1 U481 ( .A(G85GAT), .B(G148GAT), .Z(n427) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G162GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U489 ( .A(n437), .B(n436), .Z(n476) );
  NAND2_X1 U490 ( .A1(n438), .A2(n476), .ZN(n440) );
  XOR2_X1 U491 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n457) );
  XOR2_X1 U493 ( .A(KEYINPUT81), .B(KEYINPUT65), .Z(n442) );
  XNOR2_X1 U494 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n456) );
  XOR2_X1 U497 ( .A(G99GAT), .B(G190GAT), .Z(n446) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(G43GAT), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U500 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U503 ( .A(n451), .B(G176GAT), .Z(n454) );
  XNOR2_X1 U504 ( .A(n452), .B(KEYINPUT20), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U506 ( .A(n456), .B(n455), .Z(n535) );
  INV_X1 U507 ( .A(n535), .ZN(n526) );
  NAND2_X1 U508 ( .A1(n457), .A2(n526), .ZN(n458) );
  XOR2_X1 U509 ( .A(KEYINPUT122), .B(n458), .Z(n565) );
  NAND2_X1 U510 ( .A1(n538), .A2(n565), .ZN(n461) );
  XOR2_X1 U511 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n459) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n465) );
  NAND2_X1 U513 ( .A1(n544), .A2(n565), .ZN(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n462) );
  XNOR2_X1 U515 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U516 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XOR2_X1 U517 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n484) );
  NAND2_X1 U518 ( .A1(n563), .A2(n577), .ZN(n497) );
  NOR2_X1 U519 ( .A1(n544), .A2(n580), .ZN(n466) );
  XNOR2_X1 U520 ( .A(n466), .B(KEYINPUT16), .ZN(n482) );
  NAND2_X1 U521 ( .A1(n526), .A2(n524), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n467), .A2(n479), .ZN(n468) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT98), .ZN(n474) );
  XOR2_X1 U525 ( .A(n524), .B(KEYINPUT95), .Z(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT27), .B(n470), .ZN(n477) );
  NOR2_X1 U527 ( .A1(n526), .A2(n479), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT97), .B(n471), .Z(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT26), .B(n472), .ZN(n571) );
  NAND2_X1 U530 ( .A1(n477), .A2(n571), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n475), .A2(n476), .ZN(n481) );
  INV_X1 U533 ( .A(n476), .ZN(n570) );
  NAND2_X1 U534 ( .A1(n477), .A2(n570), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT96), .ZN(n551) );
  XOR2_X1 U536 ( .A(n479), .B(KEYINPUT28), .Z(n529) );
  NOR2_X1 U537 ( .A1(n551), .A2(n529), .ZN(n533) );
  NAND2_X1 U538 ( .A1(n533), .A2(n535), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n493) );
  NAND2_X1 U540 ( .A1(n482), .A2(n493), .ZN(n510) );
  NOR2_X1 U541 ( .A1(n497), .A2(n510), .ZN(n490) );
  NAND2_X1 U542 ( .A1(n490), .A2(n570), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n490), .A2(n524), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT100), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U549 ( .A1(n490), .A2(n526), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  XOR2_X1 U551 ( .A(G22GAT), .B(KEYINPUT101), .Z(n492) );
  NAND2_X1 U552 ( .A1(n490), .A2(n529), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  NAND2_X1 U554 ( .A1(n580), .A2(n493), .ZN(n494) );
  NOR2_X1 U555 ( .A1(n584), .A2(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n522) );
  NOR2_X1 U558 ( .A1(n522), .A2(n497), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT38), .ZN(n506) );
  NAND2_X1 U560 ( .A1(n506), .A2(n570), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(KEYINPUT103), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n506), .A2(n524), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n504) );
  NAND2_X1 U567 ( .A1(n526), .A2(n506), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U569 ( .A(G43GAT), .B(n505), .Z(G1330GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n508) );
  NAND2_X1 U571 ( .A1(n529), .A2(n506), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n509), .ZN(G1331GAT) );
  NAND2_X1 U574 ( .A1(n538), .A2(n573), .ZN(n521) );
  NOR2_X1 U575 ( .A1(n521), .A2(n510), .ZN(n511) );
  XOR2_X1 U576 ( .A(KEYINPUT109), .B(n511), .Z(n518) );
  NAND2_X1 U577 ( .A1(n518), .A2(n570), .ZN(n515) );
  XOR2_X1 U578 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n513) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n524), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n526), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U587 ( .A1(n518), .A2(n529), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n570), .A2(n530), .ZN(n523) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U595 ( .A1(n530), .A2(n526), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n549), .A2(n533), .ZN(n534) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n545), .A2(n563), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT114), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U606 ( .A1(n545), .A2(n538), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n541), .Z(G1341GAT) );
  NAND2_X1 U609 ( .A1(n545), .A2(n566), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n549), .A2(n571), .ZN(n550) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(n552), .Z(n561) );
  NAND2_X1 U619 ( .A1(n563), .A2(n561), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(n556), .Z(n558) );
  NAND2_X1 U625 ( .A1(n561), .A2(n345), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n566), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(G183GAT), .B(KEYINPUT123), .Z(n568) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n583) );
  NOR2_X1 U638 ( .A1(n573), .A2(n583), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n583), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n583), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

