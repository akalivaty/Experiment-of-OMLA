//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  OAI211_X1 g005(.A(KEYINPUT64), .B(KEYINPUT1), .C1(new_n189), .C2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT64), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n188), .A3(new_n190), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n200), .A2(G137), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n200), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .A4(new_n201), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n191), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT0), .A4(G128), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(new_n208), .A3(new_n201), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n199), .A2(new_n212), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT65), .B1(new_n221), .B2(KEYINPUT30), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(KEYINPUT66), .A3(new_n210), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n217), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n211), .B1(new_n195), .B2(new_n198), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(KEYINPUT30), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(G116), .B(G119), .Z(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT30), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n215), .A2(new_n216), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n210), .B2(new_n219), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n237), .B(new_n238), .C1(new_n240), .C2(new_n227), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n222), .A2(new_n229), .A3(new_n236), .A4(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n232), .B(new_n230), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n226), .A2(new_n243), .A3(new_n228), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n242), .A2(new_n244), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT31), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n242), .A2(KEYINPUT31), .A3(new_n244), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n244), .B(KEYINPUT28), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n236), .B1(new_n240), .B2(new_n227), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n250), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G472), .A2(G902), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(KEYINPUT32), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n262), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n255), .B2(new_n260), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT32), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n242), .A2(new_n244), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n259), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n272), .B(new_n273), .C1(new_n258), .C2(new_n259), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n226), .A2(new_n228), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n236), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n256), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n259), .A2(new_n273), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n274), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G472), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n267), .A2(KEYINPUT67), .A3(KEYINPUT32), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n265), .A2(new_n270), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(G234), .B2(new_n280), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT71), .A2(KEYINPUT25), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G137), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(G119), .B(G128), .Z(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT24), .B(G110), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n296));
  OAI211_X1 g110(.A(G119), .B(new_n196), .C1(new_n296), .C2(KEYINPUT23), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(G128), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT68), .B1(new_n299), .B2(G128), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n295), .B1(G110), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  INV_X1    g119(.A(G125), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G140), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(KEYINPUT69), .A3(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(KEYINPUT16), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT16), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G146), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n187), .B1(new_n311), .B2(new_n313), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(G146), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n293), .A2(new_n294), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n302), .B2(G110), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n305), .A2(new_n307), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n187), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n317), .A2(KEYINPUT70), .A3(new_n323), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n292), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n292), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n317), .B2(new_n323), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n280), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(KEYINPUT71), .A2(KEYINPUT25), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n289), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI221_X1 g147(.A(new_n280), .B1(KEYINPUT71), .B2(KEYINPUT25), .C1(new_n328), .C2(new_n330), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n287), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n328), .A2(new_n330), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n287), .A2(new_n280), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT72), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n284), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G214), .B1(G237), .B2(G902), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT80), .ZN(new_n345));
  OAI21_X1  g159(.A(G210), .B1(G237), .B2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n299), .A3(G116), .ZN(new_n349));
  OAI211_X1 g163(.A(G113), .B(new_n349), .C1(new_n234), .C2(new_n348), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT74), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G104), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT76), .B(G101), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n351), .A2(new_n356), .A3(new_n352), .A4(G104), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n352), .A2(G104), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n354), .A2(new_n355), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G104), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G107), .ZN(new_n362));
  OAI21_X1  g176(.A(G101), .B1(new_n362), .B2(new_n358), .ZN(new_n363));
  AND4_X1   g177(.A1(new_n233), .A2(new_n350), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G101), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(KEYINPUT75), .A3(G101), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n358), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(new_n357), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n243), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n364), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G122), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n239), .A2(G125), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n199), .B2(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n246), .A2(G224), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT81), .B1(new_n377), .B2(new_n378), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n377), .B2(new_n378), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  INV_X1    g201(.A(new_n378), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n236), .B1(new_n366), .B2(KEYINPUT4), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT75), .B1(new_n365), .B2(G101), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n389), .B1(new_n392), .B2(new_n370), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n387), .B(new_n388), .C1(new_n393), .C2(new_n364), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n384), .A2(new_n386), .A3(new_n397), .A4(new_n394), .ZN(new_n398));
  AOI211_X1 g212(.A(new_n379), .B(new_n383), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n378), .B(KEYINPUT8), .ZN(new_n400));
  INV_X1    g214(.A(new_n364), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n360), .A2(new_n363), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n350), .A2(new_n233), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n400), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n377), .A2(new_n378), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n382), .A2(KEYINPUT7), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n381), .B(new_n409), .Z(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n280), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n347), .B1(new_n399), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n396), .A2(new_n398), .ZN(new_n414));
  INV_X1    g228(.A(new_n379), .ZN(new_n415));
  INV_X1    g229(.A(new_n383), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n412), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n346), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n345), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT9), .B(G234), .ZN(new_n421));
  OAI21_X1  g235(.A(G221), .B1(new_n421), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n224), .A2(new_n225), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n239), .B1(new_n375), .B2(new_n372), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n360), .A2(new_n363), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n371), .A2(new_n425), .B1(new_n199), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT77), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n198), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n432));
  OAI21_X1  g246(.A(G128), .B1(new_n432), .B2(KEYINPUT78), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT1), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(G143), .B2(new_n187), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT78), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n191), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n426), .B1(new_n431), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n439), .A2(KEYINPUT79), .A3(KEYINPUT10), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n196), .B1(new_n435), .B2(new_n436), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(KEYINPUT78), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n442), .A2(new_n443), .B1(new_n188), .B2(new_n190), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n198), .B(KEYINPUT77), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n403), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n441), .B1(new_n446), .B2(new_n427), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n424), .B(new_n429), .C1(new_n440), .C2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G140), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n246), .A2(G227), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n429), .B1(new_n440), .B2(new_n447), .ZN(new_n453));
  INV_X1    g267(.A(new_n424), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n199), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n426), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n424), .B1(new_n457), .B2(new_n446), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n439), .B1(new_n456), .B2(new_n426), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n220), .A2(KEYINPUT12), .ZN(new_n460));
  OAI22_X1  g274(.A1(new_n458), .A2(KEYINPUT12), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n448), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n451), .B(KEYINPUT73), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n452), .A2(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G469), .B1(new_n464), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(G469), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n451), .B1(new_n455), .B2(new_n448), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n461), .A2(new_n448), .A3(new_n451), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n466), .B(new_n280), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n423), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G475), .ZN(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n361), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n245), .A2(new_n246), .A3(G214), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n189), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n245), .A2(new_n246), .A3(G143), .A4(G214), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT17), .A3(G131), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(G131), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n475), .A2(new_n209), .A3(new_n476), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n483), .A2(KEYINPUT17), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n315), .A2(new_n316), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(KEYINPUT18), .A2(G131), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n476), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n309), .A2(G146), .A3(new_n310), .ZN(new_n491));
  INV_X1    g305(.A(new_n487), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n491), .A2(new_n322), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n473), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n486), .A2(new_n473), .A3(new_n494), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n471), .B1(new_n498), .B2(new_n280), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n309), .B2(new_n310), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n321), .A2(KEYINPUT19), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n318), .B(new_n483), .C1(G146), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n494), .A3(KEYINPUT85), .ZN(new_n505));
  INV_X1    g319(.A(new_n473), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT85), .B1(new_n504), .B2(new_n494), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n494), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT85), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n506), .A3(new_n505), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n512), .B1(new_n516), .B2(new_n497), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n511), .B1(new_n517), .B2(KEYINPUT20), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT20), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n509), .A2(new_n512), .A3(new_n519), .A4(new_n510), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n499), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT21), .B(G898), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT92), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(G234), .A2(G237), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n525), .A2(G902), .A3(G953), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n525), .A2(G952), .A3(new_n246), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n421), .A2(new_n285), .A3(G953), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n189), .A2(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n196), .A2(G143), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n200), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n536), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G116), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G122), .ZN(new_n541));
  INV_X1    g355(.A(G122), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n542), .A2(KEYINPUT88), .A3(G116), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT88), .B1(new_n542), .B2(G116), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G107), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n352), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n539), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n536), .A2(G134), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n535), .A2(new_n200), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n541), .A2(KEYINPUT14), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n543), .A2(new_n544), .B1(KEYINPUT14), .B2(new_n541), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n559), .B2(G107), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n532), .B1(new_n550), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n554), .B(KEYINPUT89), .ZN(new_n562));
  OAI21_X1  g376(.A(G107), .B1(new_n562), .B2(new_n557), .ZN(new_n563));
  INV_X1    g377(.A(new_n553), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n565), .A2(KEYINPUT90), .A3(new_n549), .A4(new_n531), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n563), .A2(new_n564), .B1(new_n548), .B2(new_n539), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT90), .B1(new_n568), .B2(new_n531), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n280), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n568), .A2(new_n531), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n561), .A3(new_n566), .ZN(new_n581));
  INV_X1    g395(.A(new_n576), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n280), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n521), .A2(new_n530), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n420), .A2(new_n470), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n343), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(new_n355), .ZN(G3));
  NAND2_X1  g404(.A1(new_n518), .A2(new_n520), .ZN(new_n591));
  INV_X1    g405(.A(new_n497), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n280), .B1(new_n592), .B2(new_n495), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G475), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n581), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n561), .A2(new_n578), .A3(KEYINPUT33), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n597), .A2(G478), .A3(new_n280), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n570), .A2(new_n571), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT93), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT93), .B1(new_n570), .B2(new_n571), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n529), .B2(new_n527), .ZN(new_n606));
  INV_X1    g420(.A(new_n344), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n413), .B2(new_n419), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(G469), .A2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n462), .A2(new_n463), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n455), .A2(new_n448), .A3(new_n451), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(G469), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n469), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n422), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n253), .A2(new_n254), .B1(new_n258), .B2(new_n259), .ZN(new_n617));
  OAI21_X1  g431(.A(G472), .B1(new_n617), .B2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n268), .A2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n341), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  XOR2_X1   g437(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n624));
  NAND3_X1  g438(.A1(new_n509), .A2(new_n510), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n509), .B2(new_n510), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n584), .B(new_n594), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n530), .B(KEYINPUT95), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n620), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n292), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT97), .Z(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n327), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT70), .B1(new_n317), .B2(new_n323), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n326), .A2(new_n327), .A3(new_n640), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n339), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT98), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n645), .A3(new_n648), .A4(new_n339), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n615), .B(new_n422), .C1(new_n335), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n619), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n420), .A3(new_n587), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT37), .B(G110), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT99), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n526), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n529), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n628), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n399), .A2(new_n412), .A3(new_n347), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n346), .B1(new_n417), .B2(new_n418), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n661), .B(new_n344), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT67), .B1(new_n267), .B2(KEYINPUT32), .ZN(new_n666));
  NOR4_X1   g480(.A1(new_n617), .A2(new_n264), .A3(new_n269), .A4(new_n266), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n268), .A2(new_n269), .B1(new_n281), .B2(G472), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n651), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n608), .A2(new_n671), .A3(new_n661), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n665), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n196), .ZN(G30));
  XNOR2_X1  g488(.A(new_n659), .B(KEYINPUT39), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n470), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT40), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n333), .A2(new_n334), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n650), .B1(new_n679), .B2(new_n286), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n521), .A2(new_n585), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n680), .A2(new_n681), .A3(new_n344), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n677), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n413), .A2(new_n419), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT38), .Z(new_n685));
  AND2_X1   g499(.A1(new_n276), .A2(new_n244), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n251), .B1(new_n250), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n280), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n268), .A2(new_n269), .B1(new_n688), .B2(G472), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n668), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  OR3_X1    g505(.A1(new_n683), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  INV_X1    g507(.A(new_n651), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n595), .A2(new_n604), .A3(new_n659), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n284), .A2(new_n694), .A3(new_n608), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  OAI21_X1  g512(.A(new_n280), .B1(new_n467), .B2(new_n468), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G469), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n469), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n423), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n284), .A2(new_n342), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n610), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n633), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NOR2_X1   g523(.A1(new_n586), .A2(new_n680), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n284), .A2(new_n710), .A3(new_n608), .A4(new_n702), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  OAI211_X1 g530(.A(new_n681), .B(new_n344), .C1(new_n662), .C2(new_n663), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n608), .A2(new_n719), .A3(new_n681), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n255), .B1(new_n250), .B2(new_n277), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n262), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n618), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AND4_X1   g539(.A1(new_n342), .A2(new_n702), .A3(new_n629), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n721), .A2(new_n726), .A3(KEYINPUT103), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NOR2_X1   g546(.A1(new_n724), .A2(new_n680), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(new_n608), .A3(new_n696), .A4(new_n702), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  INV_X1    g549(.A(new_n343), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n413), .A2(new_n419), .A3(new_n344), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n616), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n695), .A2(KEYINPUT42), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n341), .B1(new_n669), .B2(new_n263), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n738), .A3(new_n696), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND4_X1  g559(.A1(new_n738), .A2(new_n284), .A3(new_n342), .A4(new_n661), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  NAND2_X1  g561(.A1(new_n464), .A2(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n612), .A2(new_n613), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n751), .A3(G469), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n752), .B2(new_n611), .ZN(new_n753));
  INV_X1    g567(.A(new_n469), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n611), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n423), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n675), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT104), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT43), .B1(new_n521), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n521), .A2(new_n604), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n680), .B1(new_n268), .B2(new_n618), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT44), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(KEYINPUT44), .A3(new_n763), .ZN(new_n766));
  INV_X1    g580(.A(new_n737), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n757), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT106), .Z(new_n772));
  NAND2_X1  g586(.A1(new_n757), .A2(new_n770), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT105), .Z(new_n774));
  AND2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n284), .A2(new_n342), .A3(new_n737), .A4(new_n695), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  NOR4_X1   g592(.A1(new_n341), .A2(new_n761), .A3(new_n423), .A4(new_n345), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n701), .B(KEYINPUT49), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n779), .B2(new_n780), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n783), .A3(new_n691), .A4(new_n685), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n737), .A2(new_n423), .A3(new_n701), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT115), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(KEYINPUT115), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n787), .A3(new_n529), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n342), .A3(new_n691), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n595), .A3(new_n604), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n741), .A3(new_n762), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT48), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n246), .A2(G952), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n342), .A2(new_n762), .A3(new_n528), .A4(new_n725), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n608), .A2(new_n702), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n793), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT118), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n793), .A2(new_n802), .A3(new_n795), .A4(new_n799), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n797), .A2(new_n767), .ZN(new_n806));
  INV_X1    g620(.A(new_n775), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n701), .A2(new_n422), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT114), .Z(new_n809));
  AOI21_X1  g623(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n595), .A2(new_n604), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n791), .A2(new_n792), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n788), .A2(new_n733), .A3(new_n762), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n797), .A2(new_n607), .A3(new_n685), .A4(new_n702), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n805), .B1(new_n810), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT117), .B1(new_n775), .B2(new_n808), .ZN(new_n821));
  INV_X1    g635(.A(new_n806), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n775), .A2(KEYINPUT117), .A3(new_n808), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n804), .B(new_n820), .C1(new_n825), .C2(new_n819), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n284), .B(new_n694), .C1(new_n664), .C2(KEYINPUT100), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n671), .B1(new_n608), .B2(new_n661), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n697), .B(new_n734), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n659), .B(KEYINPUT110), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n470), .A2(new_n680), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n668), .B2(new_n689), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n719), .B1(new_n608), .B2(new_n681), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n721), .A2(KEYINPUT111), .A3(new_n832), .ZN(new_n838));
  AOI211_X1 g652(.A(KEYINPUT52), .B(new_n829), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n838), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n697), .A2(new_n734), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n673), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n605), .B1(new_n595), .B2(new_n585), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n620), .A2(new_n420), .A3(new_n629), .A4(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n653), .C1(new_n343), .C2(new_n588), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n627), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n499), .B1(new_n850), .B2(new_n625), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT108), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n584), .A2(new_n660), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n284), .A2(new_n767), .A3(new_n856), .A4(new_n694), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n695), .A2(new_n724), .A3(new_n680), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n738), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n746), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT109), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n737), .A2(new_n854), .A3(new_n855), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n863), .A2(new_n670), .B1(new_n738), .B2(new_n858), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT109), .B1(new_n864), .B2(new_n746), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n849), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n703), .B1(new_n609), .B2(new_n632), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n713), .B2(new_n714), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n731), .A2(new_n870), .A3(new_n744), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT112), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n731), .A2(new_n870), .A3(new_n744), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n845), .A2(new_n868), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  INV_X1    g690(.A(new_n838), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT111), .B1(new_n721), .B2(new_n832), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n843), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n841), .A2(new_n840), .A3(new_n843), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n860), .A2(new_n861), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n864), .A2(KEYINPUT109), .A3(new_n746), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n848), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n731), .A3(new_n744), .A4(new_n870), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n867), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n875), .A2(new_n876), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n871), .A2(new_n866), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n876), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT113), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT113), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n875), .A2(new_n887), .A3(new_n876), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n887), .A2(new_n890), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n876), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n826), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n784), .B1(new_n897), .B2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n379), .B1(new_n396), .B2(new_n398), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n416), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n280), .B1(new_n875), .B2(new_n887), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(G210), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n902), .B1(new_n904), .B2(KEYINPUT56), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n246), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n903), .A2(KEYINPUT119), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n903), .A2(KEYINPUT119), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n347), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G51));
  NAND2_X1  g727(.A1(new_n872), .A2(new_n874), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n880), .A2(KEYINPUT53), .A3(new_n881), .A4(new_n885), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n845), .B2(new_n889), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT54), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n894), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n611), .B(KEYINPUT57), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n920), .A2(new_n921), .B1(new_n467), .B2(new_n468), .ZN(new_n922));
  INV_X1    g736(.A(new_n752), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n909), .A2(new_n923), .A3(new_n910), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n906), .B1(new_n922), .B2(new_n924), .ZN(G54));
  AND2_X1   g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n909), .A2(new_n910), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n497), .A3(new_n516), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n909), .A2(new_n509), .A3(new_n910), .A4(new_n926), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n928), .A2(new_n907), .A3(new_n929), .ZN(G60));
  AND2_X1   g744(.A1(new_n597), .A2(new_n598), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n876), .B1(new_n875), .B2(new_n887), .ZN(new_n936));
  OAI211_X1 g750(.A(KEYINPUT120), .B(new_n935), .C1(new_n888), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n907), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT120), .B1(new_n919), .B2(new_n935), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT121), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n935), .B1(new_n888), .B2(new_n936), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n943), .A2(new_n944), .A3(new_n907), .A4(new_n937), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n892), .A2(new_n896), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n932), .B1(new_n946), .B2(new_n934), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n940), .A2(new_n945), .A3(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n875), .B2(new_n887), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n951), .A2(new_n645), .A3(new_n644), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n907), .B1(new_n951), .B2(new_n337), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  OAI22_X1  g768(.A1(new_n952), .A2(new_n953), .B1(KEYINPUT122), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G66));
  AOI21_X1  g771(.A(new_n246), .B1(new_n523), .B2(G224), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n731), .A2(new_n870), .A3(new_n849), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n246), .ZN(new_n960));
  INV_X1    g774(.A(G898), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n900), .B1(new_n961), .B2(G953), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  NAND4_X1  g777(.A1(new_n721), .A2(new_n757), .A3(new_n675), .A4(new_n741), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n744), .A2(new_n843), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n746), .A2(new_n768), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n777), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n246), .A2(G900), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n967), .B2(new_n971), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n222), .A2(new_n229), .A3(new_n241), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(new_n503), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n692), .A2(new_n843), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n981));
  INV_X1    g795(.A(new_n676), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n736), .A2(new_n982), .A3(new_n767), .A4(new_n846), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n768), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n777), .A2(new_n980), .A3(new_n981), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n246), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n978), .B1(new_n986), .B2(new_n975), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n977), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n977), .B2(new_n987), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(G72));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT126), .Z(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n985), .B2(new_n959), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n271), .B(KEYINPUT127), .Z(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n250), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n887), .A2(new_n890), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n272), .A2(new_n251), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n998), .A2(new_n993), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n777), .A2(new_n966), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n994), .B1(new_n1001), .B2(new_n959), .ZN(new_n1002));
  INV_X1    g816(.A(new_n996), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1002), .A2(new_n259), .A3(new_n1003), .ZN(new_n1004));
  AND4_X1   g818(.A1(new_n907), .A2(new_n997), .A3(new_n1000), .A4(new_n1004), .ZN(G57));
endmodule


