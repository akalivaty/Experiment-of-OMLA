//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT66), .B(G131), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT11), .A2(G134), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT11), .A2(G134), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT64), .A2(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(new_n190), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n190), .A3(KEYINPUT65), .A4(new_n195), .ZN(new_n199));
  AOI211_X1 g013(.A(new_n189), .B(new_n193), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G128), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n202), .B(new_n204), .C1(KEYINPUT1), .C2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT64), .A2(G137), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT64), .A2(G137), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n210), .A2(new_n211), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n213), .B2(new_n192), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n207), .B(new_n209), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n200), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT0), .A4(G128), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n202), .A2(new_n204), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G128), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n193), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n210), .A2(new_n211), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT65), .B1(new_n222), .B2(new_n190), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT11), .A2(G134), .ZN(new_n224));
  NOR4_X1   g038(.A1(new_n210), .A2(new_n211), .A3(new_n224), .A4(new_n197), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n198), .A2(new_n199), .ZN(new_n228));
  INV_X1    g042(.A(new_n189), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n221), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n220), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n216), .B1(new_n231), .B2(KEYINPUT67), .ZN(new_n232));
  INV_X1    g046(.A(new_n220), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n228), .B2(new_n221), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n235), .B2(new_n200), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n188), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT2), .A2(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(KEYINPUT2), .B2(G113), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n241), .A2(new_n243), .B1(KEYINPUT2), .B2(G113), .ZN(new_n244));
  XNOR2_X1  g058(.A(G116), .B(G119), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(new_n245), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n200), .A2(new_n215), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n227), .A2(new_n230), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n220), .B(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT30), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(new_n248), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n248), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G210), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n260), .B(KEYINPUT27), .Z(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n261), .B(new_n262), .Z(new_n263));
  NAND3_X1  g077(.A1(new_n255), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT31), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n255), .A2(KEYINPUT31), .A3(new_n257), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n263), .B(KEYINPUT70), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n249), .B1(new_n236), .B2(new_n237), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n256), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI211_X1 g088(.A(new_n248), .B(new_n249), .C1(new_n250), .C2(new_n252), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT28), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n256), .B1(new_n253), .B2(KEYINPUT72), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n279));
  AOI211_X1 g093(.A(new_n279), .B(new_n249), .C1(new_n250), .C2(new_n252), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n271), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n248), .B1(new_n232), .B2(new_n238), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n257), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT71), .B1(new_n284), .B2(KEYINPUT28), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n270), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n268), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n268), .B2(new_n286), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT74), .B(new_n187), .C1(new_n288), .C2(new_n289), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n187), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n268), .A2(new_n286), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n268), .A2(new_n286), .A3(new_n287), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n253), .A2(new_n256), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT28), .B1(new_n301), .B2(new_n275), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n281), .A2(new_n302), .A3(KEYINPUT29), .A4(new_n263), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT76), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n276), .A2(new_n281), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT71), .ZN(new_n308));
  INV_X1    g122(.A(new_n285), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT75), .A4(new_n269), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n255), .A2(new_n257), .ZN(new_n312));
  INV_X1    g126(.A(new_n263), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n282), .A2(new_n285), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT75), .B1(new_n316), .B2(new_n269), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n306), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n300), .A2(KEYINPUT32), .B1(new_n318), .B2(G472), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n295), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(G234), .B2(new_n304), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT22), .B(G137), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT81), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT82), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n208), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT24), .B(G110), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n333), .B2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n334), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(G110), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G140), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(KEYINPUT77), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(G125), .A3(G140), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT16), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n350), .B2(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G146), .ZN(new_n358));
  XNOR2_X1  g172(.A(G125), .B(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n201), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n348), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n201), .A3(new_n356), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n344), .A2(G110), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(new_n336), .C2(new_n337), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT80), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n368), .A3(new_n365), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n332), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n330), .A2(new_n331), .B1(new_n361), .B2(new_n365), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT83), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n332), .ZN(new_n373));
  INV_X1    g187(.A(new_n369), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n368), .B1(new_n361), .B2(new_n365), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n377));
  INV_X1    g191(.A(new_n371), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n324), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n304), .B1(new_n370), .B2(new_n371), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT25), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT25), .B(new_n304), .C1(new_n370), .C2(new_n371), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n380), .B1(new_n385), .B2(new_n322), .ZN(new_n386));
  OR2_X1    g200(.A1(G475), .A2(G902), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT20), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n258), .A2(new_n259), .A3(G214), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n203), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n189), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n390), .B(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n229), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n351), .A2(new_n353), .ZN(new_n396));
  MUX2_X1   g210(.A(new_n359), .B(new_n396), .S(KEYINPUT19), .Z(new_n397));
  OAI211_X1 g211(.A(new_n395), .B(new_n358), .C1(new_n397), .C2(G146), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(G146), .ZN(new_n399));
  NAND3_X1  g213(.A1(KEYINPUT91), .A2(KEYINPUT18), .A3(G131), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n399), .A2(new_n360), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n393), .A2(new_n400), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(G113), .B(G122), .Z(new_n405));
  XOR2_X1   g219(.A(KEYINPUT92), .B(G104), .Z(new_n406));
  XOR2_X1   g220(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n392), .A2(new_n394), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n189), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n362), .A3(new_n358), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n403), .A3(new_n407), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n389), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n415), .A2(KEYINPUT94), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(KEYINPUT94), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n418));
  INV_X1    g232(.A(new_n414), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n407), .B1(new_n398), .B2(new_n403), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n409), .A2(KEYINPUT93), .A3(new_n414), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n387), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n416), .B(new_n417), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n392), .A2(new_n394), .A3(new_n410), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n412), .A2(new_n362), .A3(new_n358), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n403), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n407), .B1(new_n428), .B2(KEYINPUT95), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n413), .A2(new_n430), .A3(new_n403), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(KEYINPUT96), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n414), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT96), .B1(new_n429), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n304), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G475), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n208), .A2(G143), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n203), .A2(G128), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n213), .A3(new_n440), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n441), .A2(KEYINPUT98), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(KEYINPUT98), .ZN(new_n443));
  XNOR2_X1  g257(.A(G116), .B(G122), .ZN(new_n444));
  INV_X1    g258(.A(G107), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n439), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n440), .B(KEYINPUT13), .Z(new_n448));
  OAI21_X1  g262(.A(G134), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n442), .A2(new_n443), .A3(new_n446), .A4(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G122), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G116), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n445), .B1(new_n452), .B2(KEYINPUT14), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n444), .ZN(new_n454));
  INV_X1    g268(.A(new_n441), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n213), .B1(new_n439), .B2(new_n440), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n458), .A2(new_n321), .A3(G953), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n450), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n450), .B2(new_n457), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n304), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G478), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT99), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n468), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n304), .B(new_n470), .C1(new_n460), .C2(new_n461), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G952), .ZN(new_n473));
  AOI211_X1 g287(.A(G953), .B(new_n473), .C1(G234), .C2(G237), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT21), .B(G898), .Z(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT100), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n304), .B(new_n259), .C1(G234), .C2(G237), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n425), .A2(new_n436), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G140), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT84), .ZN(new_n483));
  INV_X1    g297(.A(G227), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G953), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n483), .B(new_n485), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G104), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n488), .A2(KEYINPUT3), .A3(G107), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n445), .A2(G104), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT3), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(G107), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G101), .ZN(new_n494));
  INV_X1    g308(.A(G101), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n489), .A2(new_n491), .A3(new_n495), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(KEYINPUT4), .A3(new_n496), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n252), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n490), .A2(new_n492), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G101), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(KEYINPUT85), .A3(G101), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n207), .A2(new_n209), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT10), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT86), .B1(new_n507), .B2(KEYINPUT10), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT10), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n511), .B(new_n512), .C1(new_n505), .C2(new_n506), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n250), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n515), .B1(new_n509), .B2(new_n514), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n487), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n505), .A2(new_n506), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n507), .B2(KEYINPUT87), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT87), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n505), .A2(new_n521), .A3(new_n506), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n250), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT12), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n527), .A3(new_n250), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n486), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n518), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G469), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n304), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n304), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OR3_X1    g348(.A1(new_n516), .A2(new_n517), .A3(new_n487), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n487), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n537), .A3(G469), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G214), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G210), .B1(G237), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n248), .A2(new_n497), .A3(new_n498), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n333), .A2(G116), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n545), .B(G113), .C1(KEYINPUT5), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n244), .A2(new_n245), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n549), .A2(new_n505), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G110), .B(G122), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n544), .A2(new_n552), .A3(new_n550), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(KEYINPUT6), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n506), .A2(new_n350), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n220), .A2(G125), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n259), .A2(G224), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT88), .Z(new_n561));
  XNOR2_X1  g375(.A(new_n559), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n563), .A3(new_n553), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n556), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  OR3_X1    g379(.A1(new_n549), .A2(new_n505), .A3(KEYINPUT89), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n549), .A2(new_n505), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT89), .B1(new_n549), .B2(new_n505), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n552), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT90), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n558), .A2(new_n573), .B1(KEYINPUT7), .B2(new_n560), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(new_n559), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n559), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n555), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n304), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n543), .B1(new_n565), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n577), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n580), .B2(new_n571), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n556), .A2(new_n562), .A3(new_n564), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n542), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n541), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G221), .ZN(new_n585));
  INV_X1    g399(.A(new_n458), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(new_n304), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n481), .A2(new_n539), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n320), .A2(new_n386), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND3_X1  g406(.A1(new_n386), .A2(new_n588), .A3(new_n539), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n304), .B1(new_n288), .B2(new_n289), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(G472), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n462), .A2(new_n463), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n460), .B2(new_n461), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n304), .A2(G478), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n596), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n425), .A2(new_n436), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n479), .ZN(new_n606));
  INV_X1    g420(.A(new_n583), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n542), .B1(new_n581), .B2(new_n582), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n540), .B(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n595), .A2(new_n292), .A3(new_n294), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  AND2_X1   g427(.A1(new_n292), .A2(new_n294), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n421), .A2(new_n422), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT102), .B1(new_n615), .B2(new_n388), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n388), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n424), .B2(new_n423), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n618), .B2(KEYINPUT102), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n436), .A2(new_n472), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n609), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n595), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NAND2_X1  g438(.A1(new_n594), .A2(G472), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n332), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(KEYINPUT103), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(KEYINPUT103), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OAI22_X1  g444(.A1(new_n628), .A2(new_n630), .B1(new_n375), .B2(new_n374), .ZN(new_n631));
  INV_X1    g445(.A(new_n628), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n632), .A2(new_n367), .A3(new_n369), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n323), .A2(new_n634), .B1(new_n385), .B2(new_n322), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n589), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n292), .A2(new_n625), .A3(new_n636), .A4(new_n294), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(new_n635), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n641), .A2(new_n584), .A3(new_n588), .A4(new_n539), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n295), .B2(new_n319), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n474), .B1(new_n478), .B2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n619), .A2(new_n620), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  OAI211_X1 g462(.A(KEYINPUT32), .B(new_n187), .C1(new_n288), .C2(new_n289), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n270), .B1(new_n275), .B2(new_n301), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n264), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n304), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G472), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n295), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n645), .B(KEYINPUT39), .Z(new_n655));
  NAND3_X1  g469(.A1(new_n539), .A2(new_n588), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n579), .A2(new_n583), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT38), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n540), .A3(new_n635), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n604), .A2(new_n472), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n654), .A2(new_n657), .A3(new_n658), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NOR2_X1   g479(.A1(new_n605), .A2(new_n645), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n643), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G146), .ZN(G48));
  NAND2_X1  g482(.A1(new_n530), .A2(new_n304), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G469), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(KEYINPUT105), .A3(new_n532), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(new_n672), .A3(G469), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n587), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n610), .A3(new_n386), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n295), .B2(new_n319), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT41), .B(G113), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  INV_X1    g492(.A(new_n674), .ZN(new_n679));
  INV_X1    g493(.A(new_n386), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n320), .A2(new_n621), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  INV_X1    g497(.A(new_n481), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n635), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n674), .A3(new_n584), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n320), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  XNOR2_X1  g503(.A(KEYINPUT106), .B(G472), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n594), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n268), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n269), .B1(new_n281), .B2(new_n302), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n187), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n386), .A3(new_n694), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n541), .B(new_n479), .C1(new_n579), .C2(new_n583), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n674), .A2(new_n604), .A3(new_n472), .A4(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT107), .B(G122), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G24));
  NAND3_X1  g514(.A1(new_n691), .A2(new_n641), .A3(new_n694), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n674), .A2(new_n666), .A3(new_n584), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n350), .ZN(G27));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n535), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n535), .A2(new_n537), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n532), .B(new_n534), .C1(new_n708), .C2(new_n531), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n588), .A2(new_n540), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n659), .A2(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n666), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n680), .B1(new_n295), .B2(new_n319), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n318), .A2(G472), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n649), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n300), .A2(KEYINPUT32), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n386), .B(new_n712), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n714), .A2(new_n715), .B1(new_n719), .B2(KEYINPUT42), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G131), .ZN(G33));
  AND2_X1   g535(.A1(new_n709), .A2(new_n711), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n646), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  NAND2_X1  g538(.A1(new_n614), .A2(new_n625), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n603), .A2(new_n436), .A3(new_n425), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n641), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n659), .A2(new_n541), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n708), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n707), .B2(KEYINPUT45), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n533), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n532), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n588), .B(new_n655), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G137), .ZN(G39));
  OR2_X1    g558(.A1(new_n739), .A2(new_n740), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n588), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(KEYINPUT47), .B(new_n588), .C1(new_n739), .C2(new_n740), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n320), .ZN(new_n751));
  INV_X1    g565(.A(new_n733), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n752), .A2(new_n605), .A3(new_n386), .A4(new_n645), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  NAND2_X1  g569(.A1(new_n728), .A2(new_n674), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n733), .A2(new_n474), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT119), .ZN(new_n759));
  INV_X1    g573(.A(new_n718), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n680), .B1(new_n760), .B2(new_n319), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n763));
  AOI211_X1 g577(.A(new_n473), .B(G953), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n762), .A2(KEYINPUT121), .A3(KEYINPUT48), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n691), .A2(new_n386), .A3(new_n694), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(new_n474), .A3(new_n728), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n584), .A3(new_n674), .ZN(new_n768));
  OR4_X1    g582(.A1(new_n680), .A2(new_n654), .A3(new_n679), .A4(new_n757), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(new_n605), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n764), .A2(new_n765), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n767), .A2(new_n733), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n750), .A2(KEYINPUT116), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT47), .B1(new_n745), .B2(new_n588), .ZN(new_n774));
  INV_X1    g588(.A(new_n749), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT116), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n671), .A2(new_n673), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT117), .Z(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n588), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n772), .B1(new_n773), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT118), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n772), .C1(new_n773), .C2(new_n781), .ZN(new_n785));
  INV_X1    g599(.A(new_n701), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n759), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n603), .A2(new_n604), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n769), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n756), .A2(new_n540), .A3(new_n660), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n474), .A3(new_n766), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT50), .Z(new_n793));
  AND2_X1   g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n783), .A2(new_n785), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n772), .B1(new_n750), .B2(new_n779), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n789), .A2(KEYINPUT120), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n793), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n789), .A2(KEYINPUT120), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT51), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n771), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n425), .A2(new_n436), .A3(new_n472), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n696), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n425), .A2(new_n436), .A3(new_n472), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n609), .A2(new_n806), .A3(KEYINPUT110), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n595), .A2(new_n292), .A3(new_n294), .A4(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n611), .A2(new_n809), .A3(new_n637), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n591), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n680), .B(new_n589), .C1(new_n295), .C2(new_n319), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n611), .A2(new_n809), .A3(new_n637), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT111), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n674), .A2(new_n386), .A3(new_n621), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n295), .A2(new_n319), .B1(new_n817), .B2(new_n686), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n676), .A3(new_n698), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n472), .A2(new_n645), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n733), .A2(new_n436), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n539), .A2(new_n588), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n821), .A2(new_n635), .A3(new_n822), .A4(new_n619), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n320), .A2(new_n823), .B1(new_n786), .B2(new_n712), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n819), .A2(new_n720), .A3(new_n723), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n802), .B1(new_n816), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n720), .A2(new_n723), .A3(new_n824), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n812), .A2(new_n815), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT112), .A4(new_n819), .ZN(new_n829));
  INV_X1    g643(.A(new_n645), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n587), .B1(new_n830), .B2(KEYINPUT114), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(KEYINPUT114), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n641), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n584), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n662), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n833), .A2(new_n709), .A3(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n643), .A2(new_n666), .B1(new_n654), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n703), .B1(new_n643), .B2(new_n646), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n826), .A2(new_n829), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n838), .A2(new_n845), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n837), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n840), .B1(new_n848), .B2(KEYINPUT52), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n826), .A4(new_n829), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n844), .A2(new_n851), .A3(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n843), .A2(new_n850), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n854));
  INV_X1    g668(.A(new_n675), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n320), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n695), .A2(new_n697), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n854), .B1(new_n858), .B2(new_n818), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n676), .A2(new_n698), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(KEYINPUT115), .A3(new_n682), .A4(new_n688), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n714), .A2(new_n715), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT53), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n824), .A2(new_n723), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n862), .A2(new_n828), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n849), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n801), .B(new_n852), .C1(KEYINPUT54), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n473), .A2(new_n259), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n680), .A2(new_n710), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n660), .B(new_n726), .C1(new_n875), .C2(KEYINPUT109), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(KEYINPUT109), .B2(new_n875), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n777), .B(KEYINPUT49), .Z(new_n878));
  OR3_X1    g692(.A1(new_n877), .A2(new_n654), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n556), .A2(new_n564), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n562), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  AND3_X1   g697(.A1(new_n870), .A2(G210), .A3(G902), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(KEYINPUT56), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n259), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n884), .A2(KEYINPUT56), .A3(new_n883), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(G51));
  XNOR2_X1  g704(.A(new_n533), .B(KEYINPUT57), .ZN(new_n891));
  AOI221_X4 g705(.A(KEYINPUT54), .B1(new_n849), .B2(new_n868), .C1(new_n843), .C2(new_n850), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n853), .B2(new_n869), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(KEYINPUT122), .B(new_n891), .C1(new_n892), .C2(new_n894), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n530), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n870), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n304), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n737), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n886), .B1(new_n899), .B2(new_n902), .ZN(G54));
  AND2_X1   g717(.A1(KEYINPUT58), .A2(G475), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n901), .A2(new_n615), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n615), .B1(new_n901), .B2(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n886), .ZN(G60));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT59), .Z(new_n909));
  NOR2_X1   g723(.A1(new_n601), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n892), .B2(new_n894), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n911), .A2(KEYINPUT123), .A3(new_n887), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT123), .B1(new_n911), .B2(new_n887), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n852), .B1(new_n870), .B2(KEYINPUT54), .ZN(new_n914));
  INV_X1    g728(.A(new_n909), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n600), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n912), .A2(new_n913), .A3(new_n916), .ZN(G63));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n372), .A2(new_n379), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n900), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n887), .ZN(new_n924));
  INV_X1    g738(.A(new_n634), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n900), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n918), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n926), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n887), .A4(new_n923), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(G66));
  INV_X1    g744(.A(G224), .ZN(new_n931));
  OAI21_X1  g745(.A(G953), .B1(new_n477), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n828), .A2(new_n819), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n881), .B1(G898), .B2(new_n259), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G69));
  NAND2_X1  g750(.A1(new_n239), .A2(new_n254), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT124), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n397), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n846), .A2(new_n847), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n664), .A3(new_n667), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n752), .B(new_n656), .C1(new_n605), .C2(new_n806), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n715), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n774), .A2(new_n775), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n751), .A2(new_n753), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n743), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n259), .B1(new_n941), .B2(KEYINPUT62), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n939), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n484), .A2(G900), .A3(G953), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n742), .A2(new_n761), .A3(new_n835), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n754), .A2(new_n720), .A3(new_n723), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n940), .A2(new_n667), .A3(new_n743), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n955), .B1(new_n962), .B2(G953), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n954), .B1(new_n939), .B2(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  OAI21_X1  g780(.A(new_n933), .B1(new_n941), .B2(KEYINPUT62), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n950), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n312), .B(KEYINPUT126), .Z(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n263), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n966), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n962), .B2(new_n933), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n969), .A2(new_n263), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n970), .B(new_n887), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n314), .B2(new_n264), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n844), .A2(new_n851), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(G57));
endmodule


