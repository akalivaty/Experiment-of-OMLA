

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U556 ( .A(n711), .B(n710), .ZN(n718) );
  XNOR2_X1 U557 ( .A(n740), .B(KEYINPUT32), .ZN(n746) );
  NOR2_X1 U558 ( .A1(n749), .A2(n780), .ZN(n526) );
  OR2_X1 U559 ( .A1(n745), .A2(n744), .ZN(n527) );
  OR2_X1 U560 ( .A1(n745), .A2(n720), .ZN(n721) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n710) );
  XNOR2_X1 U562 ( .A(KEYINPUT31), .B(KEYINPUT93), .ZN(n729) );
  XNOR2_X1 U563 ( .A(n730), .B(n729), .ZN(n731) );
  AND2_X1 U564 ( .A1(n746), .A2(n527), .ZN(n783) );
  NAND2_X1 U565 ( .A1(n773), .A2(n771), .ZN(n733) );
  NAND2_X1 U566 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U567 ( .A1(G164), .A2(G1384), .ZN(n773) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n635) );
  NOR2_X1 U569 ( .A1(G651), .A2(n635), .ZN(n650) );
  INV_X1 U570 ( .A(n613), .ZN(n990) );
  XOR2_X1 U571 ( .A(KEYINPUT64), .B(n529), .Z(n651) );
  AND2_X1 U572 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U574 ( .A1(n654), .A2(G89), .ZN(n528) );
  XNOR2_X1 U575 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  INV_X1 U576 ( .A(G651), .ZN(n533) );
  OR2_X1 U577 ( .A1(n533), .A2(n635), .ZN(n529) );
  NAND2_X1 U578 ( .A1(G76), .A2(n651), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U580 ( .A(n532), .B(KEYINPUT5), .ZN(n541) );
  NOR2_X1 U581 ( .A1(G543), .A2(n533), .ZN(n535) );
  XNOR2_X1 U582 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n534) );
  XNOR2_X1 U583 ( .A(n535), .B(n534), .ZN(n649) );
  NAND2_X1 U584 ( .A1(n649), .A2(G63), .ZN(n536) );
  XNOR2_X1 U585 ( .A(n536), .B(KEYINPUT74), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G51), .A2(n650), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U588 ( .A(KEYINPUT6), .B(n539), .Z(n540) );
  NAND2_X1 U589 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U590 ( .A(n542), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U591 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n543) );
  XOR2_X2 U593 ( .A(KEYINPUT17), .B(n543), .Z(n875) );
  NAND2_X1 U594 ( .A1(G138), .A2(n875), .ZN(n545) );
  INV_X1 U595 ( .A(G2105), .ZN(n546) );
  AND2_X1 U596 ( .A1(n546), .A2(G2104), .ZN(n876) );
  NAND2_X1 U597 ( .A1(G102), .A2(n876), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n550) );
  NOR2_X1 U599 ( .A1(G2104), .A2(n546), .ZN(n879) );
  NAND2_X1 U600 ( .A1(G126), .A2(n879), .ZN(n548) );
  AND2_X1 U601 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U602 ( .A1(G114), .A2(n880), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U604 ( .A1(n550), .A2(n549), .ZN(G164) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U606 ( .A1(G99), .A2(n876), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G111), .A2(n880), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G123), .A2(n879), .ZN(n553) );
  XNOR2_X1 U610 ( .A(n553), .B(KEYINPUT18), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n554), .B(KEYINPUT75), .ZN(n555) );
  NOR2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n875), .A2(G135), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n926) );
  XNOR2_X1 U615 ( .A(G2096), .B(n926), .ZN(n559) );
  OR2_X1 U616 ( .A1(G2100), .A2(n559), .ZN(G156) );
  INV_X1 U617 ( .A(G57), .ZN(G237) );
  NAND2_X1 U618 ( .A1(G52), .A2(n650), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G64), .A2(n649), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n568) );
  XNOR2_X1 U621 ( .A(KEYINPUT9), .B(KEYINPUT68), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G77), .A2(n651), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n654), .A2(G90), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT67), .B(n562), .Z(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U626 ( .A(n566), .B(n565), .Z(n567) );
  NOR2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U628 ( .A(KEYINPUT69), .B(n569), .Z(G171) );
  NAND2_X1 U629 ( .A1(n879), .A2(G125), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G101), .A2(n876), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT23), .B(n570), .Z(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G137), .A2(n875), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G113), .A2(n880), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(G160) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U638 ( .A(n577), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U639 ( .A(G223), .B(KEYINPUT70), .Z(n821) );
  NAND2_X1 U640 ( .A1(n821), .A2(G567), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT11), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT71), .B(n579), .ZN(G234) );
  NAND2_X1 U643 ( .A1(G68), .A2(n651), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT72), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n654), .A2(G81), .ZN(n581) );
  XNOR2_X1 U646 ( .A(KEYINPUT12), .B(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n584), .B(KEYINPUT13), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G43), .A2(n650), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n649), .A2(G56), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n587), .Z(n588) );
  NOR2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n591) );
  INV_X1 U653 ( .A(KEYINPUT73), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n591), .B(n590), .ZN(n613) );
  NAND2_X1 U655 ( .A1(n613), .A2(G860), .ZN(G153) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U658 ( .A1(G54), .A2(n650), .ZN(n593) );
  NAND2_X1 U659 ( .A1(G66), .A2(n649), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U661 ( .A1(G92), .A2(n654), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G79), .A2(n651), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U665 ( .A(n598), .B(KEYINPUT15), .ZN(n978) );
  INV_X1 U666 ( .A(G868), .ZN(n614) );
  NAND2_X1 U667 ( .A1(n978), .A2(n614), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G53), .A2(n650), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G65), .A2(n649), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G91), .A2(n654), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G78), .A2(n651), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U675 ( .A1(n606), .A2(n605), .ZN(n973) );
  INV_X1 U676 ( .A(n973), .ZN(G299) );
  NOR2_X1 U677 ( .A1(G286), .A2(n614), .ZN(n608) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(G297) );
  INV_X1 U680 ( .A(G559), .ZN(n611) );
  NOR2_X1 U681 ( .A1(G860), .A2(n611), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n978), .A2(n609), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT16), .B(n610), .Z(G148) );
  INV_X1 U684 ( .A(n978), .ZN(n623) );
  NAND2_X1 U685 ( .A1(n611), .A2(n623), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n612), .A2(G868), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n990), .A2(n614), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G93), .A2(n654), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G80), .A2(n651), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G55), .A2(n650), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G67), .A2(n649), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n670) );
  XNOR2_X1 U696 ( .A(KEYINPUT76), .B(n990), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n623), .A2(G559), .ZN(n668) );
  XNOR2_X1 U698 ( .A(n624), .B(n668), .ZN(n625) );
  NOR2_X1 U699 ( .A1(G860), .A2(n625), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n670), .B(n626), .ZN(G145) );
  NAND2_X1 U701 ( .A1(G61), .A2(n649), .ZN(n633) );
  NAND2_X1 U702 ( .A1(G48), .A2(n650), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G86), .A2(n654), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n651), .A2(G73), .ZN(n629) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U713 ( .A1(n649), .A2(n638), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G49), .A2(n650), .ZN(n639) );
  XOR2_X1 U715 ( .A(KEYINPUT77), .B(n639), .Z(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G85), .A2(n654), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G60), .A2(n649), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G47), .A2(n650), .ZN(n644) );
  XOR2_X1 U721 ( .A(KEYINPUT66), .B(n644), .Z(n645) );
  NOR2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G72), .A2(n651), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(G290) );
  NAND2_X1 U725 ( .A1(G62), .A2(n649), .ZN(n659) );
  NAND2_X1 U726 ( .A1(G50), .A2(n650), .ZN(n653) );
  NAND2_X1 U727 ( .A1(G75), .A2(n651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U729 ( .A1(G88), .A2(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(KEYINPUT79), .B(n655), .ZN(n656) );
  NOR2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT80), .ZN(G303) );
  INV_X1 U734 ( .A(G303), .ZN(G166) );
  XOR2_X1 U735 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n661) );
  XNOR2_X1 U736 ( .A(G288), .B(n661), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n662), .B(G290), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n973), .B(n670), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(G166), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U741 ( .A(G305), .B(n666), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n667), .B(n990), .ZN(n850) );
  XNOR2_X1 U743 ( .A(n668), .B(n850), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n669), .A2(G868), .ZN(n672) );
  OR2_X1 U745 ( .A1(n670), .A2(G868), .ZN(n671) );
  NAND2_X1 U746 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U753 ( .A1(G132), .A2(G82), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n677), .B(KEYINPUT82), .ZN(n678) );
  XNOR2_X1 U755 ( .A(n678), .B(KEYINPUT22), .ZN(n679) );
  NOR2_X1 U756 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U757 ( .A1(G96), .A2(n680), .ZN(n825) );
  NAND2_X1 U758 ( .A1(n825), .A2(G2106), .ZN(n684) );
  NAND2_X1 U759 ( .A1(G120), .A2(G69), .ZN(n681) );
  NOR2_X1 U760 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U761 ( .A1(G108), .A2(n682), .ZN(n826) );
  NAND2_X1 U762 ( .A1(n826), .A2(G567), .ZN(n683) );
  NAND2_X1 U763 ( .A1(n684), .A2(n683), .ZN(n827) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U765 ( .A1(n827), .A2(n685), .ZN(n824) );
  NAND2_X1 U766 ( .A1(n824), .A2(G36), .ZN(G176) );
  AND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n771) );
  NAND2_X1 U768 ( .A1(G8), .A2(n733), .ZN(n780) );
  NOR2_X1 U769 ( .A1(G1976), .A2(G288), .ZN(n688) );
  NAND2_X1 U770 ( .A1(n688), .A2(KEYINPUT33), .ZN(n686) );
  NOR2_X1 U771 ( .A1(n780), .A2(n686), .ZN(n753) );
  NOR2_X1 U772 ( .A1(G303), .A2(G1971), .ZN(n687) );
  NOR2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n982) );
  INV_X1 U774 ( .A(n733), .ZN(n714) );
  NAND2_X1 U775 ( .A1(n714), .A2(G2072), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n689), .B(KEYINPUT27), .ZN(n691) );
  INV_X1 U777 ( .A(G1956), .ZN(n1004) );
  NOR2_X1 U778 ( .A1(n1004), .A2(n714), .ZN(n690) );
  NOR2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n705) );
  NOR2_X1 U780 ( .A1(n973), .A2(n705), .ZN(n693) );
  XNOR2_X1 U781 ( .A(KEYINPUT89), .B(KEYINPUT28), .ZN(n692) );
  XNOR2_X1 U782 ( .A(n693), .B(n692), .ZN(n709) );
  INV_X1 U783 ( .A(G1996), .ZN(n792) );
  NOR2_X1 U784 ( .A1(n733), .A2(n792), .ZN(n694) );
  XOR2_X1 U785 ( .A(n694), .B(KEYINPUT26), .Z(n696) );
  NAND2_X1 U786 ( .A1(n733), .A2(G1341), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U788 ( .A1(n990), .A2(n697), .ZN(n701) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n733), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n714), .A2(G2067), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U792 ( .A1(n978), .A2(n702), .ZN(n700) );
  OR2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n978), .A2(n702), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n973), .A2(n705), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U799 ( .A1(n714), .A2(G1961), .ZN(n712) );
  XNOR2_X1 U800 ( .A(n712), .B(KEYINPUT87), .ZN(n716) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n713), .B(KEYINPUT88), .ZN(n956) );
  NAND2_X1 U803 ( .A1(n956), .A2(n714), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n725) );
  NAND2_X1 U805 ( .A1(n725), .A2(G171), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n732) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n780), .ZN(n745) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n733), .ZN(n741) );
  INV_X1 U809 ( .A(n741), .ZN(n719) );
  NAND2_X1 U810 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U811 ( .A(n721), .B(KEYINPUT30), .ZN(n722) );
  XNOR2_X1 U812 ( .A(n722), .B(KEYINPUT90), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n723), .A2(G168), .ZN(n724) );
  XOR2_X1 U814 ( .A(KEYINPUT91), .B(n724), .Z(n728) );
  NOR2_X1 U815 ( .A1(G171), .A2(n725), .ZN(n726) );
  XNOR2_X1 U816 ( .A(KEYINPUT92), .B(n726), .ZN(n727) );
  NOR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U818 ( .A1(n732), .A2(n731), .ZN(n743) );
  NAND2_X1 U819 ( .A1(n743), .A2(G286), .ZN(n738) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n780), .ZN(n735) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U825 ( .A1(G8), .A2(n739), .ZN(n740) );
  NAND2_X1 U826 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n743), .A2(n742), .ZN(n744) );
  INV_X1 U828 ( .A(n783), .ZN(n747) );
  NAND2_X1 U829 ( .A1(n982), .A2(n747), .ZN(n750) );
  NAND2_X1 U830 ( .A1(G288), .A2(G1976), .ZN(n748) );
  XNOR2_X1 U831 ( .A(n748), .B(KEYINPUT94), .ZN(n974) );
  INV_X1 U832 ( .A(n974), .ZN(n749) );
  AND2_X1 U833 ( .A1(n750), .A2(n526), .ZN(n751) );
  NOR2_X1 U834 ( .A1(KEYINPUT33), .A2(n751), .ZN(n752) );
  NOR2_X1 U835 ( .A1(n753), .A2(n752), .ZN(n776) );
  XOR2_X1 U836 ( .A(G1981), .B(G305), .Z(n985) );
  NAND2_X1 U837 ( .A1(G95), .A2(n876), .ZN(n755) );
  NAND2_X1 U838 ( .A1(G107), .A2(n880), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n761) );
  NAND2_X1 U840 ( .A1(G131), .A2(n875), .ZN(n756) );
  XNOR2_X1 U841 ( .A(n756), .B(KEYINPUT86), .ZN(n759) );
  NAND2_X1 U842 ( .A1(G119), .A2(n879), .ZN(n757) );
  XOR2_X1 U843 ( .A(KEYINPUT85), .B(n757), .Z(n758) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U845 ( .A1(n761), .A2(n760), .ZN(n893) );
  INV_X1 U846 ( .A(G1991), .ZN(n949) );
  NOR2_X1 U847 ( .A1(n893), .A2(n949), .ZN(n770) );
  NAND2_X1 U848 ( .A1(n876), .A2(G105), .ZN(n762) );
  XNOR2_X1 U849 ( .A(n762), .B(KEYINPUT38), .ZN(n764) );
  NAND2_X1 U850 ( .A1(G129), .A2(n879), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U852 ( .A1(G141), .A2(n875), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G117), .A2(n880), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n886) );
  NOR2_X1 U856 ( .A1(n886), .A2(n792), .ZN(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n796) );
  XOR2_X1 U858 ( .A(G1986), .B(G290), .Z(n977) );
  NAND2_X1 U859 ( .A1(n796), .A2(n977), .ZN(n774) );
  INV_X1 U860 ( .A(n771), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n817) );
  NAND2_X1 U862 ( .A1(n774), .A2(n817), .ZN(n777) );
  AND2_X1 U863 ( .A1(n985), .A2(n777), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n791) );
  INV_X1 U865 ( .A(n777), .ZN(n789) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U867 ( .A(n778), .B(KEYINPUT24), .Z(n779) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n787) );
  INV_X1 U869 ( .A(n780), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G166), .A2(G8), .ZN(n781) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n781), .ZN(n782) );
  NOR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  AND2_X1 U876 ( .A1(n791), .A2(n790), .ZN(n815) );
  AND2_X1 U877 ( .A1(n792), .A2(n886), .ZN(n936) );
  AND2_X1 U878 ( .A1(n893), .A2(n949), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n793), .B(KEYINPUT96), .ZN(n929) );
  NOR2_X1 U880 ( .A1(G1986), .A2(G290), .ZN(n794) );
  XOR2_X1 U881 ( .A(n794), .B(KEYINPUT95), .Z(n795) );
  NOR2_X1 U882 ( .A1(n929), .A2(n795), .ZN(n797) );
  INV_X1 U883 ( .A(n796), .ZN(n923) );
  NOR2_X1 U884 ( .A1(n797), .A2(n923), .ZN(n798) );
  NOR2_X1 U885 ( .A1(n936), .A2(n798), .ZN(n799) );
  XNOR2_X1 U886 ( .A(KEYINPUT39), .B(n799), .ZN(n800) );
  NAND2_X1 U887 ( .A1(n800), .A2(n817), .ZN(n813) );
  XOR2_X1 U888 ( .A(G2067), .B(KEYINPUT37), .Z(n816) );
  NAND2_X1 U889 ( .A1(G140), .A2(n875), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G104), .A2(n876), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(KEYINPUT34), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n804), .B(KEYINPUT83), .ZN(n810) );
  XNOR2_X1 U894 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G128), .A2(n879), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G116), .A2(n880), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U898 ( .A(n808), .B(n807), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(KEYINPUT36), .B(n811), .ZN(n896) );
  NOR2_X1 U901 ( .A1(n816), .A2(n896), .ZN(n932) );
  NAND2_X1 U902 ( .A1(n932), .A2(n817), .ZN(n812) );
  AND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n819) );
  AND2_X1 U905 ( .A1(n816), .A2(n896), .ZN(n924) );
  NAND2_X1 U906 ( .A1(n924), .A2(n817), .ZN(n818) );
  XNOR2_X1 U907 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U910 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U912 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U913 ( .A(G69), .B(KEYINPUT100), .Z(G235) );
  INV_X1 U915 ( .A(G132), .ZN(G219) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G82), .ZN(G220) );
  NOR2_X1 U918 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  INV_X1 U920 ( .A(n827), .ZN(G319) );
  XOR2_X1 U921 ( .A(KEYINPUT101), .B(G2090), .Z(n829) );
  XNOR2_X1 U922 ( .A(G2067), .B(G2084), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U924 ( .A(n830), .B(G2100), .Z(n832) );
  XNOR2_X1 U925 ( .A(G2078), .B(G2072), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U927 ( .A(G2096), .B(G2678), .Z(n834) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U930 ( .A(n836), .B(n835), .Z(G227) );
  XOR2_X1 U931 ( .A(KEYINPUT41), .B(KEYINPUT103), .Z(n838) );
  XNOR2_X1 U932 ( .A(KEYINPUT105), .B(G2474), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U934 ( .A(n839), .B(KEYINPUT104), .Z(n841) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n849) );
  XOR2_X1 U937 ( .A(G1981), .B(G1971), .Z(n843) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1956), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U940 ( .A(KEYINPUT102), .B(G1976), .Z(n845) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1961), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n847), .B(n846), .Z(n848) );
  XNOR2_X1 U944 ( .A(n849), .B(n848), .ZN(G229) );
  XNOR2_X1 U945 ( .A(G286), .B(n978), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n852), .B(G171), .ZN(n853) );
  NOR2_X1 U948 ( .A1(G37), .A2(n853), .ZN(G397) );
  NAND2_X1 U949 ( .A1(G124), .A2(n879), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n854), .B(KEYINPUT106), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G136), .A2(n875), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U954 ( .A1(G100), .A2(n876), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G112), .A2(n880), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U957 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U958 ( .A(KEYINPUT107), .B(n862), .Z(G162) );
  NAND2_X1 U959 ( .A1(n876), .A2(G106), .ZN(n863) );
  XOR2_X1 U960 ( .A(KEYINPUT109), .B(n863), .Z(n865) );
  NAND2_X1 U961 ( .A1(n875), .A2(G142), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n866), .B(KEYINPUT45), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G130), .A2(n879), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U966 ( .A1(n880), .A2(G118), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT108), .B(n869), .Z(n870) );
  NOR2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n874) );
  XOR2_X1 U969 ( .A(G160), .B(G162), .Z(n872) );
  XNOR2_X1 U970 ( .A(n926), .B(n872), .ZN(n873) );
  XOR2_X1 U971 ( .A(n874), .B(n873), .Z(n888) );
  NAND2_X1 U972 ( .A1(G139), .A2(n875), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G103), .A2(n876), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U975 ( .A1(G127), .A2(n879), .ZN(n882) );
  NAND2_X1 U976 ( .A1(G115), .A2(n880), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U979 ( .A1(n885), .A2(n884), .ZN(n919) );
  XNOR2_X1 U980 ( .A(n886), .B(n919), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U982 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n890) );
  XNOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U985 ( .A(n892), .B(n891), .Z(n895) );
  XNOR2_X1 U986 ( .A(G164), .B(n893), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U988 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U989 ( .A1(G37), .A2(n898), .ZN(n899) );
  XNOR2_X1 U990 ( .A(KEYINPUT112), .B(n899), .ZN(G395) );
  XOR2_X1 U991 ( .A(KEYINPUT97), .B(G2446), .Z(n901) );
  XNOR2_X1 U992 ( .A(G2430), .B(G2451), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U994 ( .A(n902), .B(KEYINPUT98), .Z(n904) );
  XNOR2_X1 U995 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U997 ( .A(KEYINPUT99), .B(G2438), .Z(n906) );
  XNOR2_X1 U998 ( .A(G2435), .B(G2454), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1000 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1001 ( .A(G2443), .B(G2427), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(n911), .A2(G14), .ZN(n918) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n912) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n912), .Z(n913) );
  XNOR2_X1 U1007 ( .A(n913), .B(KEYINPUT113), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1009 ( .A1(G397), .A2(G395), .ZN(n916) );
  NAND2_X1 U1010 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1018 ( .A(KEYINPUT50), .B(n922), .Z(n942) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n934) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(KEYINPUT114), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1024 ( .A(KEYINPUT115), .B(n930), .ZN(n931) );
  NOR2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1026 ( .A1(n934), .A2(n933), .ZN(n939) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(n937), .B(KEYINPUT51), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1031 ( .A(KEYINPUT116), .B(n940), .Z(n941) );
  NOR2_X1 U1032 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n943), .ZN(n944) );
  XNOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n967) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n967), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n945), .A2(G29), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT118), .B(n946), .ZN(n1030) );
  XNOR2_X1 U1038 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(n947), .B(G34), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G2084), .B(n948), .ZN(n966) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G35), .ZN(n964) );
  XNOR2_X1 U1042 ( .A(n949), .B(G25), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n951), .B(KEYINPUT119), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n961) );
  XOR2_X1 U1049 ( .A(n956), .B(G27), .Z(n958) );
  XNOR2_X1 U1050 ( .A(G32), .B(G1996), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT120), .B(n959), .Z(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(KEYINPUT122), .B(n967), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(n969), .B(n968), .ZN(n971) );
  INV_X1 U1059 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1061 ( .A1(n972), .A2(G11), .ZN(n1028) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XNOR2_X1 U1063 ( .A(n973), .B(G1956), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n984) );
  NAND2_X1 U1065 ( .A1(G303), .A2(G1971), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n978), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n994) );
  XNOR2_X1 U1071 ( .A(G171), .B(G1961), .ZN(n989) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(n987), .B(KEYINPUT57), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1076 ( .A(G1341), .B(n990), .ZN(n991) );
  NOR2_X1 U1077 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1078 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1079 ( .A1(n996), .A2(n995), .ZN(n1026) );
  INV_X1 U1080 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1081 ( .A(G1986), .B(G24), .ZN(n1001) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G22), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(G1976), .B(G23), .ZN(n997) );
  NOR2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(KEYINPUT127), .B(n999), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(KEYINPUT58), .B(n1002), .ZN(n1018) );
  XOR2_X1 U1088 ( .A(G1981), .B(G6), .Z(n1003) );
  XNOR2_X1 U1089 ( .A(KEYINPUT123), .B(n1003), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(G1341), .B(G19), .Z(n1006) );
  XNOR2_X1 U1091 ( .A(n1004), .B(G20), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(KEYINPUT124), .B(n1009), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(G1348), .B(KEYINPUT59), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1010), .B(G4), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1013), .B(KEYINPUT125), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1014), .Z(n1016) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G5), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XNOR2_X1 U1103 ( .A(KEYINPUT126), .B(G1966), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(G21), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1109 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1110 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

