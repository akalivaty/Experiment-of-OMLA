//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT78), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n187), .A2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n196), .B(KEYINPUT3), .C1(new_n187), .C2(G107), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G101), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n194), .B1(new_n191), .B2(new_n190), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n189), .A4(new_n197), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n204));
  INV_X1    g018(.A(G113), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT68), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(KEYINPUT2), .B2(G113), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n206), .A2(new_n208), .B1(KEYINPUT2), .B2(G113), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G116), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G119), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n209), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n198), .A2(new_n216), .A3(G101), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n203), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n190), .B2(new_n194), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n202), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(KEYINPUT5), .ZN(new_n221));
  OAI21_X1  g035(.A(G113), .B1(new_n211), .B2(KEYINPUT5), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n221), .A2(new_n223), .B1(new_n209), .B2(new_n214), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n218), .A2(new_n225), .A3(new_n227), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(KEYINPUT6), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT6), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n232), .A3(new_n228), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G128), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT64), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G143), .ZN(new_n238));
  INV_X1    g052(.A(G143), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n241), .A2(new_n242), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n234), .A2(KEYINPUT0), .A3(G128), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G125), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n239), .B(G146), .C1(new_n249), .C2(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n237), .A3(G143), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n234), .A2(new_n253), .A3(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n248), .B1(G125), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G224), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n258), .B(KEYINPUT81), .Z(new_n259));
  XNOR2_X1  g073(.A(new_n256), .B(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n231), .A2(new_n233), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n258), .A2(KEYINPUT7), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n256), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n209), .A2(new_n214), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n221), .B1(KEYINPUT82), .B2(new_n222), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n222), .A2(KEYINPUT82), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n220), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n227), .B(KEYINPUT8), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n202), .A2(new_n219), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n224), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n269), .A2(new_n272), .A3(KEYINPUT83), .A4(new_n270), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n264), .A2(new_n275), .A3(new_n230), .A4(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n261), .A2(new_n262), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(G210), .B1(G237), .B2(G902), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT84), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n261), .A2(new_n262), .A3(new_n279), .A4(new_n277), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n283), .A2(new_n282), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G214), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT9), .B(G234), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n247), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n203), .A2(new_n294), .A3(new_n217), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n250), .A2(new_n251), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n254), .B1(KEYINPUT79), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(KEYINPUT79), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n202), .B(new_n219), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n255), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n295), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G137), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(G137), .ZN(new_n307));
  INV_X1    g121(.A(G137), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT11), .A3(G134), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G131), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(KEYINPUT66), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n312), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n303), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(G110), .B(G140), .Z(new_n317));
  INV_X1    g131(.A(G227), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G953), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n313), .A2(new_n314), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n295), .A2(new_n301), .A3(new_n302), .A4(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(KEYINPUT80), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(KEYINPUT80), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n316), .B(new_n320), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n255), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n271), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n321), .B1(new_n327), .B2(new_n299), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n322), .A2(KEYINPUT80), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n322), .A2(KEYINPUT80), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(new_n320), .B(KEYINPUT77), .Z(new_n334));
  OAI211_X1 g148(.A(new_n325), .B(G469), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G469), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n262), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n331), .A2(new_n332), .B1(new_n315), .B2(new_n303), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n340), .A2(new_n320), .B1(new_n341), .B2(new_n330), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n336), .A3(new_n262), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n293), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n289), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n215), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n306), .A2(new_n309), .A3(new_n311), .A4(new_n307), .ZN(new_n347));
  INV_X1    g161(.A(new_n307), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n305), .A2(G137), .ZN(new_n349));
  OAI21_X1  g163(.A(G131), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n255), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n346), .B(new_n351), .C1(new_n321), .C2(new_n247), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT28), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n321), .B2(new_n247), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n215), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(G101), .ZN(new_n358));
  NOR2_X1   g172(.A1(G237), .A2(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G210), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT29), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n262), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n366));
  INV_X1    g180(.A(new_n351), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT65), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n247), .A2(new_n368), .B1(new_n313), .B2(new_n314), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n236), .A2(new_n245), .A3(KEYINPUT65), .A4(new_n246), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n366), .B1(new_n371), .B2(KEYINPUT30), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n247), .A2(new_n368), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n315), .A3(new_n370), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n351), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(KEYINPUT67), .A3(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n354), .A2(new_n376), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n372), .A2(new_n377), .A3(new_n215), .A4(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n361), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n352), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n352), .B(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n371), .A2(new_n346), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n361), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G472), .B1(new_n365), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n352), .A2(new_n361), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n379), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT31), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT69), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT31), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n379), .A2(new_n392), .A3(new_n388), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n379), .B2(new_n388), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT69), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT32), .ZN(new_n400));
  NOR2_X1   g214(.A1(G472), .A2(G902), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n387), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(G125), .A2(G140), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(G125), .A2(G140), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT16), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G125), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n409), .A2(KEYINPUT16), .A3(G140), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n411), .A3(G146), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n406), .A2(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n249), .A2(G119), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT73), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n416), .A2(KEYINPUT23), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(KEYINPUT23), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n417), .B(new_n418), .C1(G119), .C2(new_n249), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G110), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n414), .B(KEYINPUT72), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(G119), .B2(new_n249), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT24), .B(G110), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI221_X1 g238(.A(new_n412), .B1(G146), .B2(new_n413), .C1(new_n420), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(G110), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT16), .ZN(new_n427));
  INV_X1    g241(.A(G140), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n409), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n429), .B2(new_n405), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n237), .B1(new_n430), .B2(new_n410), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n412), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n426), .B(new_n432), .C1(new_n422), .C2(new_n423), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT22), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(G137), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n425), .B2(new_n433), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n439), .A3(G902), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT71), .B(G217), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(G234), .B2(new_n262), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT76), .ZN(new_n446));
  INV_X1    g260(.A(new_n439), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT25), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(KEYINPUT74), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n447), .A2(new_n262), .A3(new_n437), .A4(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n450), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n443), .B(new_n452), .C1(new_n440), .C2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT76), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n440), .A2(new_n455), .A3(new_n444), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n446), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n359), .A2(G143), .A3(G214), .ZN(new_n458));
  AOI21_X1  g272(.A(G143), .B1(new_n359), .B2(G214), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT17), .B(G131), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n431), .A3(new_n412), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G131), .B1(new_n458), .B2(new_n459), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT17), .ZN(new_n465));
  INV_X1    g279(.A(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n257), .A3(G214), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n239), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n359), .A2(G143), .A3(G214), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n311), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n460), .A2(new_n431), .A3(KEYINPUT86), .A4(new_n412), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n413), .B(G146), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT18), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n468), .B(new_n469), .C1(new_n475), .C2(new_n311), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n474), .B(new_n476), .C1(new_n475), .C2(new_n464), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G113), .B(G122), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(G104), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n458), .A2(new_n459), .A3(G131), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n311), .B1(new_n468), .B2(new_n469), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT85), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n413), .A2(KEYINPUT19), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n413), .A2(KEYINPUT19), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n237), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n464), .A2(new_n490), .A3(new_n470), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n486), .A2(new_n412), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n477), .A3(new_n480), .ZN(new_n493));
  NOR2_X1   g307(.A1(G475), .A2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n495), .A2(KEYINPUT88), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n482), .A2(new_n483), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(KEYINPUT88), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT89), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n480), .B1(new_n473), .B2(new_n477), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n492), .A2(new_n480), .A3(new_n477), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n501), .A2(new_n502), .A3(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT87), .B1(new_n503), .B2(new_n483), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT20), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n498), .A4(new_n496), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n482), .A2(new_n494), .A3(new_n493), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT87), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT20), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n500), .A2(new_n504), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G122), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G116), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT91), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n193), .B1(new_n514), .B2(KEYINPUT14), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(G116), .B2(new_n512), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G128), .B(G143), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n305), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n516), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(KEYINPUT13), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n249), .A2(KEYINPUT13), .A3(G143), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(new_n305), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n522), .A2(new_n524), .B1(new_n305), .B2(new_n518), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n516), .A2(G107), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n516), .A2(G107), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n291), .A2(G953), .A3(new_n442), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n521), .A2(new_n528), .A3(new_n530), .ZN(new_n533));
  AOI21_X1  g347(.A(G902), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n534), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(G234), .A2(G237), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(G952), .A3(new_n257), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT21), .B(G898), .Z(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(G902), .A3(G953), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n480), .A2(KEYINPUT90), .ZN(new_n543));
  AOI21_X1  g357(.A(G902), .B1(new_n478), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n543), .B2(new_n478), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G475), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n511), .A2(new_n537), .A3(new_n542), .A4(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(KEYINPUT92), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(KEYINPUT92), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n345), .A2(new_n404), .A3(new_n457), .A4(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(G101), .ZN(G3));
  NAND2_X1  g366(.A1(new_n399), .A2(new_n401), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n396), .A2(new_n397), .ZN(new_n554));
  AOI211_X1 g368(.A(KEYINPUT69), .B(new_n392), .C1(new_n379), .C2(new_n388), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n393), .A2(new_n394), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G472), .B1(new_n557), .B2(G902), .ZN(new_n558));
  AND4_X1   g372(.A1(new_n553), .A2(new_n344), .A3(new_n558), .A4(new_n457), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n532), .A2(new_n533), .ZN(new_n560));
  AND2_X1   g374(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n561));
  NOR2_X1   g375(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n561), .B1(new_n532), .B2(new_n533), .ZN(new_n565));
  OAI21_X1  g379(.A(G478), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n534), .A2(new_n535), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n535), .A2(new_n262), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n500), .A2(new_n507), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n504), .A2(new_n510), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n546), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n288), .B1(new_n281), .B2(new_n283), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n542), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n559), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT34), .B(G104), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(G6));
  INV_X1    g395(.A(new_n536), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n534), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n505), .A2(new_n494), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n504), .A2(new_n510), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n546), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n559), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G107), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G9));
  NAND2_X1  g404(.A1(new_n558), .A2(new_n553), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n425), .A2(new_n433), .ZN(new_n593));
  INV_X1    g407(.A(new_n436), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(KEYINPUT36), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(KEYINPUT36), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n425), .A2(new_n433), .A3(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n595), .A2(new_n262), .A3(new_n444), .A4(new_n597), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n454), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n345), .A2(new_n550), .A3(new_n592), .A4(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT37), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G110), .ZN(G12));
  NAND2_X1  g418(.A1(new_n339), .A2(new_n343), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n605), .A2(new_n292), .A3(new_n576), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n539), .B(KEYINPUT96), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT95), .B(G900), .Z(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n541), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n583), .A2(new_n585), .A3(new_n546), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT97), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n404), .A2(new_n606), .A3(new_n601), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G128), .ZN(G30));
  AOI21_X1  g429(.A(new_n380), .B1(new_n379), .B2(new_n352), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n355), .A2(new_n352), .A3(new_n380), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n262), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n402), .B2(new_n403), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n284), .A2(new_n621), .A3(new_n285), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n284), .B2(new_n285), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n599), .A2(new_n454), .A3(new_n600), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n583), .A3(new_n574), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n620), .A2(new_n624), .A3(new_n627), .A4(new_n287), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n401), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT32), .B1(new_n557), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n626), .B1(new_n634), .B2(new_n619), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(KEYINPUT98), .A3(new_n287), .A4(new_n624), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n610), .B(KEYINPUT39), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n344), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n630), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G143), .ZN(G45));
  NOR2_X1   g457(.A1(new_n575), .A2(new_n610), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n404), .A2(new_n606), .A3(new_n601), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G146), .ZN(G48));
  NAND2_X1  g460(.A1(new_n342), .A2(new_n262), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(G469), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n343), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n293), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n404), .A2(new_n578), .A3(new_n457), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT41), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G113), .ZN(G15));
  NAND4_X1  g467(.A1(new_n404), .A2(new_n457), .A3(new_n587), .A4(new_n650), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G116), .ZN(G18));
  AOI21_X1  g469(.A(new_n625), .B1(new_n634), .B2(new_n387), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n648), .A2(new_n576), .A3(new_n292), .A4(new_n343), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n548), .B2(new_n549), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n656), .A2(KEYINPUT99), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  INV_X1    g478(.A(new_n574), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n537), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n666), .A2(new_n542), .A3(new_n576), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n356), .A2(new_n380), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n393), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n401), .B1(new_n669), .B2(new_n396), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(KEYINPUT100), .B(new_n401), .C1(new_n669), .C2(new_n396), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n399), .B2(new_n262), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n667), .A2(new_n457), .A3(new_n650), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT101), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G122), .ZN(G24));
  NOR3_X1   g494(.A1(new_n674), .A2(new_n676), .A3(new_n625), .ZN(new_n681));
  INV_X1    g495(.A(new_n657), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n644), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  AND2_X1   g498(.A1(new_n404), .A2(new_n457), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n288), .B1(new_n284), .B2(new_n285), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n344), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n644), .A4(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n404), .A2(new_n687), .A3(new_n457), .A4(new_n644), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n387), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n687), .A2(new_n644), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n457), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G131), .ZN(G33));
  NAND4_X1  g514(.A1(new_n404), .A2(new_n687), .A3(new_n457), .A4(new_n613), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT104), .B(G134), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G36));
  INV_X1    g517(.A(new_n343), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n325), .B1(new_n333), .B2(new_n334), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n325), .B(KEYINPUT45), .C1(new_n333), .C2(new_n334), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(G469), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n338), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n704), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n709), .A2(KEYINPUT46), .A3(new_n338), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n293), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n638), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n574), .A2(new_n570), .A3(KEYINPUT43), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n574), .A2(KEYINPUT105), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n511), .A2(new_n719), .A3(new_n546), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n570), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n554), .A2(new_n555), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n631), .B1(new_n724), .B2(new_n395), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n601), .B1(new_n676), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT106), .B(new_n601), .C1(new_n676), .C2(new_n725), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n715), .B1(KEYINPUT44), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n718), .A2(new_n720), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n571), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n716), .B1(new_n733), .B2(KEYINPUT43), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT106), .B1(new_n591), .B2(new_n601), .ZN(new_n735));
  INV_X1    g549(.A(new_n729), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT107), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n730), .A2(new_n740), .A3(KEYINPUT44), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n686), .B(new_n731), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G137), .ZN(G39));
  NAND2_X1  g557(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n714), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n714), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n686), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n404), .A2(new_n457), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n745), .A2(new_n747), .A3(new_n644), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  OAI21_X1  g565(.A(new_n721), .B1(KEYINPUT49), .B2(new_n649), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(KEYINPUT49), .B2(new_n649), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n457), .A2(new_n287), .A3(new_n292), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n756), .A2(new_n624), .A3(new_n620), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n734), .A2(new_n607), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n677), .A2(new_n457), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n748), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n745), .A2(new_n747), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n649), .A2(new_n292), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n650), .A2(new_n686), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n681), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n620), .ZN(new_n770));
  INV_X1    g584(.A(new_n539), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n457), .A3(new_n771), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n772), .A2(new_n574), .A3(new_n571), .ZN(new_n773));
  INV_X1    g587(.A(new_n650), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n758), .A2(new_n774), .A3(new_n759), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n624), .A2(new_n287), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n775), .A2(KEYINPUT50), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT50), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n769), .B(new_n773), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT51), .B1(new_n766), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n761), .B1(new_n762), .B2(new_n765), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n783));
  OAI211_X1 g597(.A(G952), .B(new_n257), .C1(new_n783), .C2(new_n779), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n697), .A2(new_n681), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n537), .A2(new_n585), .A3(new_n546), .A4(new_n611), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n656), .A2(new_n687), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(new_n791), .A3(new_n701), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n693), .B2(new_n698), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n559), .A2(new_n542), .A3(new_n289), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n665), .A2(new_n583), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n602), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n575), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n559), .A2(new_n542), .A3(new_n289), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n551), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT111), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n551), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n796), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n678), .A2(new_n651), .A3(new_n654), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n663), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n804), .B1(new_n663), .B2(new_n805), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n793), .B(new_n803), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n620), .A2(new_n606), .A3(new_n627), .A4(new_n611), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n614), .A2(new_n645), .A3(new_n811), .A4(new_n683), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT52), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n812), .B(KEYINPUT52), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n816), .B(KEYINPUT54), .C1(new_n810), .C2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n772), .A2(new_n575), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n810), .B1(new_n808), .B2(new_n817), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n663), .A2(new_n805), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n699), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT114), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n792), .A2(new_n810), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n803), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n822), .A2(new_n699), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n826), .A3(new_n815), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n785), .A2(new_n819), .A3(new_n820), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n760), .A2(new_n657), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n696), .A2(new_n457), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n768), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT48), .Z(new_n836));
  NOR3_X1   g650(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(G952), .A2(G953), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT116), .Z(new_n839));
  OAI21_X1  g653(.A(new_n757), .B1(new_n837), .B2(new_n839), .ZN(G75));
  NOR2_X1   g654(.A1(new_n257), .A2(G952), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n821), .A2(new_n829), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(G902), .ZN(new_n843));
  INV_X1    g657(.A(G210), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n231), .A2(new_n233), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(new_n260), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT55), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n843), .A2(new_n844), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n262), .B1(new_n821), .B2(new_n829), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT118), .B1(new_n851), .B2(G210), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n849), .B(new_n850), .C1(new_n845), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n848), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n841), .B1(new_n853), .B2(new_n855), .ZN(G51));
  NAND2_X1  g670(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n831), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n842), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n337), .B(KEYINPUT57), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n342), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n843), .A2(new_n709), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n841), .B1(new_n863), .B2(new_n864), .ZN(G54));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(KEYINPUT58), .B2(G475), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n843), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n501), .A2(new_n502), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n841), .ZN(G60));
  INV_X1    g687(.A(new_n841), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n568), .B(KEYINPUT59), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n819), .B2(new_n831), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n564), .A2(new_n565), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n859), .A2(new_n860), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n564), .A2(new_n565), .A3(new_n875), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(G63));
  NAND2_X1  g695(.A1(G217), .A2(G902), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT60), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n821), .B2(new_n829), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n597), .A3(new_n595), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n438), .A2(new_n439), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n885), .B(new_n874), .C1(new_n886), .C2(new_n884), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(G66));
  NAND2_X1  g703(.A1(new_n540), .A2(G224), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT121), .ZN(new_n893));
  OAI211_X1 g707(.A(KEYINPUT122), .B(new_n891), .C1(new_n893), .C2(G953), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n893), .A2(G953), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(KEYINPUT122), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n846), .B1(G898), .B2(new_n257), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n896), .B(new_n897), .Z(G69));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n614), .A2(new_n645), .A3(new_n683), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n614), .A2(new_n645), .A3(new_n683), .A4(KEYINPUT124), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n642), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n903), .A2(new_n642), .A3(KEYINPUT62), .A4(new_n904), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n639), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n795), .A2(new_n575), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n685), .A2(new_n910), .A3(new_n686), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n742), .A2(new_n750), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n900), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n742), .A2(new_n750), .A3(new_n912), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n907), .A2(new_n908), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(KEYINPUT125), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(G953), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n372), .A2(new_n377), .A3(new_n378), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n487), .A2(new_n488), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n899), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n909), .A2(new_n900), .A3(new_n913), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT125), .B1(new_n915), .B2(new_n916), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n257), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n922), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(KEYINPUT126), .A3(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n666), .A2(new_n576), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n834), .A2(new_n638), .A3(new_n929), .A4(new_n714), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n742), .A2(new_n701), .A3(new_n750), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n699), .A2(new_n903), .A3(new_n904), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n257), .ZN(new_n934));
  INV_X1    g748(.A(G900), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n934), .B(new_n922), .C1(new_n935), .C2(new_n257), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n923), .A2(new_n928), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n318), .B2(new_n935), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT127), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n923), .A2(new_n928), .A3(new_n939), .A4(new_n936), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(G72));
  NAND2_X1  g757(.A1(G472), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT63), .Z(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n893), .B2(new_n933), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n874), .B1(new_n947), .B2(new_n381), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n816), .B1(new_n810), .B2(new_n818), .ZN(new_n949));
  INV_X1    g763(.A(new_n381), .ZN(new_n950));
  NOR4_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n616), .A4(new_n946), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n893), .A2(new_n914), .A3(new_n917), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n945), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n948), .B(new_n951), .C1(new_n616), .C2(new_n953), .ZN(G57));
endmodule


