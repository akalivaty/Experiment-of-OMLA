//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n459), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  OAI21_X1  g044(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G112), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G2105), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT65), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n460), .A2(new_n461), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n459), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n475), .A2(G136), .B1(G124), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n473), .A2(new_n479), .ZN(G162));
  OAI211_X1 g055(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(new_n459), .A3(G138), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n474), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n476), .A2(new_n477), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n484), .A2(new_n459), .A3(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(KEYINPUT67), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n482), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n459), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT66), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n459), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(new_n492), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n494), .A2(new_n497), .B1(new_n478), .B2(G126), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n490), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n510), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n508), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n509), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(new_n516), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n521), .B(new_n523), .C1(new_n527), .C2(KEYINPUT69), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n527), .A2(KEYINPUT69), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n507), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n510), .A2(new_n533), .B1(new_n516), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  INV_X1    g111(.A(new_n516), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT70), .B(G81), .Z(new_n538));
  AOI22_X1  g113(.A1(G43), .A2(new_n522), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n507), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n549));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n510), .B2(new_n550), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n522), .A2(KEYINPUT71), .A3(G53), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .A3(new_n551), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n516), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n505), .A2(new_n509), .A3(KEYINPUT72), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(G91), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n507), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n552), .A2(new_n554), .A3(new_n558), .A4(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  NAND3_X1  g138(.A1(new_n556), .A2(G87), .A3(new_n557), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n522), .A2(G49), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  OAI211_X1 g142(.A(G48), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(G61), .B1(new_n513), .B2(new_n512), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n507), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n569), .B1(new_n572), .B2(KEYINPUT73), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n507), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n556), .A2(G86), .A3(new_n557), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n507), .ZN(new_n580));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n510), .A2(new_n581), .B1(new_n516), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n556), .A2(G92), .A3(new_n557), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT10), .Z(new_n589));
  NAND2_X1  g164(.A1(new_n505), .A2(G66), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n507), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(G54), .B2(new_n522), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G321));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G299), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G168), .B2(new_n598), .ZN(G280));
  XOR2_X1   g175(.A(G280), .B(KEYINPUT75), .Z(G297));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n542), .A2(new_n598), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n594), .A2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n598), .ZN(G323));
  XOR2_X1   g181(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n607));
  XNOR2_X1  g182(.A(G323), .B(new_n607), .ZN(G282));
  NAND2_X1  g183(.A1(new_n487), .A2(new_n466), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n475), .A2(G135), .B1(G123), .B2(new_n478), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n616));
  NOR3_X1   g191(.A1(new_n616), .A2(new_n459), .A3(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n459), .B2(G111), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n615), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND3_X1  g196(.A1(new_n613), .A2(new_n614), .A3(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT78), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT17), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT80), .Z(new_n647));
  INV_X1    g222(.A(new_n643), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n645), .A2(new_n641), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n643), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n644), .B1(new_n648), .B2(new_n641), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2096), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT81), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n663), .B1(new_n661), .B2(new_n662), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n670), .A2(new_n666), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT84), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n670), .A3(new_n666), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G35), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G162), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G2090), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT92), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(G27), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G164), .B2(new_n681), .ZN(new_n688));
  INV_X1    g263(.A(G2078), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G4), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n595), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT87), .B(G1348), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n684), .A2(G2090), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(G21), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G168), .B2(new_n691), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(G1966), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(G1966), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n686), .A2(new_n690), .A3(new_n695), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(G19), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n543), .B2(new_n691), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT88), .B(G1341), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n681), .A2(G33), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT25), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n487), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n459), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n709), .B(new_n711), .C1(G139), .C2(new_n475), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n707), .B1(new_n712), .B2(new_n681), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2072), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n620), .A2(new_n681), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT30), .B(G28), .ZN(new_n716));
  OR2_X1    g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  NAND2_X1  g292(.A1(KEYINPUT31), .A2(G11), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n716), .A2(new_n681), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n706), .A2(new_n714), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n691), .A2(G5), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G171), .B2(new_n691), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n681), .B1(new_n725), .B2(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G160), .B2(G29), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n724), .B1(G2084), .B2(new_n728), .C1(G2072), .C2(new_n713), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n475), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n478), .A2(G129), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  NAND3_X1  g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(new_n681), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT91), .B1(G29), .B2(G32), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n728), .A2(G2084), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT90), .Z(new_n743));
  NOR4_X1   g318(.A1(new_n720), .A2(new_n729), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G299), .A2(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n691), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT93), .B(G1956), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n681), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n475), .A2(G140), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n478), .A2(G128), .ZN(new_n755));
  OR2_X1    g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(new_n681), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT89), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n744), .A2(new_n751), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n749), .A2(new_n750), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n702), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT95), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n691), .A2(G22), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G166), .B2(new_n691), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1971), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT33), .B(G1976), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G23), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT85), .Z(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G288), .B2(new_n691), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n769), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  MUX2_X1   g349(.A(G6), .B(G305), .S(G16), .Z(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n774), .B(new_n777), .C1(new_n770), .C2(new_n773), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT34), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(KEYINPUT34), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n691), .A2(G24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n584), .B2(new_n691), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1986), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n475), .A2(G131), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n478), .A2(G119), .ZN(new_n785));
  OR2_X1    g360(.A1(G95), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G25), .B(new_n788), .S(G29), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT35), .B(G1991), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n779), .A2(new_n780), .A3(new_n783), .A4(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT86), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT86), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n793), .A2(KEYINPUT36), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(KEYINPUT36), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n766), .A2(new_n795), .A3(new_n796), .ZN(G311));
  NAND3_X1  g372(.A1(new_n766), .A2(new_n795), .A3(new_n796), .ZN(G150));
  AOI22_X1  g373(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n507), .ZN(new_n800));
  INV_X1    g375(.A(G55), .ZN(new_n801));
  INV_X1    g376(.A(G93), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n510), .A2(new_n801), .B1(new_n516), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT97), .Z(new_n805));
  INV_X1    g380(.A(G860), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT37), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n594), .A2(new_n602), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n542), .A2(new_n804), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n805), .A2(new_n542), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n810), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n806), .B1(new_n817), .B2(KEYINPUT39), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n808), .B1(new_n818), .B2(new_n819), .ZN(G145));
  XOR2_X1   g395(.A(new_n610), .B(new_n788), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n475), .A2(G142), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT99), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n478), .A2(G130), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n459), .A2(G118), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n821), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n759), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n712), .B(new_n734), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n499), .A2(KEYINPUT98), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n490), .A2(new_n832), .A3(new_n498), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n830), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n829), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n620), .B(G160), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G162), .ZN(new_n838));
  AOI21_X1  g413(.A(G37), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n836), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g416(.A(KEYINPUT101), .B1(new_n805), .B2(G868), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n815), .B(new_n605), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n594), .A2(G299), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n594), .A2(G299), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n846), .A2(KEYINPUT41), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(KEYINPUT41), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n847), .B1(new_n850), .B2(new_n843), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT100), .ZN(new_n852));
  XOR2_X1   g427(.A(G303), .B(G288), .Z(new_n853));
  XNOR2_X1  g428(.A(G305), .B(new_n584), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT42), .Z(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n851), .B2(KEYINPUT100), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n598), .B1(new_n852), .B2(new_n857), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n842), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(G295));
  AOI21_X1  g438(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(G331));
  XNOR2_X1  g439(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n866));
  XNOR2_X1  g441(.A(G168), .B(G301), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n815), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n868), .A2(new_n846), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n813), .A2(new_n814), .ZN(new_n870));
  INV_X1    g445(.A(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(KEYINPUT103), .A3(new_n871), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n875), .A2(new_n876), .B1(new_n815), .B2(new_n867), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n855), .B(new_n873), .C1(new_n877), .C2(new_n850), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n873), .B1(new_n877), .B2(new_n850), .ZN(new_n881));
  INV_X1    g456(.A(new_n855), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n866), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n850), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n872), .A2(new_n868), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n875), .A2(new_n876), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n885), .A2(new_n886), .B1(new_n887), .B2(new_n869), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n878), .B(new_n879), .C1(new_n888), .C2(new_n855), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n865), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n883), .A2(new_n879), .A3(new_n878), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n892), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(G397));
  XNOR2_X1  g470(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n834), .B2(G1384), .ZN(new_n897));
  INV_X1    g472(.A(G40), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n464), .A2(new_n468), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G1996), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n734), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT105), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n758), .B(G2067), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(G1996), .B2(new_n734), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n897), .A2(new_n900), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n788), .B(new_n790), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT106), .Z(new_n913));
  OAI211_X1 g488(.A(new_n905), .B(new_n911), .C1(new_n909), .C2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n584), .B(G1986), .Z(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n901), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT63), .ZN(new_n917));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n831), .A2(KEYINPUT45), .A3(new_n918), .A4(new_n833), .ZN(new_n919));
  AOI21_X1  g494(.A(G1384), .B1(new_n500), .B2(new_n502), .ZN(new_n920));
  INV_X1    g495(.A(new_n896), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n899), .B(new_n919), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1971), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(G1384), .B1(new_n490), .B2(new_n498), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n899), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n490), .A2(new_n501), .A3(new_n498), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n501), .B1(new_n490), .B2(new_n498), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n927), .B1(new_n931), .B2(KEYINPUT109), .ZN(new_n932));
  INV_X1    g507(.A(G2090), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n503), .A2(new_n934), .A3(new_n928), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G8), .ZN(new_n938));
  NAND2_X1  g513(.A1(G303), .A2(G8), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI211_X1 g516(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n498), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n918), .B1(new_n929), .B2(new_n930), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n900), .B(new_n942), .C1(new_n943), .C2(KEYINPUT50), .ZN(new_n944));
  INV_X1    g519(.A(G2084), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n899), .B1(new_n925), .B2(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT110), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n948), .B(new_n899), .C1(new_n925), .C2(KEYINPUT45), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n918), .B(new_n921), .C1(new_n929), .C2(new_n930), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1966), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n944), .A2(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n954), .A3(G286), .ZN(new_n955));
  INV_X1    g530(.A(new_n942), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n900), .A2(G2090), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n956), .B(new_n957), .C1(new_n920), .C2(new_n926), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n942), .B1(new_n943), .B2(KEYINPUT50), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(KEYINPUT107), .A3(new_n957), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n924), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n940), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(G8), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n499), .A2(new_n899), .A3(new_n918), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G8), .ZN(new_n967));
  INV_X1    g542(.A(G1976), .ZN(new_n968));
  NOR2_X1   g543(.A1(G288), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT52), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n954), .B1(new_n925), .B2(new_n899), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n968), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n971), .B(new_n972), .C1(new_n968), .C2(G288), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n975));
  INV_X1    g550(.A(G1981), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n573), .A2(new_n576), .A3(new_n577), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G86), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n568), .B1(new_n516), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(G1981), .B1(new_n979), .B2(new_n572), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n967), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(KEYINPUT49), .A3(new_n980), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n975), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n984), .A3(new_n971), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT108), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n974), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n941), .A2(new_n955), .A3(new_n965), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n917), .B1(new_n990), .B2(KEYINPUT111), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n963), .A2(G8), .A3(new_n964), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n954), .B1(new_n924), .B2(new_n936), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n989), .B1(new_n994), .B2(new_n964), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n996), .B2(new_n955), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT112), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n992), .A3(new_n955), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n990), .A2(KEYINPUT111), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n917), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n955), .A2(KEYINPUT63), .A3(new_n989), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n964), .B1(new_n963), .B2(G8), .ZN(new_n1004));
  OR3_X1    g579(.A1(new_n1003), .A2(new_n993), .A3(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n998), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(G1976), .B(G288), .C1(new_n985), .C2(new_n988), .ZN(new_n1007));
  INV_X1    g582(.A(new_n977), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n971), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n974), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n983), .B1(new_n982), .B2(new_n984), .ZN(new_n1011));
  AND4_X1   g586(.A1(new_n983), .A2(new_n986), .A3(new_n984), .A4(new_n971), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1009), .B1(new_n965), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n943), .A2(new_n896), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1015), .A2(new_n689), .A3(new_n899), .A4(new_n919), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n956), .B(new_n899), .C1(new_n920), .C2(new_n926), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1016), .A2(new_n1017), .B1(new_n1018), .B2(new_n723), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n689), .A2(KEYINPUT53), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n951), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G301), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n941), .A2(new_n965), .A3(new_n1022), .A4(new_n989), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT51), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n951), .A2(new_n952), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n961), .A2(new_n945), .A3(new_n899), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n954), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G168), .A2(new_n954), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT120), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1025), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1029), .B(KEYINPUT120), .Z(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1032), .B(new_n1033), .C1(new_n953), .C2(new_n954), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n953), .A2(new_n1032), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT62), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1023), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1014), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n694), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n961), .B2(new_n899), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n966), .A2(G2067), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1043), .A2(KEYINPUT115), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1018), .B2(new_n694), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT60), .B(new_n594), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT61), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G299), .A2(KEYINPUT113), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT57), .Z(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(G2072), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1015), .A2(new_n899), .A3(new_n919), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1956), .B1(new_n932), .B2(new_n935), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1052), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1051), .B(KEYINPUT57), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n932), .A2(new_n935), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1062), .B2(new_n1055), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1050), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1015), .A2(new_n902), .A3(new_n899), .A4(new_n919), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(G1341), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n966), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n542), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1069), .A2(KEYINPUT59), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1062), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1071), .A2(KEYINPUT61), .B1(KEYINPUT59), .B2(new_n1069), .ZN(new_n1072));
  AND4_X1   g647(.A1(new_n1049), .A2(new_n1064), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT60), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT115), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n595), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1062), .A2(new_n1080), .A3(new_n1055), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1052), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT118), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1075), .A2(new_n1076), .A3(new_n595), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1081), .A2(new_n1082), .A3(new_n1087), .A4(new_n1052), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1075), .A2(new_n1076), .A3(new_n1089), .A4(new_n595), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1073), .A2(new_n1079), .B1(new_n1091), .B2(new_n1071), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1017), .B1(new_n922), .B2(G2078), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1018), .A2(new_n723), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT53), .B1(new_n1095), .B2(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1095), .B2(G2078), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n897), .A2(new_n899), .A3(new_n919), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G171), .B(KEYINPUT54), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1100), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1019), .A2(new_n1102), .A3(new_n1021), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1013), .B1(new_n938), .B2(new_n940), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n965), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1036), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n996), .A2(new_n1039), .A3(new_n1108), .A4(new_n1104), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1041), .B1(new_n1092), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n916), .B1(new_n1006), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n788), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n905), .A2(new_n790), .A3(new_n1113), .A4(new_n911), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n758), .A2(G2067), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1114), .A2(KEYINPUT124), .A3(new_n1116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n901), .A3(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n909), .A2(G1986), .A3(G290), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT48), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n914), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n901), .B1(new_n734), .B2(new_n907), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n903), .A2(KEYINPUT46), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n903), .A2(KEYINPUT46), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1128), .A2(KEYINPUT126), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(KEYINPUT126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1124), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1121), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1112), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g713(.A1(G227), .A2(new_n457), .ZN(new_n1140));
  NOR2_X1   g714(.A1(G229), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g715(.A1(new_n639), .A2(new_n1141), .A3(new_n840), .ZN(new_n1142));
  NAND2_X1  g716(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n1143));
  OR2_X1    g717(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n1144));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(G308));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1143), .ZN(new_n1146));
  NAND4_X1  g720(.A1(new_n1146), .A2(new_n639), .A3(new_n840), .A4(new_n1141), .ZN(G225));
endmodule


