//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n232), .A2(G20), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n213), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n252), .B(new_n253), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT75), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT10), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n202), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n208), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G58), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(KEYINPUT72), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT8), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n258), .B1(new_n259), .B2(new_n261), .C1(new_n262), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n230), .A2(new_n231), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n230), .A2(new_n270), .A3(new_n231), .A4(new_n267), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n207), .B2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n270), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n272), .A2(new_n274), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n257), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G223), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n287), .B1(new_n221), .B2(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n232), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(G1), .A2(G13), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n291), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n207), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G226), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n298), .B2(new_n291), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n207), .C1(G41), .C2(G45), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n294), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G190), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(G200), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n256), .A2(KEYINPUT10), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n277), .A2(new_n278), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n280), .A2(new_n314), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n277), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n310), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G179), .B2(new_n310), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n317), .A2(new_n312), .A3(new_n313), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n315), .B1(new_n323), .B2(new_n279), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n261), .A2(new_n273), .B1(new_n208), .B2(G68), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n262), .A2(new_n221), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n268), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT11), .ZN(new_n329));
  OAI21_X1  g0129(.A(G68), .B1(new_n208), .B2(G1), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n328), .A2(new_n329), .B1(new_n271), .B2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n328), .A2(new_n329), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n270), .A2(G68), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT12), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n285), .A2(G226), .A3(new_n286), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n282), .A2(new_n284), .A3(G232), .A4(G1698), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n293), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n297), .A2(G238), .A3(new_n299), .A4(new_n300), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n342), .A2(new_n308), .A3(KEYINPUT76), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT76), .B1(new_n342), .B2(new_n308), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT13), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n341), .B(new_n347), .C1(new_n344), .C2(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(G169), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n346), .A2(G179), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n350), .B1(new_n349), .B2(G169), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n336), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT77), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT77), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n346), .A2(new_n358), .A3(G190), .A4(new_n348), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n349), .A2(G200), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n335), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  XNOR2_X1  g0164(.A(G58), .B(G68), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n283), .A2(KEYINPUT78), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT78), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n369), .A3(G33), .ZN(new_n370));
  AOI21_X1  g0170(.A(G20), .B1(new_n370), .B2(new_n282), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  OAI21_X1  g0172(.A(G68), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n282), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(G33), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT79), .B(KEYINPUT7), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n376), .A2(G20), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT16), .B(new_n366), .C1(new_n373), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n366), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n284), .B1(new_n375), .B2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n372), .A2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n377), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n285), .B2(G20), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n380), .B1(new_n386), .B2(G68), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n379), .B(new_n268), .C1(new_n387), .C2(KEYINPUT16), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n265), .B1(new_n207), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n272), .B1(new_n275), .B2(new_n265), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  MUX2_X1   g0191(.A(G223), .B(G226), .S(G1698), .Z(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(new_n370), .A3(new_n282), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G87), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n292), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n297), .A2(G232), .A3(new_n299), .A4(new_n300), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n308), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n395), .A2(new_n397), .A3(G179), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n396), .A2(new_n308), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT80), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n393), .A2(new_n394), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n399), .B(new_n400), .C1(new_n401), .C2(new_n292), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT80), .B1(new_n395), .B2(new_n397), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n398), .B1(new_n404), .B2(new_n320), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n364), .B1(new_n391), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n395), .A2(new_n397), .A3(G190), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n388), .A4(new_n390), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n391), .A2(new_n405), .A3(new_n364), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n388), .B(new_n390), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n407), .A2(new_n411), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n285), .A2(G232), .A3(new_n286), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n417), .B1(new_n223), .B2(new_n285), .C1(new_n288), .C2(new_n216), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n293), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n301), .A2(G244), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n308), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n320), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT15), .B(G87), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n262), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT8), .B(G58), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n261), .B1(new_n208), .B2(new_n221), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(KEYINPUT73), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(KEYINPUT73), .B2(new_n426), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n268), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n221), .B1(new_n207), .B2(G20), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n272), .A2(new_n430), .B1(new_n221), .B2(new_n275), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n420), .A2(new_n308), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n418), .B2(new_n293), .ZN(new_n434));
  INV_X1    g0234(.A(G179), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n422), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT74), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n421), .A2(G200), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(G190), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n432), .A2(new_n438), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n437), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n325), .A2(new_n363), .A3(new_n416), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G116), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT84), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G116), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(new_n270), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n281), .A2(G1), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n271), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(new_n449), .A3(G20), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(G33), .B2(G283), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n281), .A2(G97), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n268), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT20), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT84), .B(G116), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(G20), .B1(new_n456), .B2(new_n455), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n268), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n451), .B(new_n453), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(G257), .A2(G1698), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n224), .B2(G1698), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n370), .A3(new_n282), .ZN(new_n467));
  XOR2_X1   g0267(.A(KEYINPUT87), .B(G303), .Z(new_n468));
  NAND2_X1  g0268(.A1(new_n282), .A2(new_n284), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n292), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n207), .B(G45), .C1(new_n472), .C2(KEYINPUT5), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G41), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(KEYINPUT5), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n474), .A2(new_n304), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n299), .B(G270), .C1(new_n473), .C2(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n471), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G190), .ZN(new_n485));
  OAI21_X1  g0285(.A(G200), .B1(new_n471), .B2(new_n483), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n464), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT89), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n464), .A2(new_n485), .A3(KEYINPUT89), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n467), .A2(new_n470), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n293), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n481), .A2(new_n482), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(G169), .B1(new_n471), .B2(new_n483), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n435), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n453), .ZN(new_n500));
  INV_X1    g0300(.A(new_n451), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT20), .B1(new_n462), .B2(new_n268), .ZN(new_n502));
  AND4_X1   g0302(.A1(KEYINPUT20), .A2(new_n268), .A3(new_n457), .A4(new_n454), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT88), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n320), .B1(new_n494), .B2(new_n495), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n504), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(new_n498), .ZN(new_n509));
  AOI211_X1 g0309(.A(KEYINPUT88), .B(KEYINPUT21), .C1(new_n507), .C2(new_n504), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT90), .B1(new_n492), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n498), .B1(new_n464), .B2(new_n497), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n506), .A3(new_n498), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT90), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n491), .A3(new_n517), .A4(new_n505), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n474), .A2(new_n478), .B1(new_n298), .B2(new_n291), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G257), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n481), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n370), .A2(G244), .A3(new_n286), .A4(new_n282), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT4), .A2(G244), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n282), .A2(new_n284), .A3(new_n526), .A4(new_n286), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n292), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n524), .B2(new_n523), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT81), .B1(new_n535), .B2(new_n292), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n522), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G200), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT83), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n481), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(G257), .B2(new_n520), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n531), .A2(new_n532), .ZN(new_n542));
  AOI211_X1 g0342(.A(KEYINPUT81), .B(new_n292), .C1(new_n525), .C2(new_n530), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(G200), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n223), .B1(new_n383), .B2(new_n385), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n548), .A2(new_n549), .A3(G107), .ZN(new_n550));
  XNOR2_X1  g0350(.A(G97), .B(G107), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n552), .A2(new_n208), .B1(new_n221), .B2(new_n261), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n268), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n270), .A2(G97), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n271), .A2(new_n452), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n531), .A2(new_n522), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(G190), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n539), .A2(new_n546), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n435), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n541), .B1(new_n292), .B2(new_n535), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n320), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n564), .A3(new_n558), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n268), .ZN(new_n567));
  XOR2_X1   g0367(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n568));
  NAND2_X1  g0368(.A1(new_n370), .A2(new_n282), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT22), .ZN(new_n570));
  NOR4_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(G20), .A4(new_n217), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n208), .A2(G87), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n469), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n450), .A2(new_n208), .A3(G33), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT92), .B1(new_n223), .B2(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT23), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n575), .A2(KEYINPUT23), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n573), .A2(new_n574), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n568), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n574), .A2(new_n577), .A3(new_n576), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n376), .A2(KEYINPUT22), .A3(new_n208), .A4(G87), .ZN(new_n581));
  INV_X1    g0381(.A(new_n568), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n573), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n567), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT93), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT25), .ZN(new_n586));
  AOI211_X1 g0386(.A(G107), .B(new_n270), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n589), .A2(new_n590), .B1(new_n556), .B2(G107), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n520), .A2(G264), .ZN(new_n594));
  MUX2_X1   g0394(.A(G250), .B(G257), .S(G1698), .Z(new_n595));
  AOI22_X1  g0395(.A1(new_n376), .A2(new_n595), .B1(G33), .B2(G294), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n481), .B(new_n594), .C1(new_n596), .C2(new_n292), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G190), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(G200), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n435), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n320), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n602), .B(new_n603), .C1(new_n584), .C2(new_n592), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n207), .A2(new_n303), .A3(G45), .ZN(new_n605));
  INV_X1    g0405(.A(G45), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n218), .B1(new_n606), .B2(G1), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n299), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(G238), .A2(G1698), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n222), .B2(G1698), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n370), .A3(new_n282), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n450), .A2(G33), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n614), .B2(new_n293), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n435), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n338), .B2(new_n208), .ZN(new_n618));
  NOR4_X1   g0418(.A1(KEYINPUT85), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  NOR2_X1   g0420(.A1(G87), .A2(G97), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n223), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n618), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n370), .A2(new_n208), .A3(G68), .A4(new_n282), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n617), .B1(new_n262), .B2(new_n549), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n268), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n423), .A2(new_n275), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n452), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n567), .A2(new_n270), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT86), .B1(new_n631), .B2(new_n423), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT86), .ZN(new_n633));
  INV_X1    g0433(.A(new_n423), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n556), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  OAI221_X1 g0436(.A(new_n616), .B1(G169), .B2(new_n615), .C1(new_n629), .C2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n626), .A2(new_n268), .B1(new_n275), .B2(new_n423), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n556), .A2(G87), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n615), .A2(G190), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n640), .B(new_n641), .C1(new_n538), .C2(new_n615), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n601), .A2(new_n604), .A3(new_n637), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n566), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n445), .A2(new_n519), .A3(new_n644), .ZN(G372));
  NAND2_X1  g0445(.A1(new_n361), .A2(new_n335), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n359), .B2(new_n357), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n355), .B1(new_n647), .B2(new_n437), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n413), .B(KEYINPUT17), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n391), .A2(new_n405), .A3(new_n364), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n406), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n324), .A3(new_n318), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n322), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT96), .B1(new_n516), .B2(new_n505), .ZN(new_n656));
  OAI211_X1 g0456(.A(KEYINPUT96), .B(new_n505), .C1(new_n509), .C2(new_n510), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n604), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT94), .B1(new_n614), .B2(new_n293), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT94), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n661), .B(new_n292), .C1(new_n612), .C2(new_n613), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n608), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n320), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT95), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n632), .A2(new_n635), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n666), .A2(new_n638), .B1(new_n435), .B2(new_n615), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT95), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n663), .A2(new_n668), .A3(new_n320), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n641), .A2(new_n638), .A3(new_n639), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(G200), .B2(new_n663), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n601), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n566), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n659), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n562), .A2(new_n564), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT98), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n562), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n558), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n670), .A2(new_n673), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n677), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n642), .A2(new_n637), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n685), .A2(new_n677), .A3(new_n565), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT97), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n670), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n616), .B1(new_n629), .B2(new_n636), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n664), .B2(KEYINPUT95), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT97), .A3(new_n669), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n676), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n445), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n655), .A2(new_n696), .ZN(G369));
  NAND3_X1  g0497(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n464), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n512), .B2(new_n518), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT96), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n511), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(new_n657), .A3(new_n705), .ZN(new_n709));
  OAI21_X1  g0509(.A(G330), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n604), .A2(new_n703), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n601), .B1(new_n593), .B2(new_n704), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n604), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n511), .A2(new_n704), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n604), .B2(new_n703), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT99), .ZN(G399));
  INV_X1    g0522(.A(KEYINPUT100), .ZN(new_n723));
  INV_X1    g0523(.A(new_n211), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(G41), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n211), .A2(KEYINPUT100), .A3(new_n472), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G1), .ZN(new_n728));
  OR3_X1    g0528(.A1(new_n619), .A2(new_n622), .A3(G116), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n728), .A2(new_n729), .B1(new_n233), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n376), .A2(new_n611), .B1(G33), .B2(new_n450), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n608), .B1(new_n732), .B2(new_n292), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n594), .B1(new_n596), .B2(new_n292), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n563), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT101), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n484), .A2(new_n736), .A3(G179), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT101), .B1(new_n496), .B2(new_n435), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n598), .A2(G179), .A3(new_n484), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n544), .A3(new_n663), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n734), .A2(new_n733), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n738), .A2(new_n742), .A3(new_n737), .A4(new_n559), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n746), .B2(new_n703), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT102), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n703), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT102), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n519), .A2(new_n644), .A3(new_n704), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n749), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT29), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n561), .A2(new_n565), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n672), .B1(new_n692), .B2(new_n669), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n516), .A2(new_n505), .A3(new_n604), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n761), .A2(new_n601), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n685), .A2(KEYINPUT26), .A3(new_n565), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n690), .A2(new_n693), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(KEYINPUT103), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT103), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n690), .A2(new_n768), .A3(new_n693), .ZN(new_n769));
  INV_X1    g0569(.A(new_n558), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n678), .B2(new_n679), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n762), .A2(new_n681), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT26), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n764), .A2(new_n767), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n760), .B1(new_n774), .B2(new_n704), .ZN(new_n775));
  INV_X1    g0575(.A(new_n604), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n708), .B2(new_n657), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n762), .A2(new_n565), .A3(new_n561), .A4(new_n601), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n694), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n686), .B1(new_n772), .B2(new_n677), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n760), .B(new_n704), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n759), .A2(new_n775), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n731), .B1(new_n783), .B2(G1), .ZN(G364));
  INV_X1    g0584(.A(new_n727), .ZN(new_n785));
  INV_X1    g0585(.A(G13), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n207), .B1(new_n787), .B2(G45), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n711), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n706), .A2(new_n709), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(G330), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n232), .B1(new_n208), .B2(G169), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n208), .A2(new_n435), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(new_n356), .A3(G200), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  OAI221_X1 g0601(.A(new_n469), .B1(new_n798), .B2(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n208), .A2(G179), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n803), .A2(new_n797), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT104), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT104), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n802), .B1(new_n808), .B2(G329), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n803), .A2(G190), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT105), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G303), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n356), .A2(G179), .A3(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n208), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n803), .A2(new_n356), .A3(G200), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n819), .A2(G294), .B1(new_n821), .B2(G283), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n796), .A2(G190), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G200), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n538), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G322), .A2(new_n824), .B1(new_n825), .B2(G326), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n809), .A2(new_n816), .A3(new_n822), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G159), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n807), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT32), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n815), .A2(G87), .ZN(new_n831));
  INV_X1    g0631(.A(new_n825), .ZN(new_n832));
  INV_X1    g0632(.A(new_n824), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n273), .A2(new_n832), .B1(new_n833), .B2(new_n263), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n285), .B1(new_n798), .B2(new_n221), .C1(new_n215), .C2(new_n800), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n818), .A2(new_n549), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n820), .A2(new_n223), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n830), .A2(new_n831), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n827), .B1(new_n840), .B2(KEYINPUT106), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT106), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n795), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n790), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n724), .A2(new_n376), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n606), .B2(new_n234), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n606), .B2(new_n254), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n724), .A2(new_n469), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n850), .A2(G355), .B1(new_n446), .B2(new_n724), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(G13), .A2(G33), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(G20), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n795), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n845), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n855), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n844), .B(new_n857), .C1(new_n792), .C2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n793), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G396));
  NOR2_X1   g0661(.A1(new_n795), .A2(new_n853), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n790), .B1(G77), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(G303), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n832), .A2(new_n865), .B1(new_n820), .B2(new_n217), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n836), .B(new_n866), .C1(G294), .C2(new_n824), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n815), .A2(G107), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n808), .A2(G311), .ZN(new_n869));
  INV_X1    g0669(.A(G283), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n469), .B1(new_n800), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n798), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n450), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n800), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n875), .A2(G150), .B1(new_n872), .B2(G159), .ZN(new_n876));
  INV_X1    g0676(.A(G143), .ZN(new_n877));
  INV_X1    g0677(.A(G137), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n876), .B1(new_n833), .B2(new_n877), .C1(new_n878), .C2(new_n832), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT34), .Z(new_n880));
  NOR2_X1   g0680(.A1(new_n820), .A2(new_n215), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n569), .B(new_n881), .C1(G58), .C2(new_n819), .ZN(new_n882));
  INV_X1    g0682(.A(G132), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n882), .B1(new_n273), .B2(new_n814), .C1(new_n883), .C2(new_n807), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n874), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n864), .B1(new_n885), .B2(new_n795), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n437), .A2(new_n703), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n442), .A2(new_n443), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n704), .B1(new_n429), .B2(new_n431), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n437), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n886), .B1(new_n894), .B2(new_n854), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n695), .B2(new_n704), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n444), .A2(new_n703), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n779), .B2(new_n780), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT107), .B(new_n897), .C1(new_n779), .C2(new_n780), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n759), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n845), .B1(new_n902), .B2(new_n759), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(G384));
  NAND3_X1  g0706(.A1(new_n232), .A2(G20), .A3(G116), .ZN(new_n907));
  INV_X1    g0707(.A(new_n552), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(KEYINPUT35), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(KEYINPUT35), .B2(new_n908), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT36), .ZN(new_n911));
  OAI21_X1  g0711(.A(G77), .B1(new_n263), .B2(new_n215), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n912), .A2(new_n233), .B1(G50), .B2(new_n215), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(G1), .A3(new_n786), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT108), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n379), .A2(new_n268), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n371), .A2(new_n384), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(G68), .C1(new_n372), .C2(new_n371), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT16), .B1(new_n920), .B2(new_n366), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n390), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n701), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n416), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n405), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n924), .A3(new_n413), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n391), .A2(new_n405), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n391), .A2(new_n923), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT37), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n413), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n926), .A2(new_n934), .A3(KEYINPUT38), .ZN(new_n935));
  INV_X1    g0735(.A(new_n931), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n416), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n931), .A3(new_n413), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT37), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n933), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n917), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n354), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n352), .A3(new_n351), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n336), .A3(new_n704), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT109), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT38), .ZN(new_n947));
  INV_X1    g0747(.A(new_n934), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n924), .B1(new_n649), .B2(new_n652), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n926), .A2(new_n934), .A3(KEYINPUT38), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n942), .B(new_n946), .C1(new_n917), .C2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n701), .B1(new_n651), .B2(new_n406), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT107), .B1(new_n695), .B2(new_n897), .ZN(new_n957));
  INV_X1    g0757(.A(new_n901), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n888), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n336), .B(new_n703), .C1(new_n647), .C2(new_n944), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n336), .A2(new_n703), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n355), .A2(new_n362), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n952), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n445), .B1(new_n775), .B2(new_n782), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n655), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n965), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(G330), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n747), .A2(new_n748), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n756), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n893), .B1(new_n960), .B2(new_n962), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n935), .C2(new_n941), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT40), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT40), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n952), .A2(new_n975), .A3(new_n971), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n445), .A2(new_n971), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n969), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n978), .B2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n968), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n207), .B2(new_n787), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n968), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n916), .B1(new_n982), .B2(new_n983), .ZN(G367));
  OAI21_X1  g0784(.A(new_n761), .B1(new_n770), .B2(new_n704), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n771), .A2(new_n681), .A3(new_n703), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n718), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT42), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n987), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n565), .B1(new_n992), .B2(new_n604), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n704), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n640), .A2(new_n704), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n683), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n766), .B2(new_n996), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT43), .B1(new_n999), .B2(KEYINPUT110), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(KEYINPUT110), .B2(new_n999), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n995), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n995), .B2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n715), .A2(new_n992), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n727), .B(KEYINPUT41), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT111), .B1(new_n714), .B2(new_n717), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n711), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n710), .B(KEYINPUT111), .C1(new_n714), .C2(new_n717), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1009), .A2(new_n1010), .A3(new_n988), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n988), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n775), .A2(new_n782), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n758), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT112), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n720), .B2(new_n987), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n992), .A2(KEYINPUT44), .A3(new_n719), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n720), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT45), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n992), .B2(new_n719), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1020), .A2(new_n715), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n715), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n718), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1009), .A2(new_n1010), .A3(new_n988), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT112), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n783), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1016), .A2(new_n1027), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1007), .B1(new_n1034), .B2(new_n783), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1006), .B1(new_n1035), .B2(new_n789), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n246), .A2(new_n847), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n856), .B1(new_n211), .B2(new_n423), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n790), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n800), .A2(new_n828), .B1(new_n798), .B2(new_n273), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n877), .A2(new_n832), .B1(new_n833), .B2(new_n259), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G68), .C2(new_n819), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n808), .A2(G137), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n820), .A2(new_n221), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT113), .B1(new_n1044), .B2(new_n469), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT113), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1044), .A2(new_n469), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n815), .A2(G58), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT46), .B1(new_n815), .B2(new_n450), .ZN(new_n1050));
  INV_X1    g0850(.A(G294), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n800), .A2(new_n1051), .B1(new_n798), .B2(new_n870), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n376), .B(new_n1052), .C1(new_n808), .C2(G317), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n815), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n819), .A2(G107), .B1(new_n821), .B2(G97), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G311), .A2(new_n825), .B1(new_n824), .B2(new_n468), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1049), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT47), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1039), .B1(new_n1060), .B2(new_n795), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n999), .B2(new_n858), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1036), .A2(new_n1062), .ZN(G387));
  NAND2_X1  g0863(.A1(new_n1016), .A2(new_n1033), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n727), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n242), .A2(new_n606), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(new_n846), .B1(new_n729), .B2(new_n850), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n425), .A2(G50), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n606), .B1(new_n215), .B2(new_n221), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n729), .B(new_n1071), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1068), .A2(new_n1072), .B1(G107), .B2(new_n211), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n845), .B1(new_n1073), .B2(new_n856), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n714), .B2(new_n858), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n832), .A2(new_n828), .B1(new_n820), .B2(new_n549), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n569), .B(new_n1076), .C1(G68), .C2(new_n872), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n818), .A2(new_n423), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n265), .A2(new_n800), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G50), .C2(new_n824), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n808), .A2(G150), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n814), .A2(new_n221), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G322), .A2(new_n825), .B1(new_n875), .B2(G311), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n824), .A2(G317), .B1(new_n872), .B2(new_n468), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT48), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n814), .A2(new_n1051), .B1(new_n870), .B2(new_n818), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n808), .A2(G326), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n376), .B1(new_n450), .B2(new_n821), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT49), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1084), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1075), .B1(new_n795), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n1031), .B2(new_n789), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1066), .A2(new_n1101), .ZN(G393));
  OAI21_X1  g0902(.A(new_n1064), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n785), .A3(new_n1034), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n992), .A2(new_n855), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n251), .A2(new_n847), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n856), .B1(new_n549), .B2(new_n211), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n790), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n569), .B1(G87), .B2(new_n821), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(new_n814), .B2(new_n215), .C1(new_n807), .C2(new_n877), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT117), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G150), .A2(new_n825), .B1(new_n824), .B2(G159), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT51), .Z(new_n1113));
  OAI22_X1  g0913(.A1(new_n800), .A2(new_n273), .B1(new_n798), .B2(new_n425), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G77), .B2(new_n819), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G311), .A2(new_n824), .B1(new_n825), .B2(G317), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n468), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n469), .B1(new_n798), .B2(new_n1051), .C1(new_n1119), .C2(new_n800), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n837), .B(new_n1120), .C1(new_n450), .C2(new_n819), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n808), .A2(G322), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n870), .C2(new_n814), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1108), .B1(new_n1124), .B2(new_n795), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1027), .A2(new_n789), .B1(new_n1105), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1104), .A2(new_n1126), .ZN(G390));
  AOI21_X1  g0927(.A(new_n969), .B1(new_n756), .B2(new_n970), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n445), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n966), .A2(new_n655), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n757), .A2(G330), .A3(new_n894), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n963), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n972), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n959), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1128), .A2(new_n894), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1132), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n757), .A2(G330), .A3(new_n894), .A4(new_n963), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n891), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n437), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n764), .A2(new_n773), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n766), .A2(KEYINPUT103), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n765), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n769), .A3(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n704), .B(new_n1141), .C1(new_n1142), .C2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1138), .A2(new_n888), .A3(new_n1139), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1130), .B1(new_n1136), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n946), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n887), .B1(new_n900), .B2(new_n901), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n1132), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n942), .B1(new_n952), .B2(new_n917), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1146), .A2(new_n888), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n963), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n935), .A2(new_n941), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n946), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1134), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1132), .B1(new_n1146), .B2(new_n888), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1150), .B1(new_n935), .B2(new_n941), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1139), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1149), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1139), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n946), .B1(new_n959), .B2(new_n963), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1153), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1152), .A2(new_n1153), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1148), .B(new_n1170), .C1(new_n1171), .C2(new_n1134), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1165), .A2(new_n785), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n845), .B1(new_n265), .B2(new_n862), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n469), .B1(new_n798), .B2(new_n549), .C1(new_n223), .C2(new_n800), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n446), .A2(new_n833), .B1(new_n832), .B2(new_n870), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n818), .A2(new_n221), .ZN(new_n1177));
  OR3_X1    g0977(.A1(new_n1176), .A2(new_n881), .A3(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(G294), .C2(new_n808), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n814), .A2(new_n259), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT53), .ZN(new_n1181));
  INV_X1    g0981(.A(G125), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n285), .B1(new_n828), .B2(new_n818), .C1(new_n807), .C2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT54), .B(G143), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n800), .A2(new_n878), .B1(new_n798), .B2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT118), .Z(new_n1186));
  NOR2_X1   g0986(.A1(new_n820), .A2(new_n273), .ZN(new_n1187));
  INV_X1    g0987(.A(G128), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1188), .A2(new_n832), .B1(new_n833), .B2(new_n883), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1183), .A2(new_n1186), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1179), .A2(new_n831), .B1(new_n1181), .B2(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1174), .B1(new_n794), .B2(new_n1191), .C1(new_n1169), .C2(new_n854), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1170), .A2(new_n789), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1160), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT119), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1170), .B(new_n789), .C1(new_n1171), .C2(new_n1134), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT119), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n1192), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1173), .A2(new_n1195), .A3(new_n1198), .ZN(G378));
  XNOR2_X1  g0999(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT121), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n325), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n277), .A2(new_n923), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT120), .Z(new_n1204));
  INV_X1    g1004(.A(new_n1201), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n318), .A2(new_n322), .A3(new_n324), .A4(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1202), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1204), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n853), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n472), .B1(new_n798), .B2(new_n423), .C1(new_n549), .C2(new_n800), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n376), .B(new_n1211), .C1(G68), .C2(new_n819), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n870), .B2(new_n807), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G107), .A2(new_n824), .B1(new_n825), .B2(G116), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n263), .B2(new_n820), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1213), .A2(new_n1082), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n472), .B1(new_n375), .B2(new_n281), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1216), .A2(KEYINPUT58), .B1(new_n273), .B2(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n800), .A2(new_n883), .B1(new_n798), .B2(new_n878), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G125), .B2(new_n825), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G150), .A2(new_n819), .B1(new_n824), .B2(G128), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n814), .C2(new_n1184), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n281), .B(new_n472), .C1(new_n820), .C2(new_n828), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n808), .B2(G124), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1218), .B1(KEYINPUT58), .B2(new_n1216), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n795), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n862), .A2(new_n273), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1210), .A2(new_n790), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1209), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n977), .B2(G330), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n969), .B(new_n1209), .C1(new_n974), .C2(new_n976), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n959), .A2(new_n952), .A3(new_n963), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1234), .A2(new_n1235), .B1(new_n1236), .B2(new_n955), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n971), .A2(new_n972), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT40), .B1(new_n950), .B2(new_n951), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(KEYINPUT40), .A2(new_n973), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1209), .B1(new_n1240), .B2(new_n969), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n977), .A2(G330), .A3(new_n1233), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n956), .A4(new_n964), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1237), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1232), .B1(new_n1244), .B2(new_n789), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1159), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1164), .B1(new_n1246), .B2(new_n1135), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1136), .A2(new_n1147), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1130), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(KEYINPUT57), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n785), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1130), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1172), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1244), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1245), .B1(new_n1251), .B2(new_n1254), .ZN(G375));
  OAI21_X1  g1055(.A(new_n790), .B1(G68), .B2(new_n863), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT122), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1078), .A2(new_n1044), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1258), .B1(new_n870), .B2(new_n833), .C1(new_n1051), .C2(new_n832), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n285), .B1(new_n875), .B2(new_n450), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n223), .B2(new_n798), .C1(new_n807), .C2(new_n865), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1259), .B(new_n1261), .C1(G97), .C2(new_n815), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1184), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n875), .A2(new_n1263), .B1(new_n872), .B2(G150), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n376), .B(new_n1264), .C1(new_n807), .C2(new_n1188), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n819), .A2(G50), .B1(new_n821), .B2(G58), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1266), .B1(new_n883), .B2(new_n832), .C1(new_n878), .C2(new_n833), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1265), .B(new_n1267), .C1(G159), .C2(new_n815), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n795), .B1(new_n1262), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1257), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1132), .B2(new_n853), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1248), .B2(new_n789), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT123), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1272), .B(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1007), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1136), .A2(new_n1130), .A3(new_n1147), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1149), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(G381));
  INV_X1    g1078(.A(G390), .ZN(new_n1279));
  INV_X1    g1079(.A(G384), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(G381), .ZN(new_n1283));
  OR4_X1    g1083(.A1(G387), .A2(new_n1283), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1084(.A1(new_n702), .A2(G213), .ZN(new_n1285));
  OR3_X1    g1085(.A1(G375), .A2(G378), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(G407), .A2(G213), .A3(new_n1286), .ZN(G409));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n788), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1007), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1232), .B(new_n1289), .C1(new_n1253), .C2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1288), .B1(new_n1291), .B2(G378), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1245), .C1(new_n1254), .C2(new_n1251), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1198), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1197), .B1(new_n1196), .B2(new_n1192), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1244), .A2(new_n1275), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1245), .B1(new_n1249), .B2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1296), .A2(KEYINPUT124), .A3(new_n1298), .A4(new_n1173), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1292), .A2(new_n1293), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1276), .B1(new_n1148), .B2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n1130), .A4(new_n1147), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n785), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1274), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1280), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1274), .A2(new_n1304), .A3(G384), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1300), .A2(new_n1285), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1300), .A2(new_n1285), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n702), .A2(G213), .A3(G2897), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1306), .A2(new_n1307), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1300), .A2(new_n1319), .A3(new_n1285), .A4(new_n1309), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1311), .A2(new_n1317), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(G387), .A2(KEYINPUT126), .A3(G390), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n860), .B1(new_n1066), .B2(new_n1101), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1281), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1322), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G390), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1036), .A2(KEYINPUT125), .A3(new_n1062), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1324), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G387), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1279), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(G387), .A2(new_n1331), .A3(G390), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1330), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1328), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1321), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT61), .B1(new_n1312), .B2(new_n1316), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1310), .A2(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1285), .A4(new_n1309), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1339), .A2(new_n1341), .A3(new_n1336), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1338), .A2(new_n1343), .ZN(G405));
  INV_X1    g1144(.A(new_n1327), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(new_n1325), .A3(new_n1322), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1293), .A2(new_n1347), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1346), .B(new_n1348), .C1(new_n1349), .C2(new_n1330), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1348), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1351), .B1(new_n1328), .B2(new_n1335), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(G375), .A2(new_n1173), .A3(new_n1296), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1353), .B(new_n1308), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1350), .A2(new_n1352), .A3(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1354), .B1(new_n1350), .B2(new_n1352), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1356), .ZN(G402));
endmodule


