

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790;

  INV_X1 U379 ( .A(n356), .ZN(n721) );
  NAND2_X1 U380 ( .A1(n729), .A2(n383), .ZN(n382) );
  NOR2_X1 U381 ( .A1(n656), .A2(n646), .ZN(n647) );
  INV_X1 U382 ( .A(G237), .ZN(n469) );
  NOR2_X2 U383 ( .A1(G953), .A2(G237), .ZN(n536) );
  NAND2_X1 U384 ( .A1(n581), .A2(n582), .ZN(n356) );
  AND2_X1 U385 ( .A1(n739), .A2(n559), .ZN(n560) );
  BUF_X1 U386 ( .A(n719), .Z(n392) );
  BUF_X1 U387 ( .A(G143), .Z(n396) );
  NOR2_X2 U388 ( .A1(n671), .A2(n433), .ZN(n435) );
  NAND2_X2 U389 ( .A1(n753), .A2(n758), .ZN(n565) );
  XNOR2_X2 U390 ( .A(n564), .B(KEYINPUT111), .ZN(n753) );
  NOR2_X2 U391 ( .A1(n385), .A2(n382), .ZN(n649) );
  XNOR2_X2 U392 ( .A(G125), .B(G146), .ZN(n488) );
  XNOR2_X2 U393 ( .A(n522), .B(G469), .ZN(n562) );
  XNOR2_X1 U394 ( .A(n398), .B(n477), .ZN(n479) );
  XNOR2_X1 U395 ( .A(n461), .B(G902), .ZN(n665) );
  XNOR2_X1 U396 ( .A(G119), .B(G101), .ZN(n417) );
  NOR2_X1 U397 ( .A1(n673), .A2(n672), .ZN(n736) );
  BUF_X1 U398 ( .A(n621), .Z(n732) );
  NOR2_X1 U399 ( .A1(n596), .A2(n595), .ZN(n607) );
  XNOR2_X1 U400 ( .A(n380), .B(n577), .ZN(n605) );
  NAND2_X1 U401 ( .A1(n374), .A2(n372), .ZN(n380) );
  XNOR2_X1 U402 ( .A(n369), .B(n357), .ZN(n788) );
  NAND2_X1 U403 ( .A1(n668), .A2(n665), .ZN(n433) );
  NAND2_X1 U404 ( .A1(n387), .A2(n389), .ZN(n386) );
  AND2_X1 U405 ( .A1(n587), .A2(n574), .ZN(n379) );
  NOR2_X1 U406 ( .A1(KEYINPUT47), .A2(n626), .ZN(n627) );
  XNOR2_X1 U407 ( .A(n506), .B(n505), .ZN(n590) );
  NOR2_X1 U408 ( .A1(n453), .A2(n452), .ZN(n420) );
  XNOR2_X1 U409 ( .A(n630), .B(KEYINPUT30), .ZN(n452) );
  XNOR2_X1 U410 ( .A(n468), .B(n467), .ZN(n622) );
  XNOR2_X1 U411 ( .A(n682), .B(n681), .ZN(n683) );
  OR2_X1 U412 ( .A1(n700), .A2(n665), .ZN(n465) );
  NAND2_X1 U413 ( .A1(n680), .A2(n548), .ZN(n550) );
  XNOR2_X1 U414 ( .A(n447), .B(n542), .ZN(n545) );
  XNOR2_X1 U415 ( .A(n479), .B(n478), .ZN(n421) );
  XNOR2_X1 U416 ( .A(n416), .B(G104), .ZN(n492) );
  XNOR2_X1 U417 ( .A(n417), .B(KEYINPUT3), .ZN(n543) );
  XNOR2_X1 U418 ( .A(G122), .B(G113), .ZN(n416) );
  XNOR2_X1 U419 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n413) );
  INV_X1 U420 ( .A(KEYINPUT81), .ZN(n389) );
  XOR2_X1 U421 ( .A(KEYINPUT87), .B(KEYINPUT46), .Z(n653) );
  XNOR2_X2 U422 ( .A(n508), .B(n507), .ZN(n779) );
  XNOR2_X1 U423 ( .A(G131), .B(G134), .ZN(n507) );
  OR2_X1 U424 ( .A1(n739), .A2(n738), .ZN(n583) );
  XNOR2_X1 U425 ( .A(n411), .B(G116), .ZN(n482) );
  INV_X1 U426 ( .A(G107), .ZN(n411) );
  NAND2_X1 U427 ( .A1(n790), .A2(n384), .ZN(n383) );
  AND2_X1 U428 ( .A1(n636), .A2(KEYINPUT81), .ZN(n384) );
  NOR2_X1 U429 ( .A1(n788), .A2(n652), .ZN(n654) );
  INV_X1 U430 ( .A(KEYINPUT15), .ZN(n461) );
  XNOR2_X1 U431 ( .A(G110), .B(G101), .ZN(n511) );
  INV_X1 U432 ( .A(G140), .ZN(n510) );
  AND2_X1 U433 ( .A1(n376), .A2(n576), .ZN(n375) );
  NAND2_X1 U434 ( .A1(n769), .A2(n379), .ZN(n378) );
  NOR2_X1 U435 ( .A1(n622), .A2(n473), .ZN(n418) );
  INV_X1 U436 ( .A(G902), .ZN(n548) );
  XNOR2_X1 U437 ( .A(n496), .B(n495), .ZN(n688) );
  INV_X1 U438 ( .A(G146), .ZN(n509) );
  XOR2_X1 U439 ( .A(G107), .B(KEYINPUT76), .Z(n518) );
  INV_X1 U440 ( .A(n736), .ZN(n448) );
  XNOR2_X1 U441 ( .A(n371), .B(n370), .ZN(n664) );
  INV_X1 U442 ( .A(KEYINPUT39), .ZN(n370) );
  NOR2_X1 U443 ( .A1(n453), .A2(n394), .ZN(n393) );
  OR2_X1 U444 ( .A1(n582), .A2(n581), .ZN(n663) );
  INV_X1 U445 ( .A(n583), .ZN(n742) );
  XNOR2_X1 U446 ( .A(n535), .B(n359), .ZN(n395) );
  NOR2_X1 U447 ( .A1(n674), .A2(G902), .ZN(n422) );
  BUF_X1 U448 ( .A(n446), .Z(n780) );
  XNOR2_X1 U449 ( .A(n412), .B(n482), .ZN(n410) );
  XNOR2_X1 U450 ( .A(n543), .B(n492), .ZN(n415) );
  XNOR2_X1 U451 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U452 ( .A(n427), .B(n425), .ZN(n774) );
  XNOR2_X1 U453 ( .A(n426), .B(n483), .ZN(n425) );
  AND2_X1 U454 ( .A1(n677), .A2(G953), .ZN(n777) );
  INV_X1 U455 ( .A(n636), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n424), .B(n423), .ZN(n754) );
  INV_X1 U457 ( .A(KEYINPUT103), .ZN(n423) );
  NAND2_X1 U458 ( .A1(n356), .A2(n663), .ZN(n424) );
  NAND2_X1 U459 ( .A1(n404), .A2(n358), .ZN(n408) );
  NOR2_X1 U460 ( .A1(n603), .A2(KEYINPUT65), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n632), .B(n563), .ZN(n755) );
  INV_X1 U462 ( .A(G234), .ZN(n499) );
  INV_X1 U463 ( .A(G116), .ZN(n539) );
  XNOR2_X1 U464 ( .A(G137), .B(G113), .ZN(n540) );
  XOR2_X1 U465 ( .A(KEYINPUT100), .B(G131), .Z(n491) );
  XNOR2_X1 U466 ( .A(G140), .B(n396), .ZN(n490) );
  XNOR2_X1 U467 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n454) );
  XNOR2_X1 U468 ( .A(n441), .B(n362), .ZN(n471) );
  XNOR2_X1 U469 ( .A(KEYINPUT73), .B(KEYINPUT14), .ZN(n441) );
  INV_X1 U470 ( .A(n574), .ZN(n377) );
  XNOR2_X1 U471 ( .A(n573), .B(KEYINPUT74), .ZN(n381) );
  NOR2_X1 U472 ( .A1(n572), .A2(n583), .ZN(n573) );
  XNOR2_X1 U473 ( .A(n562), .B(n401), .ZN(n572) );
  INV_X1 U474 ( .A(KEYINPUT1), .ZN(n401) );
  XNOR2_X1 U475 ( .A(G110), .B(KEYINPUT16), .ZN(n414) );
  XNOR2_X1 U476 ( .A(G122), .B(G134), .ZN(n475) );
  XNOR2_X1 U477 ( .A(n481), .B(n482), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n440), .B(n439), .ZN(n767) );
  INV_X1 U479 ( .A(KEYINPUT91), .ZN(n439) );
  NAND2_X1 U480 ( .A1(n471), .A2(G952), .ZN(n440) );
  BUF_X1 U481 ( .A(n632), .Z(n659) );
  NOR2_X1 U482 ( .A1(n356), .A2(n639), .ZN(n641) );
  AND2_X1 U483 ( .A1(n381), .A2(n584), .ZN(n748) );
  XNOR2_X1 U484 ( .A(n498), .B(n497), .ZN(n581) );
  XNOR2_X1 U485 ( .A(n484), .B(G478), .ZN(n582) );
  XNOR2_X1 U486 ( .A(n533), .B(n778), .ZN(n674) );
  XNOR2_X1 U487 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U488 ( .A(n544), .B(n521), .ZN(n695) );
  XNOR2_X1 U489 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U490 ( .A(n700), .B(n701), .ZN(n702) );
  XNOR2_X1 U491 ( .A(n568), .B(n567), .ZN(n652) );
  NOR2_X1 U492 ( .A1(n664), .A2(n356), .ZN(n369) );
  NAND2_X1 U493 ( .A1(n742), .A2(n562), .ZN(n631) );
  XNOR2_X1 U494 ( .A(n776), .B(n775), .ZN(n402) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(G75) );
  XNOR2_X1 U496 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n443) );
  OR2_X1 U497 ( .A1(n772), .A2(n445), .ZN(n444) );
  NAND2_X1 U498 ( .A1(n361), .A2(n446), .ZN(n445) );
  XOR2_X1 U499 ( .A(n651), .B(KEYINPUT40), .Z(n357) );
  AND2_X1 U500 ( .A1(n403), .A2(n400), .ZN(n358) );
  XOR2_X1 U501 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n359) );
  XOR2_X1 U502 ( .A(G104), .B(KEYINPUT75), .Z(n360) );
  NAND2_X1 U503 ( .A1(n432), .A2(n668), .ZN(n733) );
  INV_X2 U504 ( .A(G953), .ZN(n446) );
  INV_X1 U505 ( .A(n504), .ZN(n587) );
  XNOR2_X1 U506 ( .A(n418), .B(n474), .ZN(n504) );
  NOR2_X1 U507 ( .A1(n771), .A2(n770), .ZN(n361) );
  OR2_X1 U508 ( .A1(n558), .A2(n557), .ZN(n638) );
  AND2_X1 U509 ( .A1(G237), .A2(G234), .ZN(n362) );
  AND2_X1 U510 ( .A1(n562), .A2(n638), .ZN(n363) );
  INV_X1 U511 ( .A(n755), .ZN(n394) );
  XNOR2_X1 U512 ( .A(n415), .B(n410), .ZN(n615) );
  BUF_X1 U513 ( .A(n624), .Z(n364) );
  AND2_X2 U514 ( .A1(n449), .A2(n448), .ZN(n699) );
  XNOR2_X1 U515 ( .A(n450), .B(KEYINPUT64), .ZN(n449) );
  NAND2_X1 U516 ( .A1(n365), .A2(n787), .ZN(n662) );
  XNOR2_X1 U517 ( .A(n366), .B(n655), .ZN(n365) );
  NAND2_X1 U518 ( .A1(n368), .A2(n367), .ZN(n366) );
  XNOR2_X1 U519 ( .A(n654), .B(n653), .ZN(n367) );
  XNOR2_X1 U520 ( .A(n650), .B(KEYINPUT69), .ZN(n368) );
  NAND2_X1 U521 ( .A1(n393), .A2(n419), .ZN(n371) );
  NAND2_X1 U522 ( .A1(n373), .A2(n377), .ZN(n372) );
  INV_X1 U523 ( .A(n769), .ZN(n373) );
  AND2_X1 U524 ( .A1(n378), .A2(n375), .ZN(n374) );
  NAND2_X1 U525 ( .A1(n504), .A2(n377), .ZN(n376) );
  NAND2_X1 U526 ( .A1(n381), .A2(n645), .ZN(n442) );
  NAND2_X1 U527 ( .A1(n388), .A2(n386), .ZN(n385) );
  NAND2_X1 U528 ( .A1(n390), .A2(n389), .ZN(n388) );
  INV_X1 U529 ( .A(n790), .ZN(n390) );
  XNOR2_X2 U530 ( .A(n635), .B(KEYINPUT108), .ZN(n790) );
  XNOR2_X1 U531 ( .A(n391), .B(n486), .ZN(n489) );
  XNOR2_X1 U532 ( .A(n487), .B(n485), .ZN(n391) );
  AND2_X1 U533 ( .A1(n430), .A2(n428), .ZN(n397) );
  XNOR2_X1 U534 ( .A(n530), .B(n529), .ZN(n533) );
  XNOR2_X1 U535 ( .A(n438), .B(n561), .ZN(n437) );
  XNOR2_X2 U536 ( .A(n422), .B(n395), .ZN(n739) );
  NAND2_X1 U537 ( .A1(n544), .A2(n545), .ZN(n546) );
  XNOR2_X2 U538 ( .A(n779), .B(n509), .ZN(n544) );
  XNOR2_X1 U539 ( .A(n436), .B(KEYINPUT109), .ZN(n624) );
  NAND2_X1 U540 ( .A1(n397), .A2(n649), .ZN(n650) );
  NAND2_X1 U541 ( .A1(n446), .A2(G234), .ZN(n398) );
  XNOR2_X2 U542 ( .A(n399), .B(KEYINPUT45), .ZN(n621) );
  NAND2_X1 U543 ( .A1(n606), .A2(n607), .ZN(n399) );
  NAND2_X1 U544 ( .A1(n597), .A2(n578), .ZN(n407) );
  NOR2_X1 U545 ( .A1(n402), .A2(n777), .ZN(G63) );
  NAND2_X1 U546 ( .A1(n605), .A2(n604), .ZN(n403) );
  OR2_X1 U547 ( .A1(n620), .A2(n603), .ZN(n409) );
  INV_X1 U548 ( .A(n620), .ZN(n404) );
  NAND2_X1 U549 ( .A1(n408), .A2(n405), .ZN(n606) );
  NAND2_X1 U550 ( .A1(n406), .A2(n409), .ZN(n405) );
  NAND2_X1 U551 ( .A1(n407), .A2(n598), .ZN(n406) );
  INV_X1 U552 ( .A(n452), .ZN(n419) );
  NAND2_X1 U553 ( .A1(n420), .A2(n634), .ZN(n635) );
  NAND2_X1 U554 ( .A1(n421), .A2(G221), .ZN(n530) );
  NAND2_X1 U555 ( .A1(n421), .A2(G217), .ZN(n427) );
  INV_X1 U556 ( .A(n663), .ZN(n724) );
  NAND2_X1 U557 ( .A1(n429), .A2(n392), .ZN(n428) );
  XNOR2_X1 U558 ( .A(n627), .B(KEYINPUT72), .ZN(n429) );
  XNOR2_X1 U559 ( .A(n431), .B(n625), .ZN(n430) );
  NOR2_X2 U560 ( .A1(n719), .A2(n628), .ZN(n431) );
  INV_X1 U561 ( .A(n672), .ZN(n432) );
  XNOR2_X1 U562 ( .A(n434), .B(KEYINPUT84), .ZN(n451) );
  NAND2_X1 U563 ( .A1(n435), .A2(n621), .ZN(n434) );
  NAND2_X1 U564 ( .A1(n437), .A2(n562), .ZN(n436) );
  NAND2_X1 U565 ( .A1(n560), .A2(n629), .ZN(n438) );
  XNOR2_X2 U566 ( .A(n442), .B(KEYINPUT33), .ZN(n769) );
  OR2_X2 U567 ( .A1(n544), .A2(n545), .ZN(n547) );
  XNOR2_X1 U568 ( .A(n543), .B(n541), .ZN(n447) );
  NAND2_X1 U569 ( .A1(n451), .A2(n667), .ZN(n450) );
  NAND2_X1 U570 ( .A1(n742), .A2(n363), .ZN(n453) );
  XNOR2_X1 U571 ( .A(n676), .B(n675), .ZN(n678) );
  NAND2_X1 U572 ( .A1(n678), .A2(n704), .ZN(n679) );
  INV_X1 U573 ( .A(n674), .ZN(n675) );
  BUF_X1 U574 ( .A(n699), .Z(n773) );
  NAND2_X1 U575 ( .A1(n699), .A2(G217), .ZN(n676) );
  INV_X1 U576 ( .A(KEYINPUT82), .ZN(n625) );
  XNOR2_X1 U577 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U578 ( .A1(n789), .A2(n578), .ZN(n580) );
  NAND2_X1 U579 ( .A1(n755), .A2(n756), .ZN(n564) );
  XNOR2_X1 U580 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U581 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n455) );
  XNOR2_X1 U582 ( .A(n455), .B(n454), .ZN(n458) );
  NAND2_X1 U583 ( .A1(n446), .A2(G224), .ZN(n456) );
  XNOR2_X1 U584 ( .A(n488), .B(n456), .ZN(n457) );
  XNOR2_X1 U585 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X2 U586 ( .A(G128), .B(G143), .ZN(n480) );
  XNOR2_X2 U587 ( .A(n480), .B(KEYINPUT4), .ZN(n508) );
  XNOR2_X1 U588 ( .A(n508), .B(n459), .ZN(n460) );
  XNOR2_X1 U589 ( .A(n615), .B(n460), .ZN(n700) );
  NAND2_X1 U590 ( .A1(n548), .A2(n469), .ZN(n466) );
  NAND2_X1 U591 ( .A1(n466), .A2(G210), .ZN(n463) );
  INV_X1 U592 ( .A(KEYINPUT90), .ZN(n462) );
  XNOR2_X1 U593 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X2 U594 ( .A(n465), .B(n464), .ZN(n632) );
  NAND2_X1 U595 ( .A1(n466), .A2(G214), .ZN(n756) );
  NAND2_X1 U596 ( .A1(n632), .A2(n756), .ZN(n468) );
  INV_X1 U597 ( .A(KEYINPUT19), .ZN(n467) );
  NOR2_X1 U598 ( .A1(G953), .A2(n767), .ZN(n470) );
  XNOR2_X1 U599 ( .A(n470), .B(KEYINPUT92), .ZN(n558) );
  NAND2_X1 U600 ( .A1(G902), .A2(n471), .ZN(n555) );
  XNOR2_X1 U601 ( .A(G898), .B(KEYINPUT93), .ZN(n612) );
  NAND2_X1 U602 ( .A1(G953), .A2(n612), .ZN(n616) );
  NOR2_X1 U603 ( .A1(n555), .A2(n616), .ZN(n472) );
  NOR2_X1 U604 ( .A1(n558), .A2(n472), .ZN(n473) );
  INV_X1 U605 ( .A(KEYINPUT0), .ZN(n474) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n476) );
  XNOR2_X1 U607 ( .A(n476), .B(n475), .ZN(n483) );
  INV_X1 U608 ( .A(KEYINPUT68), .ZN(n477) );
  XOR2_X1 U609 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n478) );
  BUF_X1 U610 ( .A(n480), .Z(n481) );
  NOR2_X1 U611 ( .A1(G902), .A2(n774), .ZN(n484) );
  XOR2_X1 U612 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n486) );
  XNOR2_X1 U613 ( .A(KEYINPUT101), .B(KEYINPUT12), .ZN(n485) );
  NAND2_X1 U614 ( .A1(G214), .A2(n536), .ZN(n487) );
  XNOR2_X1 U615 ( .A(n488), .B(KEYINPUT10), .ZN(n532) );
  XNOR2_X1 U616 ( .A(n489), .B(n532), .ZN(n496) );
  XNOR2_X1 U617 ( .A(n491), .B(n490), .ZN(n494) );
  INV_X1 U618 ( .A(n492), .ZN(n493) );
  XNOR2_X1 U619 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U620 ( .A1(n688), .A2(n548), .ZN(n498) );
  XOR2_X1 U621 ( .A(KEYINPUT13), .B(G475), .Z(n497) );
  INV_X1 U622 ( .A(n581), .ZN(n575) );
  AND2_X1 U623 ( .A1(n582), .A2(n575), .ZN(n758) );
  OR2_X1 U624 ( .A1(n665), .A2(n499), .ZN(n500) );
  XNOR2_X1 U625 ( .A(n500), .B(KEYINPUT20), .ZN(n534) );
  NAND2_X1 U626 ( .A1(n534), .A2(G221), .ZN(n502) );
  INV_X1 U627 ( .A(KEYINPUT21), .ZN(n501) );
  XNOR2_X1 U628 ( .A(n502), .B(n501), .ZN(n640) );
  NAND2_X1 U629 ( .A1(n758), .A2(n640), .ZN(n503) );
  OR2_X1 U630 ( .A1(n504), .A2(n503), .ZN(n506) );
  INV_X1 U631 ( .A(KEYINPUT22), .ZN(n505) );
  INV_X1 U632 ( .A(n590), .ZN(n554) );
  XNOR2_X1 U633 ( .A(n510), .B(G137), .ZN(n531) );
  XNOR2_X1 U634 ( .A(n360), .B(n511), .ZN(n513) );
  INV_X1 U635 ( .A(n513), .ZN(n512) );
  NAND2_X1 U636 ( .A1(n531), .A2(n512), .ZN(n516) );
  INV_X1 U637 ( .A(n531), .ZN(n514) );
  NAND2_X1 U638 ( .A1(n514), .A2(n513), .ZN(n515) );
  NAND2_X1 U639 ( .A1(n516), .A2(n515), .ZN(n520) );
  NAND2_X1 U640 ( .A1(G227), .A2(n780), .ZN(n517) );
  NAND2_X1 U641 ( .A1(n695), .A2(n548), .ZN(n522) );
  INV_X1 U642 ( .A(n572), .ZN(n743) );
  XNOR2_X1 U643 ( .A(G110), .B(G128), .ZN(n524) );
  XNOR2_X1 U644 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n523) );
  XNOR2_X1 U645 ( .A(n524), .B(n523), .ZN(n528) );
  XNOR2_X1 U646 ( .A(G119), .B(KEYINPUT94), .ZN(n526) );
  XNOR2_X1 U647 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n525) );
  XNOR2_X1 U648 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U649 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U650 ( .A(n532), .B(n531), .ZN(n778) );
  AND2_X1 U651 ( .A1(n534), .A2(G217), .ZN(n535) );
  INV_X1 U652 ( .A(n739), .ZN(n642) );
  NOR2_X1 U653 ( .A1(n743), .A2(n642), .ZN(n552) );
  XOR2_X1 U654 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n538) );
  NAND2_X1 U655 ( .A1(n536), .A2(G210), .ZN(n537) );
  XNOR2_X1 U656 ( .A(n538), .B(n537), .ZN(n542) );
  NAND2_X1 U657 ( .A1(n547), .A2(n546), .ZN(n680) );
  INV_X1 U658 ( .A(G472), .ZN(n549) );
  XNOR2_X2 U659 ( .A(n550), .B(n549), .ZN(n569) );
  XNOR2_X2 U660 ( .A(n569), .B(KEYINPUT105), .ZN(n629) );
  INV_X1 U661 ( .A(n629), .ZN(n551) );
  NAND2_X1 U662 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U663 ( .A1(n554), .A2(n553), .ZN(n603) );
  XOR2_X1 U664 ( .A(G110), .B(n603), .Z(G12) );
  NOR2_X1 U665 ( .A1(G900), .A2(n555), .ZN(n556) );
  AND2_X1 U666 ( .A1(G953), .A2(n556), .ZN(n557) );
  AND2_X1 U667 ( .A1(n638), .A2(n640), .ZN(n559) );
  INV_X1 U668 ( .A(KEYINPUT28), .ZN(n561) );
  INV_X1 U669 ( .A(KEYINPUT38), .ZN(n563) );
  XNOR2_X2 U670 ( .A(n565), .B(KEYINPUT41), .ZN(n768) );
  NAND2_X1 U671 ( .A1(n364), .A2(n768), .ZN(n568) );
  XNOR2_X1 U672 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n566) );
  XNOR2_X1 U673 ( .A(n566), .B(KEYINPUT112), .ZN(n567) );
  XOR2_X1 U674 ( .A(n652), .B(G137), .Z(G39) );
  BUF_X1 U675 ( .A(n569), .Z(n570) );
  INV_X1 U676 ( .A(n570), .ZN(n584) );
  INV_X1 U677 ( .A(KEYINPUT6), .ZN(n571) );
  XNOR2_X1 U678 ( .A(n570), .B(n571), .ZN(n637) );
  INV_X1 U679 ( .A(n640), .ZN(n738) );
  XNOR2_X1 U680 ( .A(KEYINPUT34), .B(KEYINPUT79), .ZN(n574) );
  OR2_X1 U681 ( .A1(n582), .A2(n575), .ZN(n633) );
  INV_X1 U682 ( .A(n633), .ZN(n576) );
  INV_X1 U683 ( .A(KEYINPUT35), .ZN(n577) );
  INV_X1 U684 ( .A(n605), .ZN(n789) );
  INV_X1 U685 ( .A(KEYINPUT44), .ZN(n578) );
  NOR2_X1 U686 ( .A1(KEYINPUT44), .A2(KEYINPUT65), .ZN(n579) );
  NOR2_X1 U687 ( .A1(n580), .A2(n579), .ZN(n596) );
  XNOR2_X1 U688 ( .A(KEYINPUT83), .B(n754), .ZN(n626) );
  NOR2_X1 U689 ( .A1(n631), .A2(n584), .ZN(n585) );
  NAND2_X1 U690 ( .A1(n587), .A2(n585), .ZN(n586) );
  XNOR2_X1 U691 ( .A(KEYINPUT99), .B(n586), .ZN(n713) );
  NAND2_X1 U692 ( .A1(n748), .A2(n587), .ZN(n588) );
  XNOR2_X1 U693 ( .A(n588), .B(KEYINPUT31), .ZN(n725) );
  NOR2_X1 U694 ( .A1(n713), .A2(n725), .ZN(n589) );
  NOR2_X1 U695 ( .A1(n626), .A2(n589), .ZN(n594) );
  NAND2_X1 U696 ( .A1(n590), .A2(n637), .ZN(n601) );
  INV_X1 U697 ( .A(KEYINPUT88), .ZN(n591) );
  XNOR2_X1 U698 ( .A(n601), .B(n591), .ZN(n593) );
  NOR2_X1 U699 ( .A1(n743), .A2(n739), .ZN(n592) );
  AND2_X1 U700 ( .A1(n593), .A2(n592), .ZN(n708) );
  OR2_X1 U701 ( .A1(n594), .A2(n708), .ZN(n595) );
  NAND2_X1 U702 ( .A1(KEYINPUT89), .A2(n605), .ZN(n597) );
  INV_X1 U703 ( .A(KEYINPUT65), .ZN(n598) );
  NAND2_X1 U704 ( .A1(n743), .A2(n739), .ZN(n599) );
  XNOR2_X1 U705 ( .A(n599), .B(KEYINPUT104), .ZN(n600) );
  NOR2_X1 U706 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U707 ( .A(n602), .B(KEYINPUT32), .ZN(n620) );
  NOR2_X1 U708 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n604) );
  NAND2_X1 U709 ( .A1(n732), .A2(n780), .ZN(n608) );
  XNOR2_X1 U710 ( .A(n608), .B(KEYINPUT127), .ZN(n614) );
  XOR2_X1 U711 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n610) );
  NAND2_X1 U712 ( .A1(G224), .A2(G953), .ZN(n609) );
  XNOR2_X1 U713 ( .A(n610), .B(n609), .ZN(n611) );
  NOR2_X1 U714 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U715 ( .A1(n614), .A2(n613), .ZN(n619) );
  INV_X1 U716 ( .A(n615), .ZN(n617) );
  NAND2_X1 U717 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U718 ( .A(n619), .B(n618), .ZN(G69) );
  XOR2_X1 U719 ( .A(G119), .B(n620), .Z(G21) );
  INV_X1 U720 ( .A(n622), .ZN(n623) );
  AND2_X2 U721 ( .A1(n624), .A2(n623), .ZN(n719) );
  INV_X1 U722 ( .A(KEYINPUT47), .ZN(n628) );
  OR2_X1 U723 ( .A1(n754), .A2(n628), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n629), .A2(n756), .ZN(n630) );
  INV_X1 U725 ( .A(n659), .ZN(n646) );
  NOR2_X1 U726 ( .A1(n646), .A2(n633), .ZN(n634) );
  INV_X1 U727 ( .A(n637), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n638), .A2(n756), .ZN(n639) );
  NAND2_X1 U729 ( .A1(n641), .A2(n640), .ZN(n643) );
  NOR2_X1 U730 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n647), .B(KEYINPUT36), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n648), .A2(n743), .ZN(n729) );
  INV_X1 U734 ( .A(KEYINPUT110), .ZN(n651) );
  INV_X1 U735 ( .A(KEYINPUT48), .ZN(n655) );
  XNOR2_X1 U736 ( .A(KEYINPUT106), .B(n656), .ZN(n657) );
  NOR2_X1 U737 ( .A1(n743), .A2(n657), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(KEYINPUT43), .ZN(n660) );
  NOR2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n661), .B(KEYINPUT107), .ZN(n787) );
  XNOR2_X1 U741 ( .A(n662), .B(KEYINPUT86), .ZN(n671) );
  OR2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n668) );
  INV_X1 U743 ( .A(n668), .ZN(n730) );
  XOR2_X1 U744 ( .A(KEYINPUT85), .B(n665), .Z(n666) );
  NAND2_X1 U745 ( .A1(n666), .A2(KEYINPUT2), .ZN(n667) );
  NAND2_X1 U746 ( .A1(KEYINPUT2), .A2(n668), .ZN(n669) );
  XOR2_X1 U747 ( .A(KEYINPUT80), .B(n669), .Z(n670) );
  NAND2_X1 U748 ( .A1(n732), .A2(n670), .ZN(n673) );
  BUF_X1 U749 ( .A(n671), .Z(n672) );
  INV_X1 U750 ( .A(G952), .ZN(n677) );
  INV_X1 U751 ( .A(n777), .ZN(n704) );
  XNOR2_X1 U752 ( .A(n679), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U753 ( .A1(n699), .A2(G472), .ZN(n684) );
  BUF_X1 U754 ( .A(n680), .Z(n682) );
  XNOR2_X1 U755 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n681) );
  XNOR2_X1 U756 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n685), .A2(n704), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n686), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U759 ( .A1(n699), .A2(G475), .ZN(n690) );
  XOR2_X1 U760 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n687) );
  XNOR2_X1 U761 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n691), .A2(n704), .ZN(n693) );
  INV_X1 U763 ( .A(KEYINPUT60), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n693), .B(n692), .ZN(G60) );
  NAND2_X1 U765 ( .A1(n773), .A2(G469), .ZN(n697) );
  XNOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n694) );
  XNOR2_X1 U767 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U768 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U769 ( .A1(n698), .A2(n777), .ZN(G54) );
  NAND2_X1 U770 ( .A1(n699), .A2(G210), .ZN(n703) );
  XNOR2_X1 U771 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n701) );
  XNOR2_X1 U772 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n707) );
  INV_X1 U774 ( .A(KEYINPUT56), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n707), .B(n706), .ZN(G51) );
  XOR2_X1 U776 ( .A(G101), .B(n708), .Z(G3) );
  NAND2_X1 U777 ( .A1(n713), .A2(n721), .ZN(n709) );
  XNOR2_X1 U778 ( .A(n709), .B(G104), .ZN(G6) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n711) );
  XNOR2_X1 U780 ( .A(G107), .B(KEYINPUT26), .ZN(n710) );
  XNOR2_X1 U781 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U782 ( .A(KEYINPUT115), .B(n712), .Z(n715) );
  NAND2_X1 U783 ( .A1(n713), .A2(n724), .ZN(n714) );
  XNOR2_X1 U784 ( .A(n715), .B(n714), .ZN(G9) );
  XOR2_X1 U785 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n717) );
  NAND2_X1 U786 ( .A1(n392), .A2(n724), .ZN(n716) );
  XNOR2_X1 U787 ( .A(n717), .B(n716), .ZN(n718) );
  XOR2_X1 U788 ( .A(G128), .B(n718), .Z(G30) );
  NAND2_X1 U789 ( .A1(n392), .A2(n721), .ZN(n720) );
  XNOR2_X1 U790 ( .A(n720), .B(G146), .ZN(G48) );
  NAND2_X1 U791 ( .A1(n725), .A2(n721), .ZN(n722) );
  XNOR2_X1 U792 ( .A(n722), .B(KEYINPUT118), .ZN(n723) );
  XNOR2_X1 U793 ( .A(G113), .B(n723), .ZN(G15) );
  XOR2_X1 U794 ( .A(G116), .B(KEYINPUT119), .Z(n727) );
  NAND2_X1 U795 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U796 ( .A(n727), .B(n726), .ZN(G18) );
  XOR2_X1 U797 ( .A(G125), .B(KEYINPUT37), .Z(n728) );
  XNOR2_X1 U798 ( .A(n729), .B(n728), .ZN(G27) );
  XNOR2_X1 U799 ( .A(G134), .B(KEYINPUT120), .ZN(n731) );
  XOR2_X1 U800 ( .A(n731), .B(n730), .Z(G36) );
  INV_X1 U801 ( .A(n732), .ZN(n734) );
  NOR2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U803 ( .A1(n735), .A2(KEYINPUT2), .ZN(n737) );
  NOR2_X1 U804 ( .A1(n737), .A2(n736), .ZN(n772) );
  NAND2_X1 U805 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U806 ( .A(KEYINPUT49), .B(n740), .Z(n741) );
  NAND2_X1 U807 ( .A1(n570), .A2(n741), .ZN(n746) );
  NOR2_X1 U808 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U809 ( .A(n744), .B(KEYINPUT50), .ZN(n745) );
  NOR2_X1 U810 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U811 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U812 ( .A(KEYINPUT121), .B(n749), .Z(n750) );
  XNOR2_X1 U813 ( .A(KEYINPUT51), .B(n750), .ZN(n751) );
  NAND2_X1 U814 ( .A1(n751), .A2(n768), .ZN(n752) );
  XNOR2_X1 U815 ( .A(n752), .B(KEYINPUT122), .ZN(n764) );
  NAND2_X1 U816 ( .A1(n754), .A2(n753), .ZN(n761) );
  INV_X1 U817 ( .A(n756), .ZN(n757) );
  NAND2_X1 U818 ( .A1(n394), .A2(n757), .ZN(n759) );
  NAND2_X1 U819 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U820 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U821 ( .A1(n769), .A2(n762), .ZN(n763) );
  NAND2_X1 U822 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U823 ( .A(KEYINPUT52), .B(n765), .Z(n766) );
  NOR2_X1 U824 ( .A1(n767), .A2(n766), .ZN(n771) );
  AND2_X1 U825 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U826 ( .A1(n773), .A2(G478), .ZN(n776) );
  XNOR2_X1 U827 ( .A(n774), .B(KEYINPUT124), .ZN(n775) );
  XNOR2_X1 U828 ( .A(n779), .B(n778), .ZN(n782) );
  XNOR2_X1 U829 ( .A(n733), .B(n782), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n781), .A2(n780), .ZN(n786) );
  XNOR2_X1 U831 ( .A(n782), .B(G227), .ZN(n783) );
  NAND2_X1 U832 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U833 ( .A1(n784), .A2(G953), .ZN(n785) );
  NAND2_X1 U834 ( .A1(n786), .A2(n785), .ZN(G72) );
  XNOR2_X1 U835 ( .A(G140), .B(n787), .ZN(G42) );
  XOR2_X1 U836 ( .A(n788), .B(G131), .Z(G33) );
  XOR2_X1 U837 ( .A(G122), .B(n789), .Z(G24) );
  XNOR2_X1 U838 ( .A(n790), .B(n396), .ZN(G45) );
endmodule

