//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n459), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n465), .A2(new_n459), .ZN(new_n476));
  AOI22_X1  g051(.A1(G124), .A2(new_n476), .B1(new_n466), .B2(G136), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT66), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(KEYINPUT66), .A2(G100), .A3(G2105), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G112), .B2(new_n459), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n477), .A2(new_n481), .ZN(G162));
  NAND2_X1  g057(.A1(new_n470), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G126), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n459), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n467), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n466), .A2(new_n490), .A3(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G651), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT67), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(new_n493), .A3(G651), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(KEYINPUT68), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n499), .A2(new_n506), .A3(KEYINPUT69), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT69), .B1(new_n499), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n500), .A2(KEYINPUT68), .A3(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT68), .B1(new_n500), .B2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(G50), .A2(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n518), .A2(G651), .B1(new_n499), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  INV_X1    g097(.A(G63), .ZN(new_n523));
  NAND2_X1  g098(.A1(G76), .A2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n516), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(G651), .B1(new_n527), .B2(new_n525), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  INV_X1    g104(.A(new_n494), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n497), .B1(new_n493), .B2(G651), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n495), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n535), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(G543), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n528), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n533), .B2(new_n516), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n499), .A2(new_n506), .A3(KEYINPUT69), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT73), .B(G89), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n538), .A2(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n516), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n537), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT74), .B(G90), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n540), .A2(new_n541), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(G171));
  INV_X1    g130(.A(new_n537), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G43), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT75), .B(G81), .Z(new_n558));
  NAND2_X1  g133(.A1(new_n509), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n516), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g143(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n569));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND4_X1  g147(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n536), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n503), .B1(new_n533), .B2(KEYINPUT71), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n576), .A2(KEYINPUT78), .A3(G53), .A4(new_n536), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n573), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT79), .B1(new_n507), .B2(new_n508), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n540), .A2(new_n582), .A3(new_n541), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n583), .A3(G91), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n495), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n578), .A2(new_n580), .A3(new_n584), .A4(new_n586), .ZN(G299));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n552), .B2(new_n554), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g165(.A1(new_n552), .A2(new_n554), .A3(new_n588), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(G301));
  OAI221_X1 g167(.A(new_n528), .B1(new_n529), .B2(new_n537), .C1(new_n542), .C2(new_n544), .ZN(G286));
  AND2_X1   g168(.A1(new_n581), .A2(new_n583), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G87), .ZN(new_n595));
  INV_X1    g170(.A(G74), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n495), .B1(new_n516), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n556), .B2(G49), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(KEYINPUT81), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(KEYINPUT81), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(G288));
  NAND2_X1  g177(.A1(new_n594), .A2(G86), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n499), .A2(G48), .A3(G543), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n495), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n556), .A2(G47), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n509), .A2(G85), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n609), .B(new_n610), .C1(new_n495), .C2(new_n611), .ZN(G290));
  NAND3_X1  g187(.A1(new_n581), .A2(new_n583), .A3(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT10), .A4(G92), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n495), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n516), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(KEYINPUT82), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G54), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n537), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n617), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  MUX2_X1   g205(.A(G301), .B(new_n629), .S(new_n630), .Z(G284));
  MUX2_X1   g206(.A(G301), .B(new_n629), .S(new_n630), .Z(G321));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  INV_X1    g208(.A(G299), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G868), .ZN(G297));
  OAI21_X1  g210(.A(new_n633), .B1(new_n634), .B2(G868), .ZN(G280));
  AOI21_X1  g211(.A(new_n627), .B1(new_n615), .B2(new_n616), .ZN(new_n637));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G860), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT83), .ZN(G148));
  NOR2_X1   g215(.A1(new_n565), .A2(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n638), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G868), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT84), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n470), .A2(new_n461), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  INV_X1    g223(.A(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n466), .A2(G135), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n476), .A2(G123), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n459), .A2(G111), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2096), .Z(new_n657));
  OAI211_X1 g232(.A(new_n651), .B(new_n657), .C1(new_n649), .C2(new_n648), .ZN(G156));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n664), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n678), .B2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n649), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(KEYINPUT17), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n676), .A2(new_n677), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2096), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n681), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT87), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT20), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n690), .A2(new_n691), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(new_n693), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n697), .B(new_n699), .C1(new_n689), .C2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT88), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1981), .B(G1986), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G229));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G6), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G305), .B2(G16), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n712), .A2(G23), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n599), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n711), .A2(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n716), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n714), .A2(new_n711), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n712), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n712), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1971), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(G119), .A2(new_n476), .B1(new_n466), .B2(G131), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n731));
  OAI221_X1 g306(.A(G2104), .B1(G107), .B2(new_n459), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G25), .B(new_n735), .S(G29), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT91), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n736), .B(new_n738), .Z(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G24), .ZN(new_n740));
  XNOR2_X1  g315(.A(G290), .B(KEYINPUT92), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G16), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G1986), .Z(new_n743));
  NAND4_X1  g318(.A1(new_n726), .A2(new_n727), .A3(new_n739), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT36), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G26), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n466), .A2(G140), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n476), .A2(G128), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n459), .A2(G116), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT95), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT101), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n746), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n746), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G2090), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n757), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n758), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n712), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n712), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1961), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n712), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n712), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G1966), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT100), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n764), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT26), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G129), .B2(new_n476), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n466), .A2(G141), .B1(G105), .B2(new_n461), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G29), .B2(G32), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G2090), .B2(new_n761), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n565), .A2(G16), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G16), .B2(G19), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT94), .B(G1341), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT30), .B(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n746), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT24), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n746), .B1(new_n793), .B2(G34), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n793), .B2(G34), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G160), .B2(G29), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n792), .B1(new_n746), .B2(new_n656), .C1(new_n796), .C2(G2084), .ZN(new_n797));
  NOR2_X1   g372(.A1(G27), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(G29), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(G2078), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(G2078), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n797), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n783), .A2(new_n787), .A3(new_n788), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n769), .A2(G1966), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT99), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n780), .A2(new_n781), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT97), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n746), .A2(G33), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT25), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n470), .A2(G127), .ZN(new_n811));
  NAND2_X1  g386(.A1(G115), .A2(G2104), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n459), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n810), .B(new_n813), .C1(G139), .C2(new_n466), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n746), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2072), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(G2072), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n796), .A2(G2084), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n807), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n805), .B1(new_n819), .B2(KEYINPUT98), .ZN(new_n820));
  AOI211_X1 g395(.A(new_n803), .B(new_n820), .C1(KEYINPUT98), .C2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n712), .A2(G20), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT23), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n634), .B2(new_n712), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1956), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n712), .A2(G4), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n637), .B2(new_n712), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT93), .B(G1348), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n745), .A2(new_n772), .A3(new_n821), .A4(new_n831), .ZN(G150));
  INV_X1    g407(.A(G150), .ZN(G311));
  NAND2_X1  g408(.A1(new_n637), .A2(G559), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT38), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n556), .A2(G55), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n509), .A2(G93), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n516), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G651), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n564), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n556), .A2(G43), .B1(G651), .B2(new_n562), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n509), .A2(G93), .B1(G651), .B2(new_n840), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n559), .A4(new_n836), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n835), .B(new_n847), .Z(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  AOI21_X1  g424(.A(G860), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n842), .A2(G860), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT102), .Z(G145));
  NOR2_X1   g430(.A1(new_n814), .A2(new_n777), .ZN(new_n856));
  INV_X1    g431(.A(new_n778), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(new_n814), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n735), .B(new_n647), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(G118), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(G2105), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n476), .A2(G130), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT105), .ZN(new_n864));
  AOI211_X1 g439(.A(new_n862), .B(new_n864), .C1(G142), .C2(new_n466), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n859), .A2(new_n865), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n754), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n754), .A3(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(G164), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  INV_X1    g447(.A(G164), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n872), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n858), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n872), .B2(new_n868), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(G164), .A3(new_n870), .ZN(new_n877));
  INV_X1    g452(.A(new_n858), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G162), .B(new_n656), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n882), .B(new_n883), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n875), .A2(new_n884), .A3(new_n879), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g465(.A(new_n642), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n847), .A2(KEYINPUT106), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n843), .A2(new_n846), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n843), .A2(new_n846), .A3(new_n893), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n893), .B1(new_n843), .B2(new_n846), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n642), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n617), .A2(G299), .A3(new_n628), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n637), .A2(KEYINPUT107), .A3(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n629), .A2(new_n634), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT108), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n637), .A2(G299), .ZN(new_n908));
  AOI211_X1 g483(.A(new_n907), .B(new_n908), .C1(new_n902), .C2(new_n903), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n899), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n899), .B(new_n912), .C1(new_n906), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n629), .B2(new_n634), .ZN(new_n916));
  AND4_X1   g491(.A1(KEYINPUT107), .A2(new_n617), .A3(G299), .A4(new_n628), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT107), .B1(new_n637), .B2(G299), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT110), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n905), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n915), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n904), .A2(new_n923), .A3(new_n916), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n899), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(KEYINPUT111), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND4_X1   g505(.A1(KEYINPUT112), .A2(new_n914), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT112), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n927), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n911), .A2(new_n913), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n599), .B(G305), .ZN(new_n936));
  XNOR2_X1  g511(.A(G290), .B(G303), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n936), .B(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT42), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n931), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n933), .A2(new_n934), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n941), .A2(KEYINPUT112), .A3(new_n939), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n842), .A2(new_n630), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(G331));
  NAND2_X1  g521(.A1(G171), .A2(KEYINPUT80), .ZN(new_n947));
  AOI21_X1  g522(.A(G286), .B1(new_n947), .B2(new_n589), .ZN(new_n948));
  NOR2_X1   g523(.A1(G168), .A2(G171), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n843), .B(new_n846), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(G286), .B1(new_n554), .B2(new_n552), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n847), .B(new_n951), .C1(G301), .C2(G286), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n921), .A2(new_n907), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n904), .A2(KEYINPUT108), .A3(new_n905), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n938), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n953), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n906), .B2(new_n909), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT113), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n922), .B2(new_n919), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n925), .A2(new_n953), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n921), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n938), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n888), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT115), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n963), .A2(new_n969), .A3(new_n888), .A4(new_n966), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n966), .A2(new_n888), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n938), .B1(new_n964), .B2(new_n965), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n973), .B2(new_n974), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n963), .A2(new_n976), .A3(new_n888), .A4(new_n966), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT114), .B1(new_n981), .B2(new_n972), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n983), .B(KEYINPUT44), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n978), .B1(new_n982), .B2(new_n984), .ZN(G397));
  XNOR2_X1  g560(.A(new_n754), .B(new_n756), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n777), .A2(G1996), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n986), .B(new_n987), .C1(G1996), .C2(new_n857), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(G164), .B2(G1384), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT116), .B(G40), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n990), .A2(new_n474), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT117), .ZN(new_n994));
  INV_X1    g569(.A(new_n992), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n735), .B(new_n738), .Z(new_n996));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n997), .B2(new_n996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(G290), .B(G1986), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n992), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n474), .A2(new_n991), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G164), .A2(G1384), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1976), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(new_n1008), .B2(new_n599), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n600), .A2(new_n1008), .A3(new_n601), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1012), .A2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1013), .B2(new_n1009), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n540), .A2(G86), .A3(new_n541), .ZN(new_n1015));
  OAI21_X1  g590(.A(G1981), .B1(new_n1015), .B2(new_n606), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1016), .A2(KEYINPUT119), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(KEYINPUT119), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1017), .B(new_n1018), .C1(G305), .C2(G1981), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1007), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1014), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT55), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1003), .B1(new_n1004), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1004), .A2(new_n1027), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT121), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1028), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G2090), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1004), .A2(KEYINPUT45), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1003), .A3(new_n990), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1034), .A2(new_n1035), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1026), .B1(new_n1039), .B2(new_n1006), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1036), .ZN(new_n1041));
  OR2_X1    g616(.A1(G164), .A2(G1384), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n1003), .A3(new_n1029), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n1044), .B2(G2090), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1040), .B1(new_n1026), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1024), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1966), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1038), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G2084), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1043), .A2(new_n1051), .A3(new_n1003), .A4(new_n1029), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1006), .B1(new_n1053), .B2(G168), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G286), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT123), .B1(new_n1053), .B2(new_n1006), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT51), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1006), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT51), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1054), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1066), .A2(G2078), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1038), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1038), .B2(G2078), .ZN(new_n1069));
  INV_X1    g644(.A(G1961), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1044), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G301), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1063), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1054), .A2(new_n1063), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1048), .A2(new_n1065), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1078), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1085), .A2(new_n1024), .A3(new_n1047), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(KEYINPUT126), .A3(new_n1065), .A4(new_n1081), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1046), .A2(new_n1026), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1061), .A2(G168), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(KEYINPUT63), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1040), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G305), .A2(G1981), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G288), .A2(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n1023), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1007), .B(KEYINPUT120), .Z(new_n1095));
  OAI22_X1  g670(.A1(new_n1091), .A2(new_n1024), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1089), .B1(new_n1026), .B2(new_n1046), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1014), .A2(new_n1097), .A3(new_n1023), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1096), .B1(KEYINPUT63), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1084), .A2(new_n1087), .A3(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT56), .B(G2072), .Z(new_n1101));
  OAI22_X1  g676(.A1(new_n1034), .A2(G1956), .B1(new_n1038), .B2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(G299), .B(KEYINPUT57), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1044), .A2(new_n828), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1005), .A2(new_n756), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n637), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1038), .A2(G1996), .B1(new_n1005), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n565), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n637), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1107), .B(new_n629), .ZN(new_n1118));
  OAI221_X1 g693(.A(new_n1115), .B1(new_n1107), .B2(new_n1117), .C1(new_n1118), .C2(new_n1116), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT61), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1104), .A2(KEYINPUT61), .A3(new_n1109), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1110), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  INV_X1    g699(.A(G40), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n474), .A2(new_n1125), .A3(new_n1067), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1037), .A2(new_n990), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1071), .A2(new_n1069), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1124), .B1(new_n1128), .B2(G171), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1128), .A2(new_n1073), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1124), .B1(new_n1078), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1132), .A2(new_n1134), .A3(new_n1048), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1123), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1002), .B1(new_n1100), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n735), .A2(new_n738), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n994), .A2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n754), .A2(G2067), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n995), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(G1996), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n992), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT127), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n986), .A2(new_n776), .A3(new_n775), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1148), .A2(new_n992), .B1(new_n1145), .B2(new_n1144), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT47), .Z(new_n1151));
  INV_X1    g726(.A(new_n1000), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n995), .A2(G1986), .A3(G290), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT48), .Z(new_n1154));
  AOI211_X1 g729(.A(new_n1142), .B(new_n1151), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1138), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g731(.A1(G227), .A2(new_n457), .ZN(new_n1158));
  NOR3_X1   g732(.A1(G229), .A2(G401), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n1159), .A2(new_n889), .A3(new_n981), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


