//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT33), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n210));
  OAI211_X1 g009(.A(KEYINPUT28), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT28), .A4(new_n208), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G183gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT27), .ZN(new_n220));
  INV_X1    g019(.A(new_n210), .ZN(new_n221));
  AOI21_X1  g020(.A(G190gat), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n212), .B(new_n215), .C1(new_n222), .C2(KEYINPUT28), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  INV_X1    g028(.A(G169gat), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n225), .A2(new_n226), .A3(new_n228), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT67), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n237), .A3(new_n234), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT69), .B(G113gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G120gat), .ZN(new_n241));
  INV_X1    g040(.A(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G113gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT1), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n247));
  NOR2_X1   g046(.A1(G127gat), .A2(G134gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT68), .B(G127gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n249), .B2(G134gat), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n244), .A2(new_n245), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(new_n230), .A3(new_n231), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n253), .A2(new_n254), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT24), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n234), .B(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT64), .B(G183gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(G190gat), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT25), .B(new_n255), .C1(new_n263), .C2(new_n257), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n239), .A2(new_n251), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n239), .A2(new_n265), .ZN(new_n269));
  INV_X1    g068(.A(new_n251), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n239), .A2(KEYINPUT70), .A3(new_n251), .A4(new_n265), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n273), .A2(KEYINPUT71), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT71), .B1(new_n273), .B2(new_n274), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT32), .B(new_n207), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT33), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT32), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n274), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(KEYINPUT71), .A3(new_n274), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n285));
  INV_X1    g084(.A(new_n206), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n275), .A2(new_n276), .B1(KEYINPUT32), .B2(new_n278), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT74), .B1(new_n288), .B2(new_n206), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n277), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n273), .A2(new_n274), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT34), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT31), .B(G50gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT84), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(G78gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(G106gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G228gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n302));
  INV_X1    g101(.A(G141gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(G148gat), .ZN(new_n305));
  INV_X1    g104(.A(G148gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  OR2_X1    g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(KEYINPUT2), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT82), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n306), .A2(G141gat), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n305), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n309), .B(new_n310), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n316), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G211gat), .B(G218gat), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT75), .ZN(new_n329));
  XNOR2_X1  g128(.A(G197gat), .B(G204gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(G211gat), .A2(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT22), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n329), .B(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n323), .A2(KEYINPUT86), .A3(new_n324), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n315), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n314), .B1(new_n308), .B2(new_n311), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n320), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n335), .A2(KEYINPUT29), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(KEYINPUT3), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n301), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G22gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n334), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT29), .B1(new_n346), .B2(new_n328), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n328), .B2(new_n346), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n322), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n340), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT85), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n335), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(KEYINPUT85), .A3(new_n340), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n301), .A4(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n344), .A2(new_n345), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(G22gat), .B1(new_n357), .B2(new_n343), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n300), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n298), .A2(new_n299), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT88), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT88), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n298), .A2(new_n299), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n359), .B(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n288), .A2(KEYINPUT74), .A3(new_n206), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n293), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n277), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n294), .A2(new_n366), .A3(KEYINPUT35), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n251), .A2(new_n316), .A3(new_n320), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n251), .B1(new_n340), .B2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n323), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n376), .B(new_n378), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n270), .A2(new_n340), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n373), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n385), .B2(new_n375), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n379), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n388), .A2(new_n380), .B1(new_n323), .B2(new_n377), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  NOR2_X1   g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT6), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  INV_X1    g199(.A(new_n397), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n392), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n399), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n335), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n239), .A2(new_n405), .A3(new_n265), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n239), .B2(new_n265), .ZN(new_n407));
  INV_X1    g206(.A(G226gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(KEYINPUT29), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n269), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n404), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n406), .B2(new_n407), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n239), .A2(new_n410), .A3(new_n265), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n419), .A2(new_n335), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n269), .A2(KEYINPUT76), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n239), .A2(new_n405), .A3(new_n265), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n410), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n414), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(KEYINPUT77), .A3(new_n404), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n418), .A2(new_n422), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(G36gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT78), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G8gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n418), .A2(new_n422), .A3(new_n427), .A4(new_n432), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT77), .B1(new_n426), .B2(new_n404), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n417), .B(new_n335), .C1(new_n425), .C2(new_n414), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n443), .A2(KEYINPUT79), .A3(new_n422), .A4(new_n432), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n444), .A3(new_n435), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n403), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n372), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n440), .A2(new_n444), .A3(new_n435), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n437), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n438), .A2(KEYINPUT89), .A3(new_n445), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n370), .B1(new_n369), .B2(new_n277), .ZN(new_n453));
  INV_X1    g252(.A(new_n277), .ZN(new_n454));
  AOI211_X1 g253(.A(new_n293), .B(new_n454), .C1(new_n367), .C2(new_n368), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n356), .A2(new_n358), .ZN(new_n456));
  INV_X1    g255(.A(new_n300), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n365), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI211_X1 g257(.A(new_n300), .B(new_n364), .C1(new_n356), .C2(new_n358), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n453), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT92), .B1(new_n398), .B2(KEYINPUT6), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n393), .A2(KEYINPUT91), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n397), .B1(new_n392), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n402), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  AND4_X1   g265(.A1(KEYINPUT92), .A2(new_n392), .A3(KEYINPUT6), .A4(new_n401), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n462), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n461), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n447), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n389), .A2(new_n374), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n397), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n385), .A2(new_n375), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n473), .B(KEYINPUT40), .C1(new_n477), .C2(new_n479), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n482), .A2(new_n483), .B1(new_n463), .B2(new_n465), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n450), .A2(new_n451), .A3(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n441), .A2(new_n442), .A3(new_n421), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT93), .B(new_n433), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n443), .A2(new_n487), .A3(new_n422), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n428), .A2(KEYINPUT37), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT93), .B1(new_n491), .B2(new_n433), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT38), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n426), .A2(new_n335), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n419), .A2(new_n404), .A3(new_n420), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT37), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n489), .A2(new_n494), .A3(new_n433), .A4(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n498), .A2(new_n440), .A3(new_n444), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(new_n468), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n500), .A3(new_n366), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n453), .B2(new_n455), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n294), .A2(KEYINPUT36), .A3(new_n371), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n503), .A2(new_n504), .B1(new_n446), .B2(new_n460), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n472), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  XOR2_X1   g307(.A(G15gat), .B(G22gat), .Z(new_n509));
  INV_X1    g308(.A(G1gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n511), .B2(KEYINPUT98), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(G1gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n511), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n512), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT21), .ZN(new_n518));
  NAND2_X1  g317(.A1(G71gat), .A2(G78gat), .ZN(new_n519));
  OR2_X1    g318(.A1(G71gat), .A2(G78gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(G57gat), .B(G64gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT100), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n520), .A2(new_n519), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n526), .B(KEYINPUT100), .C1(new_n522), .C2(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n520), .A2(new_n522), .ZN(new_n529));
  INV_X1    g328(.A(new_n519), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(new_n521), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G183gat), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT101), .B(KEYINPUT21), .Z(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n528), .B2(new_n532), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G127gat), .B(G155gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G211gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n534), .B(new_n216), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n540), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n546));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n542), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n542), .B2(new_n545), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT102), .B(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(G85gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT7), .ZN(new_n556));
  INV_X1    g355(.A(G99gat), .ZN(new_n557));
  INV_X1    g356(.A(G106gat), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT8), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(new_n554), .A3(new_n556), .A4(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT15), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT95), .B(G29gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G36gat), .ZN(new_n571));
  OR3_X1    g370(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n572), .A2(KEYINPUT97), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(KEYINPUT97), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n569), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n571), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT94), .B1(new_n572), .B2(new_n575), .ZN(new_n580));
  OAI211_X1 g379(.A(KEYINPUT15), .B(new_n566), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(KEYINPUT17), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n577), .B2(new_n581), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n565), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n564), .A3(new_n562), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G190gat), .B(G218gat), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n591), .A2(KEYINPUT103), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n589), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n589), .B2(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(KEYINPUT103), .ZN(new_n597));
  XOR2_X1   g396(.A(G134gat), .B(G162gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR3_X1    g399(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n595), .B2(new_n596), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n517), .B1(new_n583), .B2(new_n585), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n516), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n517), .A2(KEYINPUT99), .A3(new_n577), .A4(new_n581), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n582), .B2(new_n516), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n612), .A3(new_n606), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n605), .B(KEYINPUT13), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n606), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT11), .B(G169gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G197gat), .ZN(new_n620));
  XOR2_X1   g419(.A(G113gat), .B(G141gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n609), .A2(new_n623), .A3(new_n616), .A4(new_n617), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n533), .A2(new_n565), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n528), .A2(new_n532), .A3(new_n564), .A4(new_n562), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(KEYINPUT104), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n533), .A2(new_n632), .A3(new_n565), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT10), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G230gat), .ZN(new_n637));
  OAI22_X1  g436(.A1(new_n634), .A2(new_n636), .B1(new_n637), .B2(new_n409), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n409), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n631), .A2(new_n639), .A3(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n231), .ZN(new_n643));
  INV_X1    g442(.A(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n628), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g448(.A1(new_n507), .A2(new_n551), .A3(new_n603), .A4(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n403), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT105), .B(G1gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1324gat));
  INV_X1    g453(.A(new_n452), .ZN(new_n655));
  NAND2_X1  g454(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n513), .A2(new_n508), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n650), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT106), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n650), .A2(new_n655), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G8gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(KEYINPUT106), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n661), .A2(new_n662), .A3(new_n664), .A4(new_n665), .ZN(G1325gat));
  NOR2_X1   g465(.A1(new_n453), .A2(new_n455), .ZN(new_n667));
  AOI21_X1  g466(.A(G15gat), .B1(new_n650), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n503), .A2(new_n504), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n650), .A2(G15gat), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n650), .A2(new_n460), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(new_n603), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n507), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n507), .A2(KEYINPUT44), .A3(new_n676), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n549), .A2(new_n550), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n649), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n651), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n570), .ZN(new_n686));
  INV_X1    g485(.A(new_n683), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n507), .A2(new_n676), .A3(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n688), .A2(new_n403), .A3(new_n570), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(G1328gat));
  NAND2_X1  g490(.A1(new_n684), .A2(new_n655), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G36gat), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n688), .A2(G36gat), .A3(new_n452), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1329gat));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n507), .B2(new_n676), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n678), .B(new_n603), .C1(new_n472), .C2(new_n506), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n699), .A2(G43gat), .A3(new_n670), .A4(new_n687), .ZN(new_n700));
  INV_X1    g499(.A(new_n667), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n688), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(G43gat), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g503(.A1(new_n699), .A2(G50gat), .A3(new_n460), .A4(new_n687), .ZN(new_n705));
  INV_X1    g504(.A(G50gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n688), .B2(new_n366), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT48), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n705), .A2(new_n713), .A3(new_n707), .A4(new_n708), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n712), .A3(new_n714), .ZN(G1331gat));
  NOR3_X1   g514(.A1(new_n682), .A2(new_n676), .A3(new_n627), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n507), .A2(new_n648), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n403), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT109), .B(G57gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1332gat));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n507), .A2(KEYINPUT110), .A3(new_n648), .A4(new_n716), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n452), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT111), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n727), .B(new_n728), .Z(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n717), .B2(new_n701), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n669), .A2(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n724), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n733), .ZN(new_n735));
  AOI211_X1 g534(.A(KEYINPUT112), .B(new_n735), .C1(new_n722), .C2(new_n723), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n731), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT50), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n739), .B(new_n731), .C1(new_n734), .C2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1334gat));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n460), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g542(.A1(new_n682), .A2(new_n628), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT113), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n648), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n681), .A2(new_n553), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n507), .A2(new_n676), .A3(new_n745), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT51), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n507), .A2(new_n745), .A3(new_n750), .A4(new_n676), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n749), .A2(new_n651), .A3(new_n648), .A4(new_n751), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n747), .A2(new_n651), .B1(new_n553), .B2(new_n752), .ZN(G1336gat));
  NOR2_X1   g552(.A1(new_n452), .A2(G92gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n749), .A2(new_n648), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n681), .A2(new_n452), .A3(new_n746), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(new_n552), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n759), .B(new_n755), .C1(new_n756), .C2(new_n552), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1337gat));
  NOR3_X1   g560(.A1(new_n681), .A2(new_n669), .A3(new_n746), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n749), .A2(new_n557), .A3(new_n648), .A4(new_n751), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n762), .A2(new_n557), .B1(new_n701), .B2(new_n763), .ZN(G1338gat));
  NOR4_X1   g563(.A1(new_n697), .A2(new_n698), .A3(new_n366), .A4(new_n746), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n558), .A3(new_n648), .A4(new_n751), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n765), .A2(new_n558), .B1(new_n766), .B2(new_n366), .ZN(new_n767));
  INV_X1    g566(.A(new_n746), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n679), .A2(new_n460), .A3(new_n680), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI221_X1 g573(.A(new_n770), .B1(new_n771), .B2(KEYINPUT53), .C1(new_n366), .C2(new_n766), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1339gat));
  INV_X1    g575(.A(new_n648), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n551), .A2(new_n603), .A3(new_n777), .A4(new_n628), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT115), .B1(new_n638), .B2(KEYINPUT54), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n631), .A2(new_n633), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n635), .ZN(new_n782));
  INV_X1    g581(.A(new_n636), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n639), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n638), .A3(KEYINPUT54), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n784), .A2(new_n638), .A3(KEYINPUT115), .A4(KEYINPUT54), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n645), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n779), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n780), .A2(new_n785), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n645), .A4(new_n787), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n789), .A2(new_n646), .A3(new_n627), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n613), .A2(new_n615), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n622), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT116), .B(new_n622), .C1(new_n793), .C2(new_n794), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n797), .A2(new_n626), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n648), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n603), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n789), .A2(new_n646), .A3(new_n791), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n803), .A2(new_n676), .A3(KEYINPUT117), .A4(new_n799), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n799), .A2(new_n789), .A3(new_n646), .A4(new_n791), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n603), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n778), .B1(new_n808), .B2(new_n682), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n452), .A2(new_n461), .A3(new_n651), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n627), .ZN(new_n812));
  MUX2_X1   g611(.A(new_n240), .B(G113gat), .S(new_n812), .Z(G1340gat));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n648), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n242), .A2(KEYINPUT118), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n811), .A2(new_n648), .B1(KEYINPUT118), .B2(new_n242), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n815), .ZN(G1341gat));
  NAND2_X1  g617(.A1(new_n811), .A2(new_n551), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(new_n249), .ZN(G1342gat));
  NAND2_X1  g619(.A1(new_n811), .A2(new_n676), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(KEYINPUT56), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT119), .Z(new_n823));
  AOI21_X1  g622(.A(G134gat), .B1(new_n821), .B2(KEYINPUT56), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(G1343gat));
  NAND3_X1  g624(.A1(new_n669), .A2(new_n651), .A3(new_n452), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT120), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n808), .A2(new_n682), .ZN(new_n828));
  INV_X1    g627(.A(new_n778), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n830), .B2(new_n460), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n809), .A2(new_n832), .A3(new_n366), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G141gat), .B1(new_n834), .B2(new_n628), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n809), .A2(new_n366), .A3(new_n826), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n303), .A3(new_n627), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n837), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n834), .A2(KEYINPUT121), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n830), .A2(KEYINPUT57), .A3(new_n460), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n832), .B1(new_n809), .B2(new_n366), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n842), .B1(new_n845), .B2(new_n827), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n627), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n840), .B1(new_n847), .B2(G141gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n839), .B1(new_n848), .B2(new_n838), .ZN(G1344gat));
  NAND3_X1  g648(.A1(new_n836), .A2(new_n306), .A3(new_n648), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT121), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n845), .A2(new_n842), .A3(new_n827), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n777), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(KEYINPUT59), .A3(new_n306), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n843), .A2(KEYINPUT122), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n833), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n676), .B1(new_n792), .B2(new_n800), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n806), .A2(new_n603), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n682), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n366), .B1(new_n829), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n862), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n856), .B(new_n858), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n648), .A3(new_n827), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n855), .B1(new_n868), .B2(G148gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n850), .B1(new_n854), .B2(new_n869), .ZN(G1345gat));
  AOI21_X1  g669(.A(G155gat), .B1(new_n836), .B2(new_n551), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n682), .B1(new_n851), .B2(new_n852), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n836), .B2(new_n676), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n603), .B1(new_n851), .B2(new_n852), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(G162gat), .ZN(G1347gat));
  NOR3_X1   g675(.A1(new_n809), .A2(new_n460), .A3(new_n701), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n452), .A2(new_n651), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT124), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n230), .A3(new_n627), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT125), .B1(new_n877), .B2(new_n878), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n877), .A2(KEYINPUT125), .A3(new_n878), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n628), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n882), .B1(new_n886), .B2(new_n230), .ZN(G1348gat));
  OAI21_X1  g686(.A(new_n231), .B1(new_n880), .B2(new_n777), .ZN(new_n888));
  INV_X1    g687(.A(new_n885), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n648), .B1(new_n889), .B2(new_n883), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n231), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(G1349gat));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n213), .A3(new_n551), .A4(new_n878), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT126), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n682), .B1(new_n884), .B2(new_n885), .ZN(new_n895));
  INV_X1    g694(.A(new_n262), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n894), .B(new_n899), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n208), .A3(new_n676), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n676), .B1(new_n889), .B2(new_n883), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(G190gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n903), .B2(G190gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G1351gat));
  AND2_X1   g706(.A1(new_n878), .A2(new_n669), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n867), .A2(new_n627), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G197gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n830), .A2(new_n460), .A3(new_n908), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(G197gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n628), .B2(new_n912), .ZN(G1352gat));
  NOR3_X1   g712(.A1(new_n911), .A2(G204gat), .A3(new_n777), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT62), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n867), .A2(new_n648), .A3(new_n908), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n644), .ZN(G1353gat));
  NAND3_X1  g716(.A1(new_n867), .A2(new_n551), .A3(new_n908), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G211gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT63), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n921), .A3(G211gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n911), .A2(G211gat), .A3(new_n682), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT127), .Z(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(G1354gat));
  NAND3_X1  g724(.A1(new_n867), .A2(new_n676), .A3(new_n908), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G218gat), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n603), .A2(G218gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n911), .B2(new_n928), .ZN(G1355gat));
endmodule


