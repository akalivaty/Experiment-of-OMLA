//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960;
  INV_X1    g000(.A(G1gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT88), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT90), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(KEYINPUT90), .A3(new_n205), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI211_X1 g010(.A(G1gat), .B(new_n205), .C1(KEYINPUT89), .C2(G8gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n205), .A2(G1gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214));
  NOR3_X1   g013(.A1(new_n213), .A2(new_n214), .A3(new_n209), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n212), .B1(new_n206), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G43gat), .B(G50gat), .Z(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n218), .B1(new_n225), .B2(KEYINPUT15), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(KEYINPUT15), .B2(new_n225), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(KEYINPUT15), .A3(new_n218), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n217), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n229), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n211), .A3(new_n216), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n227), .A3(new_n229), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n235), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(new_n233), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n232), .A2(KEYINPUT18), .A3(new_n233), .A4(new_n235), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n238), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G197gat), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT11), .B(G169gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n238), .A2(new_n243), .A3(new_n250), .A4(new_n244), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT23), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT24), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n260), .B(new_n267), .C1(new_n273), .C2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n281), .A2(new_n276), .A3(new_n277), .A4(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT25), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n263), .B2(new_n266), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n256), .B1(KEYINPUT23), .B2(new_n264), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n279), .A2(KEYINPUT25), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n265), .B1(KEYINPUT26), .B2(new_n263), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n258), .A2(new_n259), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(KEYINPUT26), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G183gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n274), .A2(KEYINPUT27), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n274), .A2(KEYINPUT27), .ZN(new_n297));
  AOI21_X1  g096(.A(G190gat), .B1(new_n297), .B2(KEYINPUT67), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT28), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n300), .A2(KEYINPUT28), .A3(new_n275), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n291), .B(new_n272), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n288), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G226gat), .A2(G233gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n288), .B2(new_n302), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT22), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n308), .A3(new_n312), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n305), .B(new_n318), .C1(new_n304), .C2(new_n306), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G8gat), .B(G36gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G64gat), .B(G92gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n322), .A2(KEYINPUT30), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n322), .B2(new_n326), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n326), .B2(new_n322), .ZN(new_n331));
  INV_X1    g130(.A(G134gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(G127gat), .ZN(new_n333));
  INV_X1    g132(.A(G127gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(G134gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT69), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G120gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G113gat), .ZN(new_n338));
  INV_X1    g137(.A(G113gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G120gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT1), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n334), .A2(G134gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n332), .A2(G127gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n336), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT68), .ZN(new_n347));
  OR3_X1    g146(.A1(new_n332), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n347), .B(new_n348), .C1(KEYINPUT1), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  INV_X1    g150(.A(G155gat), .ZN(new_n352));
  INV_X1    g151(.A(G162gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G141gat), .B(G148gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n351), .B(new_n354), .C1(new_n355), .C2(KEYINPUT2), .ZN(new_n356));
  XOR2_X1   g155(.A(G141gat), .B(G148gat), .Z(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n351), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(KEYINPUT2), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n346), .A2(new_n350), .A3(new_n356), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT76), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n365), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n362), .B2(KEYINPUT75), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n371));
  AOI211_X1 g170(.A(new_n371), .B(KEYINPUT76), .C1(new_n361), .C2(KEYINPUT4), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n360), .A2(new_n356), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n356), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n346), .A2(new_n350), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT39), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n360), .A2(new_n356), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(new_n379), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT83), .A3(new_n383), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT39), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT83), .B1(new_n387), .B2(new_n383), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n380), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(new_n368), .B2(new_n373), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n393), .B2(new_n383), .ZN(new_n394));
  XOR2_X1   g193(.A(G1gat), .B(G29gat), .Z(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT40), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n328), .B(new_n331), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT5), .B1(new_n387), .B2(new_n383), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT73), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT73), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n406), .B(KEYINPUT5), .C1(new_n387), .C2(new_n383), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n369), .A2(new_n362), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(new_n383), .A3(new_n380), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n380), .A2(new_n412), .A3(new_n383), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT77), .B1(new_n374), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n374), .A2(KEYINPUT77), .A3(new_n414), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n411), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n421));
  AOI211_X1 g220(.A(new_n421), .B(new_n413), .C1(new_n368), .C2(new_n373), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n410), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n400), .B1(new_n423), .B2(KEYINPUT86), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n403), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n401), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n385), .A2(new_n394), .A3(KEYINPUT84), .A4(new_n400), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n402), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT85), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n427), .A2(KEYINPUT85), .A3(new_n402), .A4(new_n428), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n423), .A2(new_n399), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n423), .A2(KEYINPUT87), .A3(new_n399), .A4(new_n435), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n420), .A2(new_n424), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n400), .B(new_n410), .C1(new_n415), .C2(new_n422), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n434), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n322), .A2(KEYINPUT37), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n325), .B1(new_n322), .B2(KEYINPUT37), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n322), .A2(new_n326), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n440), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(G50gat), .ZN(new_n455));
  XOR2_X1   g254(.A(G78gat), .B(G106gat), .Z(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(G228gat), .A2(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459));
  INV_X1    g258(.A(new_n317), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n314), .B1(new_n312), .B2(new_n308), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n386), .B1(new_n462), .B2(new_n377), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n318), .B1(new_n378), .B2(new_n459), .ZN(new_n464));
  OAI211_X1 g263(.A(KEYINPUT80), .B(new_n458), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n378), .A2(new_n459), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n319), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT29), .B1(new_n316), .B2(new_n317), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n375), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(G22gat), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n457), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n465), .A2(G22gat), .A3(new_n472), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(new_n473), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n479), .B(new_n457), .C1(new_n473), .C2(new_n474), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n476), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n433), .A2(new_n453), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n331), .A2(new_n328), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n423), .A2(new_n399), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n434), .A3(new_n442), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n488), .B2(new_n436), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  INV_X1    g289(.A(new_n379), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n303), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G227gat), .ZN(new_n493));
  INV_X1    g292(.A(G233gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n288), .A2(new_n302), .A3(new_n379), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT32), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT70), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G43gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT33), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n497), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n497), .B(KEYINPUT32), .C1(new_n504), .C2(new_n503), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n288), .A2(new_n302), .A3(new_n379), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n379), .B1(new_n288), .B2(new_n302), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n511), .B1(new_n514), .B2(new_n495), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n492), .A2(new_n496), .ZN(new_n516));
  INV_X1    g315(.A(new_n495), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n510), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n515), .A2(new_n518), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n508), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n507), .B(new_n508), .C1(KEYINPUT71), .C2(new_n519), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT36), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n490), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n485), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n488), .A2(new_n436), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n527), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n483), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n486), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n520), .A2(new_n523), .B1(new_n331), .B2(new_n328), .ZN(new_n539));
  INV_X1    g338(.A(new_n482), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT35), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n438), .A2(new_n439), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n443), .B1(new_n420), .B2(new_n424), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n539), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n255), .B1(new_n532), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G99gat), .B(G106gat), .Z(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT7), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n554));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n555), .A2(KEYINPUT8), .ZN(new_n556));
  NOR2_X1   g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT97), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n550), .B(new_n553), .C1(new_n558), .C2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n550), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n562), .ZN(new_n565));
  INV_X1    g364(.A(new_n553), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI22_X1  g366(.A1(new_n230), .A2(new_n231), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n563), .ZN(new_n569));
  AND2_X1   g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n569), .A2(new_n234), .B1(KEYINPUT41), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(KEYINPUT98), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n549), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI211_X1 g376(.A(new_n574), .B(new_n548), .C1(new_n568), .C2(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(KEYINPUT98), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n576), .B2(new_n578), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT92), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n590), .B(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n217), .B1(new_n587), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  XOR2_X1   g397(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT20), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n596), .B(new_n597), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n607), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n607), .B2(new_n610), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n586), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n565), .A2(new_n566), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n550), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n590), .B(new_n593), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n556), .A2(new_n554), .A3(new_n557), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n561), .A2(KEYINPUT97), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n564), .B(new_n566), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n621), .A2(new_n622), .A3(KEYINPUT10), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT100), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n569), .A2(new_n628), .A3(KEYINPUT10), .A4(new_n622), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(KEYINPUT99), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n631), .B(new_n622), .C1(new_n567), .C2(new_n563), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n621), .B(new_n625), .C1(new_n595), .C2(KEYINPUT99), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT10), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G230gat), .ZN(new_n635));
  OAI22_X1  g434(.A1(new_n630), .A2(new_n634), .B1(new_n635), .B2(new_n494), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n494), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n637), .A3(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n619), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n619), .ZN(new_n642));
  AOI211_X1 g441(.A(KEYINPUT101), .B(new_n642), .C1(new_n636), .C2(new_n638), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n616), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n616), .A2(KEYINPUT102), .A3(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n533), .A2(KEYINPUT103), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n533), .A2(KEYINPUT103), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n547), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n547), .A2(new_n650), .ZN(new_n656));
  OR3_X1    g455(.A1(new_n656), .A2(KEYINPUT104), .A3(new_n536), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT104), .B1(new_n656), .B2(new_n536), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(G8gat), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n656), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT16), .B(G8gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT105), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n660), .A2(KEYINPUT42), .A3(new_n486), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n657), .B2(new_n658), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n659), .B(new_n664), .C1(new_n665), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g465(.A(new_n520), .ZN(new_n667));
  INV_X1    g466(.A(new_n523), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n660), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n530), .A2(G15gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT106), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n660), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n484), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n583), .A2(new_n585), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n532), .B2(new_n546), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n614), .A2(new_n615), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(new_n255), .A3(new_n644), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n223), .A3(new_n653), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n542), .A2(new_n539), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n440), .B2(new_n445), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT35), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n489), .B2(new_n535), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT108), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n538), .A2(new_n692), .A3(new_n545), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n691), .A2(new_n693), .B1(new_n485), .B2(new_n531), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n686), .B1(new_n694), .B2(new_n678), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n532), .A2(new_n546), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(KEYINPUT44), .A3(new_n586), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(new_n681), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n653), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n700), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n682), .A2(new_n219), .A3(new_n486), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n703));
  OAI21_X1  g502(.A(G36gat), .B1(new_n698), .B2(new_n536), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n695), .A2(new_n530), .A3(new_n697), .A4(new_n681), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G43gat), .ZN(new_n708));
  INV_X1    g507(.A(G43gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n682), .A2(new_n709), .A3(new_n670), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1330gat));
  NAND4_X1  g514(.A1(new_n695), .A2(new_n483), .A3(new_n697), .A4(new_n681), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G50gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n484), .A2(G50gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n682), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT109), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n682), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n717), .A2(new_n720), .A3(KEYINPUT48), .A4(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n717), .A2(new_n719), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g524(.A1(new_n616), .A2(new_n255), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n694), .A2(new_n645), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n653), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n694), .A2(new_n726), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n536), .A2(new_n645), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  INV_X1    g534(.A(new_n727), .ZN(new_n736));
  OAI21_X1  g535(.A(G71gat), .B1(new_n736), .B2(new_n529), .ZN(new_n737));
  INV_X1    g536(.A(G71gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n727), .A2(new_n738), .A3(new_n670), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n737), .B2(new_n739), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n483), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT111), .B(G78gat), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n744), .B(new_n745), .Z(G1335gat));
  NOR2_X1   g545(.A1(new_n680), .A2(new_n254), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n645), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n695), .A2(new_n697), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n699), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n691), .A2(new_n693), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n678), .B1(new_n752), .B2(new_n532), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n753), .B2(new_n747), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n694), .A2(new_n755), .A3(new_n678), .A4(new_n748), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n644), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n653), .A2(new_n559), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(G1336gat));
  NAND4_X1  g558(.A1(new_n695), .A2(new_n486), .A3(new_n697), .A4(new_n749), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n731), .A2(new_n560), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT112), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n754), .B2(new_n756), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n750), .B2(new_n529), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n669), .A2(G99gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n757), .B2(new_n771), .ZN(G1338gat));
  NOR2_X1   g571(.A1(new_n484), .A2(G106gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n644), .B(new_n773), .C1(new_n754), .C2(new_n756), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n695), .A2(new_n483), .A3(new_n697), .A4(new_n749), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(new_n680), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n632), .A2(new_n633), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT10), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n627), .A2(new_n629), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n637), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n783), .A2(new_n784), .B1(new_n627), .B2(new_n629), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(KEYINPUT113), .A3(new_n637), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n789), .A2(new_n791), .A3(KEYINPUT54), .A4(new_n636), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n790), .A2(new_n637), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n619), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n636), .A2(new_n638), .A3(new_n619), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n795), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n798), .A2(new_n254), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n240), .A2(new_n242), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n233), .B1(new_n232), .B2(new_n235), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n249), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT114), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n806), .B(new_n249), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n644), .A2(new_n253), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n586), .B1(new_n801), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n800), .A2(new_n799), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n805), .A2(new_n253), .A3(new_n807), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n678), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n811), .A2(new_n798), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n782), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n616), .A2(new_n255), .A3(new_n645), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n817), .A2(new_n535), .A3(new_n653), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n536), .A3(new_n254), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n484), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n653), .A2(new_n539), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n255), .A2(new_n339), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n819), .A2(new_n339), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  AOI21_X1  g623(.A(new_n337), .B1(new_n822), .B2(new_n644), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n825), .B(KEYINPUT115), .Z(new_n826));
  NAND2_X1  g625(.A1(new_n818), .A2(new_n536), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n644), .A2(new_n337), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT116), .Z(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(G1341gat));
  INV_X1    g629(.A(new_n822), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n334), .A3(new_n782), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n827), .A2(KEYINPUT117), .A3(new_n782), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(G127gat), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT117), .B1(new_n827), .B2(new_n782), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(G1342gat));
  NOR2_X1   g635(.A1(new_n486), .A2(new_n678), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT118), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(G134gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n831), .B2(new_n678), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT119), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n841), .A2(new_n842), .A3(new_n846), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1343gat));
  INV_X1    g647(.A(new_n816), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n811), .A2(new_n798), .A3(new_n813), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n812), .A2(new_n643), .A3(new_n641), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n796), .A2(new_n797), .B1(new_n252), .B2(new_n253), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n811), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n853), .B2(new_n586), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n849), .B1(new_n854), .B2(new_n782), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n529), .A2(new_n483), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n855), .A2(new_n699), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n536), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(G141gat), .A3(new_n255), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n699), .A2(new_n486), .A3(new_n530), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n817), .B2(new_n483), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n862), .B(new_n484), .C1(new_n815), .C2(new_n816), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT120), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n866), .B(new_n860), .C1(new_n861), .C2(new_n863), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n867), .A3(new_n254), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n859), .B1(new_n868), .B2(G141gat), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n864), .A2(new_n255), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n859), .A2(KEYINPUT58), .ZN(new_n873));
  OAI22_X1  g672(.A1(new_n869), .A2(new_n870), .B1(new_n872), .B2(new_n873), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n645), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(G148gat), .ZN(new_n877));
  INV_X1    g676(.A(G148gat), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n650), .A2(new_n255), .B1(new_n854), .B2(new_n782), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n862), .B1(new_n879), .B2(new_n484), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n817), .A2(KEYINPUT57), .A3(new_n483), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n644), .A3(new_n860), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(KEYINPUT59), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n865), .A2(new_n867), .A3(new_n876), .A4(new_n644), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n782), .A2(new_n352), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n865), .A2(new_n867), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n352), .B1(new_n858), .B2(new_n782), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n888), .A2(KEYINPUT121), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1346gat));
  NOR2_X1   g693(.A1(new_n838), .A2(G162gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n857), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT122), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n865), .A2(new_n867), .A3(new_n586), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n353), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n855), .A2(new_n653), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n535), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n536), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n254), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n653), .A2(new_n536), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n670), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n820), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n255), .A2(new_n261), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1348gat));
  INV_X1    g707(.A(new_n906), .ZN(new_n909));
  OAI21_X1  g708(.A(G176gat), .B1(new_n909), .B2(new_n645), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n731), .A2(new_n262), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n901), .B2(new_n911), .ZN(G1349gat));
  NAND3_X1  g711(.A1(new_n902), .A2(new_n300), .A3(new_n680), .ZN(new_n913));
  OAI21_X1  g712(.A(G183gat), .B1(new_n909), .B2(new_n782), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n275), .A3(new_n586), .ZN(new_n918));
  OAI21_X1  g717(.A(G190gat), .B1(new_n909), .B2(new_n678), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n856), .A2(new_n536), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n900), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n254), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n904), .A2(new_n529), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n880), .B2(new_n881), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n254), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n900), .A2(new_n933), .A3(new_n644), .A4(new_n923), .ZN(new_n934));
  XNOR2_X1  g733(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n934), .B(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n930), .A2(new_n644), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n933), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n934), .B(new_n935), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n933), .B1(new_n930), .B2(new_n644), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT126), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n310), .A3(new_n680), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n310), .B1(new_n930), .B2(new_n680), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(KEYINPUT63), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(KEYINPUT63), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1354gat));
  NOR2_X1   g748(.A1(new_n678), .A2(G218gat), .ZN(new_n950));
  INV_X1    g749(.A(new_n926), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n930), .A2(new_n586), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n953), .B(KEYINPUT127), .C1(new_n954), .C2(new_n311), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  INV_X1    g755(.A(new_n950), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n925), .B2(new_n926), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n311), .B1(new_n930), .B2(new_n586), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n955), .A2(new_n960), .ZN(G1355gat));
endmodule


