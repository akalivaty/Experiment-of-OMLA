

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721;

  NOR2_X1 U368 ( .A1(n639), .A2(n669), .ZN(n559) );
  AND2_X1 U369 ( .A1(n489), .A2(n488), .ZN(n490) );
  INV_X1 U370 ( .A(n676), .ZN(n639) );
  NAND2_X1 U371 ( .A1(n472), .A2(n474), .ZN(n676) );
  AND2_X2 U372 ( .A1(n457), .A2(n564), .ZN(n458) );
  AND2_X2 U373 ( .A1(n463), .A2(n554), .ZN(n484) );
  AND2_X1 U374 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U375 ( .A(n454), .B(n453), .ZN(n649) );
  NOR2_X1 U376 ( .A1(n514), .A2(n676), .ZN(n454) );
  NOR2_X1 U377 ( .A1(n603), .A2(n602), .ZN(n551) );
  XNOR2_X1 U378 ( .A(n366), .B(KEYINPUT25), .ZN(n367) );
  XNOR2_X1 U379 ( .A(n358), .B(G140), .ZN(n378) );
  XNOR2_X1 U380 ( .A(KEYINPUT10), .B(n409), .ZN(n708) );
  NOR2_X2 U381 ( .A1(n691), .A2(G902), .ZN(n368) );
  INV_X2 U382 ( .A(n597), .ZN(n564) );
  XNOR2_X1 U383 ( .A(n440), .B(n651), .ZN(n441) );
  NOR2_X1 U384 ( .A1(n505), .A2(n504), .ZN(n507) );
  XNOR2_X1 U385 ( .A(n422), .B(n421), .ZN(n468) );
  XNOR2_X1 U386 ( .A(n570), .B(n569), .ZN(n698) );
  INV_X1 U387 ( .A(KEYINPUT45), .ZN(n569) );
  XNOR2_X1 U388 ( .A(G107), .B(G122), .ZN(n413) );
  XNOR2_X1 U389 ( .A(n708), .B(n437), .ZN(n438) );
  NOR2_X1 U390 ( .A1(n493), .A2(n467), .ZN(n400) );
  BUF_X1 U391 ( .A(n468), .Z(n511) );
  INV_X1 U392 ( .A(KEYINPUT120), .ZN(n633) );
  NOR2_X1 U393 ( .A1(n583), .A2(n694), .ZN(n585) );
  XNOR2_X1 U394 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U395 ( .A(n399), .B(n398), .ZN(n493) );
  NOR2_X1 U396 ( .A1(n405), .A2(n522), .ZN(n345) );
  XOR2_X1 U397 ( .A(n490), .B(KEYINPUT82), .Z(n346) );
  INV_X2 U398 ( .A(G953), .ZN(n405) );
  OR2_X1 U399 ( .A1(G902), .A2(G237), .ZN(n347) );
  XNOR2_X1 U400 ( .A(G143), .B(G128), .ZN(n401) );
  XOR2_X1 U401 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n348) );
  AND2_X1 U402 ( .A1(n536), .A2(n598), .ZN(n349) );
  XOR2_X1 U403 ( .A(n588), .B(n587), .Z(n350) );
  XNOR2_X1 U404 ( .A(KEYINPUT17), .B(KEYINPUT92), .ZN(n407) );
  NOR2_X1 U405 ( .A1(n502), .A2(n501), .ZN(n503) );
  INV_X2 U406 ( .A(KEYINPUT4), .ZN(n379) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n428) );
  XNOR2_X1 U408 ( .A(n707), .B(G101), .ZN(n404) );
  NAND2_X1 U409 ( .A1(n598), .A2(n458), .ZN(n492) );
  XNOR2_X1 U410 ( .A(n394), .B(n393), .ZN(n395) );
  NOR2_X1 U411 ( .A1(n648), .A2(n549), .ZN(n550) );
  XNOR2_X1 U412 ( .A(n444), .B(n377), .ZN(n393) );
  XNOR2_X1 U413 ( .A(n396), .B(n395), .ZN(n586) );
  NOR2_X1 U414 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U415 ( .A(n520), .B(n519), .ZN(n622) );
  XNOR2_X1 U416 ( .A(n439), .B(n438), .ZN(n652) );
  NOR2_X1 U417 ( .A1(n622), .A2(n556), .ZN(n531) );
  XNOR2_X1 U418 ( .A(n442), .B(n441), .ZN(n475) );
  AND2_X1 U419 ( .A1(n387), .A2(n554), .ZN(n477) );
  INV_X1 U420 ( .A(n694), .ZN(n589) );
  INV_X1 U421 ( .A(KEYINPUT40), .ZN(n453) );
  INV_X1 U422 ( .A(KEYINPUT121), .ZN(n584) );
  XNOR2_X1 U423 ( .A(n585), .B(n584), .ZN(G54) );
  XOR2_X1 U424 ( .A(KEYINPUT20), .B(KEYINPUT97), .Z(n352) );
  XNOR2_X1 U425 ( .A(G902), .B(KEYINPUT15), .ZN(n572) );
  NAND2_X1 U426 ( .A1(G234), .A2(n572), .ZN(n351) );
  XNOR2_X1 U427 ( .A(n352), .B(n351), .ZN(n365) );
  AND2_X1 U428 ( .A1(n365), .A2(G221), .ZN(n353) );
  XNOR2_X1 U429 ( .A(n353), .B(KEYINPUT21), .ZN(n598) );
  XOR2_X1 U430 ( .A(G110), .B(G119), .Z(n355) );
  XNOR2_X1 U431 ( .A(G128), .B(G137), .ZN(n354) );
  XNOR2_X1 U432 ( .A(n355), .B(n354), .ZN(n364) );
  XOR2_X1 U433 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n357) );
  NAND2_X1 U434 ( .A1(G234), .A2(n405), .ZN(n356) );
  XNOR2_X1 U435 ( .A(n357), .B(n356), .ZN(n446) );
  NAND2_X1 U436 ( .A1(n446), .A2(G221), .ZN(n360) );
  INV_X1 U437 ( .A(KEYINPUT68), .ZN(n358) );
  XOR2_X1 U438 ( .A(n378), .B(KEYINPUT96), .Z(n359) );
  XNOR2_X1 U439 ( .A(n360), .B(n359), .ZN(n362) );
  XNOR2_X2 U440 ( .A(G146), .B(G125), .ZN(n409) );
  XNOR2_X1 U441 ( .A(n708), .B(n348), .ZN(n361) );
  XNOR2_X1 U442 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U443 ( .A(n364), .B(n363), .ZN(n691) );
  NAND2_X1 U444 ( .A1(G217), .A2(n365), .ZN(n366) );
  XNOR2_X2 U445 ( .A(n368), .B(n367), .ZN(n597) );
  NAND2_X1 U446 ( .A1(n598), .A2(n597), .ZN(n602) );
  INV_X1 U447 ( .A(n602), .ZN(n375) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n369) );
  XNOR2_X1 U449 ( .A(n369), .B(KEYINPUT14), .ZN(n371) );
  NAND2_X1 U450 ( .A1(n371), .A2(G952), .ZN(n628) );
  INV_X1 U451 ( .A(n628), .ZN(n370) );
  NAND2_X1 U452 ( .A1(n370), .A2(n405), .ZN(n523) );
  INV_X1 U453 ( .A(G900), .ZN(n373) );
  NAND2_X1 U454 ( .A1(n371), .A2(G902), .ZN(n372) );
  XOR2_X1 U455 ( .A(KEYINPUT95), .B(n372), .Z(n522) );
  NAND2_X1 U456 ( .A1(n373), .A2(n345), .ZN(n374) );
  NAND2_X1 U457 ( .A1(n523), .A2(n374), .ZN(n457) );
  AND2_X1 U458 ( .A1(n375), .A2(n457), .ZN(n387) );
  XNOR2_X1 U459 ( .A(n401), .B(G134), .ZN(n444) );
  XNOR2_X1 U460 ( .A(G137), .B(G131), .ZN(n376) );
  XNOR2_X1 U461 ( .A(n376), .B(KEYINPUT69), .ZN(n377) );
  XNOR2_X1 U462 ( .A(n393), .B(n378), .ZN(n711) );
  XNOR2_X2 U463 ( .A(n379), .B(KEYINPUT67), .ZN(n707) );
  XNOR2_X1 U464 ( .A(n404), .B(G146), .ZN(n394) );
  NAND2_X1 U465 ( .A1(n405), .A2(G227), .ZN(n380) );
  XNOR2_X1 U466 ( .A(n380), .B(G107), .ZN(n381) );
  XNOR2_X1 U467 ( .A(G110), .B(G104), .ZN(n415) );
  XNOR2_X1 U468 ( .A(n381), .B(n415), .ZN(n382) );
  XNOR2_X1 U469 ( .A(n394), .B(n382), .ZN(n383) );
  XNOR2_X1 U470 ( .A(n711), .B(n383), .ZN(n579) );
  INV_X1 U471 ( .A(G902), .ZN(n397) );
  NAND2_X1 U472 ( .A1(n579), .A2(n397), .ZN(n386) );
  XNOR2_X1 U473 ( .A(KEYINPUT72), .B(G469), .ZN(n384) );
  XNOR2_X1 U474 ( .A(n384), .B(KEYINPUT71), .ZN(n385) );
  XNOR2_X2 U475 ( .A(n386), .B(n385), .ZN(n499) );
  INV_X1 U476 ( .A(n499), .ZN(n554) );
  XNOR2_X1 U477 ( .A(KEYINPUT3), .B(G119), .ZN(n388) );
  XNOR2_X1 U478 ( .A(n388), .B(G113), .ZN(n414) );
  XNOR2_X1 U479 ( .A(G116), .B(KEYINPUT5), .ZN(n389) );
  XNOR2_X1 U480 ( .A(n414), .B(n389), .ZN(n392) );
  NAND2_X1 U481 ( .A1(n428), .A2(G210), .ZN(n390) );
  XNOR2_X1 U482 ( .A(n390), .B(KEYINPUT98), .ZN(n391) );
  XNOR2_X1 U483 ( .A(n392), .B(n391), .ZN(n396) );
  NAND2_X1 U484 ( .A1(n586), .A2(n397), .ZN(n399) );
  XNOR2_X1 U485 ( .A(KEYINPUT99), .B(G472), .ZN(n398) );
  XNOR2_X1 U486 ( .A(KEYINPUT76), .B(n347), .ZN(n419) );
  NAND2_X1 U487 ( .A1(n419), .A2(G214), .ZN(n616) );
  INV_X1 U488 ( .A(n616), .ZN(n467) );
  XNOR2_X1 U489 ( .A(n400), .B(KEYINPUT30), .ZN(n478) );
  NAND2_X1 U490 ( .A1(n477), .A2(n478), .ZN(n424) );
  XNOR2_X1 U491 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n402) );
  XNOR2_X1 U492 ( .A(n401), .B(n402), .ZN(n403) );
  XNOR2_X1 U493 ( .A(n404), .B(n403), .ZN(n411) );
  NAND2_X1 U494 ( .A1(n405), .A2(G224), .ZN(n406) );
  XNOR2_X1 U495 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U496 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U497 ( .A(n411), .B(n410), .ZN(n418) );
  INV_X1 U498 ( .A(G116), .ZN(n412) );
  XNOR2_X1 U499 ( .A(n413), .B(n412), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n414), .B(n447), .ZN(n417) );
  XNOR2_X1 U501 ( .A(n415), .B(KEYINPUT16), .ZN(n416) );
  XNOR2_X1 U502 ( .A(n417), .B(n416), .ZN(n695) );
  XNOR2_X1 U503 ( .A(n418), .B(n695), .ZN(n658) );
  NAND2_X1 U504 ( .A1(n658), .A2(n572), .ZN(n422) );
  NAND2_X1 U505 ( .A1(n419), .A2(G210), .ZN(n420) );
  XNOR2_X1 U506 ( .A(n420), .B(KEYINPUT80), .ZN(n421) );
  XNOR2_X1 U507 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n423) );
  XNOR2_X1 U508 ( .A(n511), .B(n423), .ZN(n614) );
  NOR2_X1 U509 ( .A1(n424), .A2(n614), .ZN(n425) );
  XNOR2_X1 U510 ( .A(n425), .B(KEYINPUT39), .ZN(n514) );
  XOR2_X1 U511 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n427) );
  XNOR2_X1 U512 ( .A(G140), .B(G104), .ZN(n426) );
  XNOR2_X1 U513 ( .A(n427), .B(n426), .ZN(n430) );
  NAND2_X1 U514 ( .A1(n428), .A2(G214), .ZN(n429) );
  XNOR2_X1 U515 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U516 ( .A(G122), .B(G113), .Z(n432) );
  XNOR2_X1 U517 ( .A(G131), .B(G143), .ZN(n431) );
  XNOR2_X1 U518 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U519 ( .A(n434), .B(n433), .ZN(n439) );
  XOR2_X1 U520 ( .A(KEYINPUT104), .B(KEYINPUT102), .Z(n436) );
  XNOR2_X1 U521 ( .A(KEYINPUT105), .B(KEYINPUT11), .ZN(n435) );
  XNOR2_X1 U522 ( .A(n436), .B(n435), .ZN(n437) );
  NOR2_X1 U523 ( .A1(G902), .A2(n652), .ZN(n442) );
  XNOR2_X1 U524 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n440) );
  INV_X1 U525 ( .A(G475), .ZN(n651) );
  XNOR2_X1 U526 ( .A(n475), .B(KEYINPUT107), .ZN(n472) );
  XOR2_X1 U527 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n443) );
  XNOR2_X1 U528 ( .A(n443), .B(KEYINPUT108), .ZN(n445) );
  XNOR2_X1 U529 ( .A(n445), .B(n444), .ZN(n450) );
  NAND2_X1 U530 ( .A1(G217), .A2(n446), .ZN(n448) );
  XNOR2_X1 U531 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U532 ( .A(n450), .B(n449), .ZN(n687) );
  OR2_X1 U533 ( .A1(n687), .A2(G902), .ZN(n452) );
  XNOR2_X1 U534 ( .A(KEYINPUT109), .B(G478), .ZN(n451) );
  XNOR2_X1 U535 ( .A(n452), .B(n451), .ZN(n474) );
  AND2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n536) );
  INV_X1 U537 ( .A(n536), .ZN(n618) );
  NOR2_X1 U538 ( .A1(n618), .A2(n467), .ZN(n455) );
  INV_X1 U539 ( .A(n614), .ZN(n617) );
  NAND2_X1 U540 ( .A1(n455), .A2(n617), .ZN(n456) );
  XNOR2_X1 U541 ( .A(n456), .B(KEYINPUT41), .ZN(n610) );
  INV_X1 U542 ( .A(n493), .ZN(n460) );
  INV_X1 U543 ( .A(n492), .ZN(n459) );
  NAND2_X1 U544 ( .A1(n460), .A2(n459), .ZN(n462) );
  INV_X1 U545 ( .A(KEYINPUT28), .ZN(n461) );
  XNOR2_X1 U546 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U547 ( .A1(n610), .A2(n484), .ZN(n465) );
  XNOR2_X1 U548 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n464) );
  XNOR2_X1 U549 ( .A(n465), .B(n464), .ZN(n644) );
  NAND2_X1 U550 ( .A1(n649), .A2(n644), .ZN(n466) );
  XNOR2_X1 U551 ( .A(n466), .B(KEYINPUT46), .ZN(n505) );
  OR2_X2 U552 ( .A1(n468), .A2(n467), .ZN(n471) );
  INV_X1 U553 ( .A(KEYINPUT77), .ZN(n469) );
  XNOR2_X1 U554 ( .A(n469), .B(KEYINPUT19), .ZN(n470) );
  XNOR2_X2 U555 ( .A(n471), .B(n470), .ZN(n526) );
  NOR2_X1 U556 ( .A1(n472), .A2(n474), .ZN(n669) );
  INV_X1 U557 ( .A(n559), .ZN(n613) );
  AND2_X1 U558 ( .A1(n526), .A2(n613), .ZN(n473) );
  NAND2_X1 U559 ( .A1(n484), .A2(n473), .ZN(n491) );
  NAND2_X1 U560 ( .A1(n491), .A2(KEYINPUT47), .ZN(n483) );
  INV_X1 U561 ( .A(KEYINPUT83), .ZN(n481) );
  NOR2_X1 U562 ( .A1(n475), .A2(n474), .ZN(n532) );
  INV_X1 U563 ( .A(n532), .ZN(n476) );
  NOR2_X1 U564 ( .A1(n476), .A2(n511), .ZN(n480) );
  AND2_X1 U565 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U566 ( .A1(n480), .A2(n479), .ZN(n647) );
  AND2_X1 U567 ( .A1(n481), .A2(n647), .ZN(n482) );
  NAND2_X1 U568 ( .A1(n483), .A2(n482), .ZN(n489) );
  NAND2_X1 U569 ( .A1(n484), .A2(n526), .ZN(n638) );
  NAND2_X1 U570 ( .A1(KEYINPUT83), .A2(KEYINPUT47), .ZN(n485) );
  NOR2_X1 U571 ( .A1(n559), .A2(n485), .ZN(n486) );
  AND2_X1 U572 ( .A1(n647), .A2(n486), .ZN(n487) );
  NAND2_X1 U573 ( .A1(n638), .A2(n487), .ZN(n488) );
  NOR2_X1 U574 ( .A1(n491), .A2(KEYINPUT47), .ZN(n502) );
  NOR2_X1 U575 ( .A1(n676), .A2(n492), .ZN(n494) );
  XNOR2_X1 U576 ( .A(n493), .B(KEYINPUT6), .ZN(n561) );
  NAND2_X1 U577 ( .A1(n494), .A2(n561), .ZN(n495) );
  XNOR2_X1 U578 ( .A(n495), .B(KEYINPUT111), .ZN(n496) );
  NAND2_X1 U579 ( .A1(n496), .A2(n616), .ZN(n508) );
  NOR2_X1 U580 ( .A1(n508), .A2(n511), .ZN(n497) );
  XNOR2_X1 U581 ( .A(n497), .B(KEYINPUT36), .ZN(n500) );
  XNOR2_X1 U582 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n498) );
  XNOR2_X2 U583 ( .A(n499), .B(n498), .ZN(n542) );
  NAND2_X1 U584 ( .A1(n500), .A2(n542), .ZN(n681) );
  INV_X1 U585 ( .A(n681), .ZN(n501) );
  NAND2_X1 U586 ( .A1(n346), .A2(n503), .ZN(n504) );
  XOR2_X1 U587 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n506) );
  XNOR2_X1 U588 ( .A(n507), .B(n506), .ZN(n517) );
  XNOR2_X1 U589 ( .A(KEYINPUT43), .B(KEYINPUT112), .ZN(n510) );
  NOR2_X1 U590 ( .A1(n508), .A2(n542), .ZN(n509) );
  XOR2_X1 U591 ( .A(n510), .B(n509), .Z(n512) );
  NAND2_X1 U592 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U593 ( .A(KEYINPUT113), .B(n513), .Z(n720) );
  INV_X1 U594 ( .A(n514), .ZN(n515) );
  NAND2_X1 U595 ( .A1(n515), .A2(n669), .ZN(n683) );
  NAND2_X1 U596 ( .A1(n720), .A2(n683), .ZN(n516) );
  NOR2_X2 U597 ( .A1(n517), .A2(n516), .ZN(n573) );
  NAND2_X1 U598 ( .A1(n573), .A2(KEYINPUT2), .ZN(n518) );
  XNOR2_X1 U599 ( .A(n518), .B(KEYINPUT86), .ZN(n571) );
  INV_X1 U600 ( .A(n542), .ZN(n603) );
  NAND2_X1 U601 ( .A1(n551), .A2(n561), .ZN(n520) );
  XNOR2_X1 U602 ( .A(KEYINPUT91), .B(KEYINPUT33), .ZN(n519) );
  XNOR2_X1 U603 ( .A(KEYINPUT93), .B(G898), .ZN(n701) );
  NAND2_X1 U604 ( .A1(n701), .A2(G953), .ZN(n521) );
  XNOR2_X1 U605 ( .A(n521), .B(KEYINPUT94), .ZN(n696) );
  OR2_X1 U606 ( .A1(n522), .A2(n696), .ZN(n524) );
  NAND2_X1 U607 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U608 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U609 ( .A(KEYINPUT90), .B(KEYINPUT0), .ZN(n527) );
  XNOR2_X1 U610 ( .A(n528), .B(n527), .ZN(n535) );
  BUF_X1 U611 ( .A(n535), .Z(n556) );
  XNOR2_X1 U612 ( .A(KEYINPUT79), .B(KEYINPUT34), .ZN(n529) );
  XNOR2_X1 U613 ( .A(n529), .B(KEYINPUT73), .ZN(n530) );
  XNOR2_X1 U614 ( .A(n531), .B(n530), .ZN(n533) );
  NAND2_X1 U615 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U616 ( .A(n534), .B(KEYINPUT35), .ZN(n648) );
  INV_X1 U617 ( .A(n535), .ZN(n537) );
  NAND2_X1 U618 ( .A1(n537), .A2(n349), .ZN(n539) );
  XNOR2_X1 U619 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n538) );
  XNOR2_X1 U620 ( .A(n539), .B(n538), .ZN(n547) );
  OR2_X2 U621 ( .A1(n547), .A2(n542), .ZN(n562) );
  NOR2_X2 U622 ( .A1(n562), .A2(n460), .ZN(n540) );
  XNOR2_X1 U623 ( .A(n540), .B(KEYINPUT64), .ZN(n541) );
  NAND2_X1 U624 ( .A1(n541), .A2(n564), .ZN(n645) );
  NAND2_X1 U625 ( .A1(n542), .A2(n564), .ZN(n543) );
  XOR2_X1 U626 ( .A(KEYINPUT110), .B(n543), .Z(n545) );
  INV_X1 U627 ( .A(n561), .ZN(n544) );
  NAND2_X1 U628 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U629 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U630 ( .A(KEYINPUT32), .B(n548), .Z(n721) );
  NAND2_X1 U631 ( .A1(n645), .A2(n721), .ZN(n549) );
  XNOR2_X1 U632 ( .A(n550), .B(KEYINPUT44), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n551), .A2(n460), .ZN(n607) );
  NOR2_X1 U634 ( .A1(n607), .A2(n556), .ZN(n552) );
  XNOR2_X1 U635 ( .A(n552), .B(KEYINPUT31), .ZN(n678) );
  NOR2_X1 U636 ( .A1(n460), .A2(n602), .ZN(n553) );
  NAND2_X1 U637 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U639 ( .A(KEYINPUT100), .B(n557), .Z(n670) );
  NAND2_X1 U640 ( .A1(n678), .A2(n670), .ZN(n558) );
  XNOR2_X1 U641 ( .A(n558), .B(KEYINPUT101), .ZN(n560) );
  NOR2_X1 U642 ( .A1(n560), .A2(n559), .ZN(n566) );
  NOR2_X1 U643 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U644 ( .A(KEYINPUT88), .B(n563), .Z(n565) );
  NOR2_X1 U645 ( .A1(n565), .A2(n564), .ZN(n666) );
  NOR2_X1 U646 ( .A1(n566), .A2(n666), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n568), .A2(n567), .ZN(n570) );
  NOR2_X1 U648 ( .A1(n571), .A2(n698), .ZN(n593) );
  NOR2_X1 U649 ( .A1(n593), .A2(n572), .ZN(n577) );
  INV_X1 U650 ( .A(n698), .ZN(n574) );
  NAND2_X1 U651 ( .A1(n574), .A2(n573), .ZN(n592) );
  INV_X1 U652 ( .A(KEYINPUT2), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n592), .A2(n575), .ZN(n576) );
  NAND2_X1 U654 ( .A1(n577), .A2(n576), .ZN(n650) );
  INV_X2 U655 ( .A(n650), .ZN(n690) );
  NAND2_X1 U656 ( .A1(n690), .A2(G469), .ZN(n581) );
  XNOR2_X1 U657 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n578) );
  XNOR2_X1 U658 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U659 ( .A(n581), .B(n580), .ZN(n583) );
  INV_X1 U660 ( .A(G952), .ZN(n582) );
  AND2_X1 U661 ( .A1(n582), .A2(G953), .ZN(n694) );
  NAND2_X1 U662 ( .A1(n690), .A2(G472), .ZN(n588) );
  XOR2_X1 U663 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  NAND2_X1 U664 ( .A1(n350), .A2(n589), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n590), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U666 ( .A(KEYINPUT2), .B(KEYINPUT81), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT85), .ZN(n632) );
  INV_X1 U668 ( .A(n622), .ZN(n596) );
  AND2_X1 U669 ( .A1(n596), .A2(n610), .ZN(n630) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U671 ( .A(KEYINPUT49), .B(n599), .Z(n600) );
  NOR2_X1 U672 ( .A1(n600), .A2(n460), .ZN(n601) );
  XOR2_X1 U673 ( .A(KEYINPUT119), .B(n601), .Z(n606) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT50), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n609), .B(KEYINPUT51), .ZN(n612) );
  INV_X1 U679 ( .A(n610), .ZN(n611) );
  NOR2_X1 U680 ( .A1(n612), .A2(n611), .ZN(n625) );
  NAND2_X1 U681 ( .A1(n613), .A2(n616), .ZN(n615) );
  NOR2_X1 U682 ( .A1(n615), .A2(n614), .ZN(n621) );
  NOR2_X1 U683 ( .A1(n617), .A2(n616), .ZN(n619) );
  NOR2_X1 U684 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U685 ( .A1(n621), .A2(n620), .ZN(n623) );
  NOR2_X1 U686 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U687 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U688 ( .A(n626), .B(KEYINPUT52), .ZN(n627) );
  NOR2_X1 U689 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U690 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U691 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U692 ( .A1(n635), .A2(n405), .ZN(n637) );
  INV_X1 U693 ( .A(KEYINPUT53), .ZN(n636) );
  XNOR2_X1 U694 ( .A(n637), .B(n636), .ZN(G75) );
  INV_X1 U695 ( .A(n638), .ZN(n641) );
  NAND2_X1 U696 ( .A1(n641), .A2(n639), .ZN(n640) );
  XNOR2_X1 U697 ( .A(n640), .B(G146), .ZN(G48) );
  NAND2_X1 U698 ( .A1(n641), .A2(n669), .ZN(n643) );
  XOR2_X1 U699 ( .A(G128), .B(KEYINPUT29), .Z(n642) );
  XNOR2_X1 U700 ( .A(n643), .B(n642), .ZN(G30) );
  XNOR2_X1 U701 ( .A(n644), .B(G137), .ZN(G39) );
  BUF_X1 U702 ( .A(n645), .Z(n646) );
  XNOR2_X1 U703 ( .A(n646), .B(G110), .ZN(G12) );
  XNOR2_X1 U704 ( .A(n647), .B(G143), .ZN(G45) );
  XOR2_X1 U705 ( .A(n648), .B(G122), .Z(G24) );
  XNOR2_X1 U706 ( .A(n649), .B(G131), .ZN(G33) );
  NOR2_X1 U707 ( .A1(n650), .A2(n651), .ZN(n654) );
  XNOR2_X1 U708 ( .A(n652), .B(KEYINPUT59), .ZN(n653) );
  XNOR2_X1 U709 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U710 ( .A1(n655), .A2(n694), .ZN(n657) );
  XNOR2_X1 U711 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n656) );
  XNOR2_X1 U712 ( .A(n657), .B(n656), .ZN(G60) );
  NAND2_X1 U713 ( .A1(n690), .A2(G210), .ZN(n662) );
  XOR2_X1 U714 ( .A(KEYINPUT89), .B(KEYINPUT54), .Z(n659) );
  XNOR2_X1 U715 ( .A(n659), .B(KEYINPUT55), .ZN(n660) );
  XNOR2_X1 U716 ( .A(n658), .B(n660), .ZN(n661) );
  XNOR2_X1 U717 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X1 U718 ( .A1(n663), .A2(n694), .ZN(n665) );
  XOR2_X1 U719 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n664) );
  XNOR2_X1 U720 ( .A(n665), .B(n664), .ZN(G51) );
  XOR2_X1 U721 ( .A(G101), .B(n666), .Z(G3) );
  NOR2_X1 U722 ( .A1(n670), .A2(n676), .ZN(n668) );
  XNOR2_X1 U723 ( .A(G104), .B(KEYINPUT115), .ZN(n667) );
  XNOR2_X1 U724 ( .A(n668), .B(n667), .ZN(G6) );
  INV_X1 U725 ( .A(n669), .ZN(n679) );
  NOR2_X1 U726 ( .A1(n670), .A2(n679), .ZN(n675) );
  XOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n672) );
  XNOR2_X1 U728 ( .A(G107), .B(KEYINPUT116), .ZN(n671) );
  XNOR2_X1 U729 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U730 ( .A(KEYINPUT26), .B(n673), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n675), .B(n674), .ZN(G9) );
  NOR2_X1 U732 ( .A1(n676), .A2(n678), .ZN(n677) );
  XOR2_X1 U733 ( .A(G113), .B(n677), .Z(G15) );
  NOR2_X1 U734 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U735 ( .A(G116), .B(n680), .Z(G18) );
  XOR2_X1 U736 ( .A(G125), .B(n681), .Z(n682) );
  XNOR2_X1 U737 ( .A(n682), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U738 ( .A(n683), .B(G134), .ZN(n684) );
  XNOR2_X1 U739 ( .A(KEYINPUT118), .B(n684), .ZN(G36) );
  NAND2_X1 U740 ( .A1(n690), .A2(G478), .ZN(n686) );
  XOR2_X1 U741 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n685) );
  XNOR2_X1 U742 ( .A(n686), .B(n685), .ZN(n688) );
  XNOR2_X1 U743 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U744 ( .A1(n694), .A2(n689), .ZN(G63) );
  NAND2_X1 U745 ( .A1(n690), .A2(G217), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U747 ( .A1(n694), .A2(n693), .ZN(G66) );
  XNOR2_X1 U748 ( .A(n695), .B(G101), .ZN(n697) );
  NAND2_X1 U749 ( .A1(n697), .A2(n696), .ZN(n706) );
  NOR2_X1 U750 ( .A1(n698), .A2(G953), .ZN(n704) );
  NAND2_X1 U751 ( .A1(G953), .A2(G224), .ZN(n699) );
  XOR2_X1 U752 ( .A(KEYINPUT61), .B(n699), .Z(n700) );
  NOR2_X1 U753 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U754 ( .A(n702), .B(KEYINPUT124), .ZN(n703) );
  NOR2_X1 U755 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n706), .B(n705), .ZN(G69) );
  XNOR2_X1 U757 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U758 ( .A(n709), .B(KEYINPUT125), .ZN(n710) );
  XNOR2_X1 U759 ( .A(n711), .B(n710), .ZN(n715) );
  XNOR2_X1 U760 ( .A(n715), .B(KEYINPUT126), .ZN(n712) );
  XNOR2_X1 U761 ( .A(n573), .B(n712), .ZN(n713) );
  NOR2_X1 U762 ( .A1(G953), .A2(n713), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n714), .B(KEYINPUT127), .ZN(n719) );
  XNOR2_X1 U764 ( .A(G227), .B(n715), .ZN(n716) );
  NAND2_X1 U765 ( .A1(n716), .A2(G900), .ZN(n717) );
  NAND2_X1 U766 ( .A1(G953), .A2(n717), .ZN(n718) );
  NAND2_X1 U767 ( .A1(n719), .A2(n718), .ZN(G72) );
  XNOR2_X1 U768 ( .A(G140), .B(n720), .ZN(G42) );
  XNOR2_X1 U769 ( .A(G119), .B(n721), .ZN(G21) );
endmodule

