//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT67), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT69), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  OR4_X1    g028(.A1(G221), .A2(G220), .A3(G219), .A4(G218), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n465), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(new_n468), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  XOR2_X1   g058(.A(KEYINPUT3), .B(G2104), .Z(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n465), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n483), .B1(new_n485), .B2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n484), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n465), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n468), .B2(new_n490), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n467), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n495), .A2(new_n465), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT72), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT72), .A2(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XOR2_X1   g078(.A(new_n503), .B(KEYINPUT74), .Z(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT72), .B(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT5), .B(G543), .Z(new_n510));
  NOR2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(G88), .ZN(new_n512));
  AOI22_X1  g087(.A1(G50), .A2(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  OAI21_X1  g090(.A(KEYINPUT76), .B1(new_n507), .B2(new_n508), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT72), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT72), .A2(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT6), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n505), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT75), .B1(new_n510), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n499), .A2(new_n528), .A3(G63), .A4(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n521), .A2(G89), .A3(new_n499), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n525), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n516), .B2(new_n523), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n510), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(new_n506), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n521), .A2(G90), .A3(new_n499), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g118(.A1(new_n537), .A2(new_n543), .A3(KEYINPUT77), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n541), .A2(new_n542), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n522), .B1(new_n521), .B2(G543), .ZN(new_n547));
  AOI211_X1 g122(.A(KEYINPUT76), .B(new_n508), .C1(new_n519), .C2(new_n520), .ZN(new_n548));
  OAI21_X1  g123(.A(G52), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n545), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n544), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n510), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n511), .A2(G81), .B1(new_n555), .B2(new_n506), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n516), .B2(new_n523), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n501), .B2(new_n502), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n567), .C2(new_n505), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT78), .B1(new_n507), .B2(new_n510), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n521), .A2(new_n571), .A3(new_n499), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(G91), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(G78), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n499), .B2(G65), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  INV_X1    g151(.A(G651), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n575), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n569), .A2(new_n573), .A3(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n525), .A2(new_n534), .ZN(G286));
  NAND3_X1  g157(.A1(new_n570), .A2(G87), .A3(new_n572), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n570), .A2(KEYINPUT80), .A3(G87), .A4(new_n572), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n521), .A2(G49), .A3(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n510), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n509), .A2(G48), .B1(new_n595), .B2(new_n506), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n570), .A2(G86), .A3(new_n572), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n524), .A2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n510), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n511), .A2(G85), .B1(new_n602), .B2(new_n506), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G290));
  NAND3_X1  g179(.A1(new_n570), .A2(G92), .A3(new_n572), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n570), .A2(KEYINPUT10), .A3(G92), .A4(new_n572), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n510), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n524), .A2(G54), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n614), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g190(.A(new_n614), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(new_n614), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n479), .A2(G135), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n485), .B2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n633), .A2(G2096), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n634), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(new_n658), .A3(G14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(KEYINPUT17), .ZN(new_n667));
  INV_X1    g242(.A(new_n661), .ZN(new_n668));
  INV_X1    g243(.A(new_n662), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n664), .A3(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n663), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n666), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  AOI211_X1 g259(.A(new_n682), .B(new_n684), .C1(new_n677), .C2(new_n681), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT84), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  NAND3_X1  g267(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n696));
  INV_X1    g271(.A(G139), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n695), .B1(new_n465), .B2(new_n696), .C1(new_n478), .C2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G33), .B(new_n698), .S(G29), .Z(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G2072), .Z(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n701), .A2(G32), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n479), .A2(G141), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n485), .A2(G129), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT26), .Z(new_n707));
  NAND4_X1  g282(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n702), .B1(new_n708), .B2(G29), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n701), .B1(new_n711), .B2(G34), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G34), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G160), .B2(G29), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n709), .A2(new_n710), .B1(G2084), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n700), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n701), .A2(G35), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT95), .Z(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n487), .B2(G29), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT97), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2090), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n701), .A2(G26), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT28), .Z(new_n726));
  OR2_X1    g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT89), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G128), .B2(new_n485), .ZN(new_n730));
  INV_X1    g305(.A(G140), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n478), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2067), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G19), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n560), .B2(G16), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1341), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(G1341), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n701), .A2(G27), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G164), .B2(new_n701), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n734), .A2(new_n737), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G4), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n621), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT88), .B(G1348), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n717), .A2(new_n724), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G5), .A2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  INV_X1    g325(.A(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(G301), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n754), .B1(G2084), .B2(new_n714), .C1(new_n709), .C2(new_n710), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n751), .A2(G20), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT23), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n618), .B2(new_n751), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT98), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n755), .A2(KEYINPUT94), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n756), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n751), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n751), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT91), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1966), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n752), .A2(new_n753), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n628), .A2(G29), .A3(new_n632), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT30), .B(G28), .ZN(new_n771));
  OR2_X1    g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NAND2_X1  g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n771), .A2(new_n701), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n748), .A2(new_n764), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G16), .A2(G23), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT85), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n587), .B2(new_n591), .ZN(new_n783));
  AOI211_X1 g358(.A(KEYINPUT86), .B(new_n590), .C1(new_n585), .C2(new_n586), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n781), .B1(new_n785), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT87), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT33), .B(G1976), .Z(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n751), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n751), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1971), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n751), .A2(G6), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G305), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT32), .B(G1981), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n795), .A2(new_n797), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n793), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n789), .A2(new_n790), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n485), .A2(G119), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n465), .A2(G107), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G131), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n804), .B1(new_n805), .B2(new_n806), .C1(new_n478), .C2(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G25), .B(new_n808), .S(G29), .Z(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1986), .ZN(new_n812));
  INV_X1    g387(.A(G290), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n751), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n751), .B2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n811), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n812), .B2(new_n815), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n802), .A2(new_n803), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(KEYINPUT36), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(KEYINPUT36), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n779), .B1(new_n820), .B2(new_n821), .ZN(G311));
  AND3_X1   g397(.A1(new_n748), .A2(new_n777), .A3(new_n778), .ZN(new_n823));
  INV_X1    g398(.A(new_n821), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n823), .B(new_n764), .C1(new_n824), .C2(new_n819), .ZN(G150));
  NOR2_X1   g400(.A1(new_n614), .A2(new_n622), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  INV_X1    g402(.A(new_n559), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n524), .A2(G55), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  INV_X1    g405(.A(new_n506), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n521), .A2(G93), .A3(new_n499), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n828), .A2(new_n829), .A3(new_n834), .A4(new_n556), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n516), .B2(new_n523), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n832), .A2(new_n833), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n557), .A2(new_n559), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n827), .B(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n842), .A2(new_n843), .A3(G860), .ZN(new_n844));
  OAI21_X1  g419(.A(G860), .B1(new_n837), .B2(new_n838), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n485), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n465), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  INV_X1    g425(.A(G142), .ZN(new_n851));
  OAI221_X1 g426(.A(new_n848), .B1(new_n849), .B2(new_n850), .C1(new_n478), .C2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n636), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n708), .B(new_n698), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n732), .B(new_n497), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n808), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(G160), .B(KEYINPUT99), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n487), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n633), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g441(.A(G303), .B(G305), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(G288), .A2(KEYINPUT86), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n587), .A2(new_n782), .A3(new_n591), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n813), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(G290), .B1(new_n783), .B2(new_n784), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT102), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n867), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n609), .A2(G299), .A3(new_n613), .ZN(new_n881));
  AOI21_X1  g456(.A(G299), .B1(new_n609), .B2(new_n613), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n614), .A2(new_n618), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n609), .A2(G299), .A3(new_n613), .ZN(new_n885));
  XOR2_X1   g460(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n885), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n624), .B(new_n840), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n889), .B(new_n890), .S(new_n891), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n879), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n879), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n837), .A2(new_n838), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(G868), .B2(new_n897), .ZN(G295));
  OAI21_X1  g473(.A(new_n896), .B1(G868), .B2(new_n897), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT77), .B1(new_n537), .B2(new_n543), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n546), .A2(new_n549), .A3(new_n545), .ZN(new_n902));
  AND3_X1   g477(.A1(G286), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G286), .B1(new_n902), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n840), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(G168), .B1(new_n544), .B2(new_n550), .ZN(new_n906));
  NAND3_X1  g481(.A1(G286), .A2(new_n901), .A3(new_n902), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n839), .A3(new_n835), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n908), .A3(new_n890), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n905), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n889), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n905), .A2(new_n908), .A3(new_n890), .A4(KEYINPUT103), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n878), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n887), .B1(new_n881), .B2(new_n882), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n884), .A2(new_n880), .A3(new_n885), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n905), .A2(new_n908), .A3(new_n890), .A4(KEYINPUT105), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n875), .A3(new_n877), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n916), .A2(new_n917), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n917), .B1(new_n916), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n910), .A2(new_n909), .B1(new_n889), .B2(new_n912), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n813), .B1(new_n869), .B2(new_n870), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n783), .A2(new_n784), .A3(G290), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n867), .B1(new_n933), .B2(new_n876), .ZN(new_n934));
  INV_X1    g509(.A(new_n877), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n914), .B(new_n929), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n875), .A3(new_n877), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n900), .B1(new_n928), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n936), .A2(new_n925), .A3(new_n937), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n944), .A2(KEYINPUT104), .B1(new_n945), .B2(new_n941), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n916), .B2(new_n939), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT44), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT107), .B1(new_n943), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n916), .A2(new_n925), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n916), .A2(new_n917), .A3(new_n925), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n941), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n942), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n947), .A2(new_n948), .B1(new_n952), .B2(KEYINPUT43), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n944), .A2(KEYINPUT104), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n900), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n951), .A2(new_n962), .ZN(G397));
  AND2_X1   g538(.A1(G160), .A2(G40), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G160), .A2(G40), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n497), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(G1996), .A3(new_n708), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT110), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n732), .B(G2067), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n708), .A2(G1996), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n810), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n808), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n808), .A2(new_n981), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n974), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(KEYINPUT127), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n974), .A2(new_n812), .A3(new_n813), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT125), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n732), .A2(G2067), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n980), .B2(new_n982), .ZN(new_n994));
  INV_X1    g569(.A(new_n974), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n994), .A2(new_n992), .A3(new_n995), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(G1996), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT46), .Z(new_n1000));
  OAI21_X1  g575(.A(new_n974), .B1(new_n977), .B2(new_n708), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT126), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT47), .Z(new_n1004));
  NOR3_X1   g579(.A1(new_n997), .A2(new_n998), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n971), .A2(new_n966), .A3(new_n968), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT113), .B(G86), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n511), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n596), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G1981), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(G305), .B2(G1981), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1007), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1007), .A2(new_n1014), .A3(KEYINPUT114), .A4(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G288), .A2(G1976), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(G1981), .B2(G305), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n785), .A2(G1976), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1007), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1976), .B1(new_n587), .B2(new_n591), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n1025), .A2(KEYINPUT52), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1027), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT55), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2090), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n497), .A2(new_n970), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n966), .B(new_n968), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n971), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n973), .B1(new_n497), .B2(new_n970), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(KEYINPUT45), .B2(new_n971), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n966), .A2(new_n968), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1971), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1034), .A2(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1033), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1023), .A2(new_n1007), .B1(new_n1029), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1035), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n497), .A2(new_n970), .A3(new_n973), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n968), .A4(new_n966), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT116), .B(G2084), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1038), .A2(new_n1040), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G168), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(new_n1048), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1051), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1031), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1027), .A2(new_n1020), .A3(new_n1028), .A4(new_n1072), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1073), .A2(KEYINPUT117), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(KEYINPUT117), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1071), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT63), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1053), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G286), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1079));
  AOI211_X1 g654(.A(G168), .B(new_n1066), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT51), .B(G8), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1063), .A2(G168), .A3(new_n1067), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1085), .A3(KEYINPUT62), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT124), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1081), .A2(new_n1085), .A3(new_n1088), .A4(KEYINPUT62), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n1090));
  NAND2_X1  g665(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1063), .A2(G286), .A3(new_n1067), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1069), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT51), .B1(new_n1082), .B2(G8), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1090), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1043), .A2(new_n1044), .A3(new_n741), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1096), .A2(new_n753), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OR3_X1    g674(.A1(new_n1057), .A2(new_n1098), .A3(G2078), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(G301), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1087), .A2(new_n1089), .A3(new_n1095), .A4(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1036), .B1(new_n497), .B2(new_n970), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n969), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT118), .B1(new_n1106), .B2(G1956), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1104), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1105), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1044), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1043), .A2(new_n1044), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT121), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1043), .A2(new_n1044), .A3(new_n1117), .A4(new_n1114), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1107), .A2(new_n1113), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n580), .A2(new_n573), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT120), .Z(new_n1121));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n569), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n569), .A2(new_n1122), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1123), .A2(new_n1124), .A3(KEYINPUT57), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1121), .A2(new_n1125), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1006), .A2(G2067), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n614), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT61), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1136));
  AND4_X1   g711(.A1(KEYINPUT61), .A2(new_n1135), .A3(new_n1126), .A4(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1006), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT122), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1006), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1141), .B(new_n1143), .C1(G1996), .C2(new_n1045), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n560), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1130), .A2(new_n1131), .A3(new_n614), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT60), .B1(new_n1148), .B2(new_n1132), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n614), .A2(KEYINPUT60), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1130), .A2(new_n1131), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1144), .A2(KEYINPUT59), .A3(new_n560), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1133), .B1(new_n1138), .B2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(G301), .B(KEYINPUT54), .Z(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT123), .B(G2078), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1043), .A2(KEYINPUT53), .A3(new_n964), .A4(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1099), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1101), .B2(new_n1155), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1093), .A2(new_n1159), .A3(new_n1094), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1154), .A2(new_n1160), .B1(new_n1077), .B2(new_n1070), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1103), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1106), .A2(new_n1034), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1031), .B1(new_n1165), .B2(new_n1048), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1029), .A2(new_n1166), .A3(new_n1051), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1078), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(G290), .B(new_n812), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n980), .B(new_n984), .C1(new_n995), .C2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1005), .B1(new_n1168), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g746(.A1(G229), .A2(new_n463), .A3(new_n659), .A4(G227), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n949), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n865), .A3(new_n1174), .ZN(G225));
  INV_X1    g749(.A(G225), .ZN(G308));
endmodule


