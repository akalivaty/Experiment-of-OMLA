//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G214), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(G237), .A2(G953), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(G143), .A3(G214), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT18), .A2(G131), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n196), .A2(new_n197), .ZN(new_n205));
  AOI21_X1  g019(.A(G143), .B1(new_n199), .B2(G214), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT18), .B(G131), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT84), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT84), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n198), .B2(new_n200), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n211), .B2(KEYINPUT18), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n193), .B(new_n204), .C1(new_n208), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT85), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(KEYINPUT84), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n209), .A3(KEYINPUT18), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT85), .A3(new_n193), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n221));
  INV_X1    g035(.A(G140), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G125), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n223), .A2(KEYINPUT16), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n221), .A2(G146), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(G146), .B1(new_n221), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G131), .B1(new_n205), .B2(new_n206), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n198), .A2(new_n210), .A3(new_n200), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n211), .A2(KEYINPUT17), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n227), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n190), .B1(new_n220), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n190), .ZN(new_n236));
  AOI211_X1 g050(.A(new_n236), .B(new_n233), .C1(new_n215), .C2(new_n219), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n187), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G475), .ZN(new_n239));
  NOR2_X1   g053(.A1(G475), .A2(G902), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT89), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G125), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G140), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n222), .A2(G125), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT19), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(G140), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT19), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n223), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n192), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT87), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n221), .A2(G146), .A3(new_n224), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n246), .A2(new_n253), .A3(new_n192), .A4(new_n249), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT88), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n251), .A2(KEYINPUT88), .A3(new_n252), .A4(new_n254), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT86), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n228), .A2(new_n259), .A3(new_n230), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n228), .B2(new_n230), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n213), .A2(new_n214), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT85), .B1(new_n218), .B2(new_n193), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n236), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n220), .A2(new_n190), .A3(new_n234), .ZN(new_n268));
  AOI211_X1 g082(.A(KEYINPUT20), .B(new_n242), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n190), .B1(new_n220), .B2(new_n263), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n241), .B1(new_n270), .B2(new_n237), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT20), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT90), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n242), .B1(new_n267), .B2(new_n268), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n239), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT91), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n276), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n267), .A2(new_n268), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n276), .B1(new_n283), .B2(new_n241), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n284), .B2(KEYINPUT90), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n277), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT91), .A3(new_n239), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT9), .B(G234), .Z(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(G217), .A3(new_n195), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n290), .B(KEYINPUT94), .Z(new_n291));
  INV_X1    g105(.A(G128), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G143), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(G143), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(KEYINPUT13), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT92), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT92), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n293), .C1(new_n294), .C2(KEYINPUT13), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G134), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n302), .A2(G122), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(G122), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G107), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n294), .ZN(new_n308));
  INV_X1    g122(.A(G134), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n293), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n301), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n197), .A2(G128), .ZN(new_n312));
  OAI21_X1  g126(.A(G134), .B1(new_n312), .B2(new_n294), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n306), .B1(new_n303), .B2(KEYINPUT14), .ZN(new_n317));
  INV_X1    g131(.A(new_n305), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n310), .A2(KEYINPUT93), .A3(new_n313), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n303), .B(new_n304), .C1(KEYINPUT14), .C2(new_n306), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n316), .A2(new_n319), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n291), .B1(new_n311), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n291), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n301), .A2(new_n307), .A3(new_n310), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(KEYINPUT95), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT95), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n326), .A2(new_n322), .A3(new_n325), .A4(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n330), .A3(new_n187), .ZN(new_n331));
  INV_X1    g145(.A(G478), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(KEYINPUT15), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G214), .B1(G237), .B2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT81), .B(G224), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n195), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT0), .A2(G128), .ZN(new_n339));
  XNOR2_X1  g153(.A(G143), .B(G146), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(KEYINPUT64), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n192), .A2(G143), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n197), .A2(G146), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G128), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT64), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n347), .A3(G125), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n341), .A2(new_n347), .A3(KEYINPUT80), .A4(G125), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n192), .A2(G143), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G128), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n192), .A2(new_n312), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT65), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n292), .A2(KEYINPUT1), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n360), .A2(new_n343), .B1(new_n293), .B2(G146), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT65), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n342), .A3(new_n343), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n359), .A2(new_n243), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n352), .A2(new_n353), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n353), .B1(new_n352), .B2(new_n364), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n338), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n352), .A2(new_n364), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT82), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(new_n195), .A3(new_n337), .A4(new_n365), .ZN(new_n371));
  XNOR2_X1  g185(.A(G116), .B(G119), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT2), .B(G113), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n376));
  INV_X1    g190(.A(G119), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(G116), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT79), .A4(G116), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n380), .A2(G113), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n372), .A2(KEYINPUT5), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n306), .A3(G104), .ZN(new_n387));
  INV_X1    g201(.A(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n189), .A2(G107), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n385), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n306), .A2(G104), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n189), .A2(G107), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n372), .B(new_n374), .Z(new_n397));
  NAND3_X1  g211(.A1(new_n385), .A2(new_n387), .A3(new_n389), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G101), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(G101), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n405));
  XOR2_X1   g219(.A(G110), .B(G122), .Z(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n406), .ZN(new_n408));
  INV_X1    g222(.A(new_n406), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n368), .A2(new_n371), .A3(new_n407), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n338), .A2(KEYINPUT7), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n369), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n384), .A2(new_n394), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n406), .B(KEYINPUT8), .Z(new_n416));
  XOR2_X1   g230(.A(new_n383), .B(KEYINPUT83), .Z(new_n417));
  AOI21_X1  g231(.A(new_n375), .B1(new_n417), .B2(new_n382), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n415), .B(new_n416), .C1(new_n418), .C2(new_n394), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n364), .A2(new_n348), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n413), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n414), .A2(new_n419), .A3(new_n421), .A4(new_n410), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n412), .A2(new_n187), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G210), .B1(G237), .B2(G902), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n412), .A2(new_n187), .A3(new_n424), .A4(new_n422), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n336), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(G234), .A2(G237), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G952), .A3(new_n195), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT21), .B(G898), .Z(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(G902), .A3(G953), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n288), .A2(new_n334), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT22), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(G137), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT24), .B(G110), .Z(new_n440));
  XNOR2_X1  g254(.A(G119), .B(G128), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT23), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n377), .B2(G128), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n292), .A2(KEYINPUT23), .A3(G119), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n445), .C1(G119), .C2(new_n292), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n442), .A2(KEYINPUT71), .B1(new_n446), .B2(G110), .ZN(new_n447));
  OAI221_X1 g261(.A(new_n447), .B1(KEYINPUT71), .B2(new_n442), .C1(new_n225), .C2(new_n226), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n446), .A2(G110), .B1(new_n441), .B2(new_n440), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n191), .A2(new_n192), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n252), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n448), .A2(KEYINPUT72), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT72), .B1(new_n448), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n439), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n448), .A2(new_n451), .A3(new_n438), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n187), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G217), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(G234), .B2(new_n187), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT25), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n462), .A2(G902), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n465), .B(KEYINPUT74), .Z(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n454), .A2(new_n467), .A3(new_n455), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(G472), .A2(G902), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n199), .A2(G210), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT27), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT26), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT26), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n474), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n388), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT68), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT68), .B1(new_n476), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n309), .A2(G137), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n309), .A2(G137), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT11), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n309), .B2(G137), .ZN(new_n490));
  INV_X1    g304(.A(G137), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT11), .A3(G134), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n490), .A2(new_n492), .A3(new_n210), .A4(new_n485), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n397), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n485), .A3(new_n492), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G131), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n493), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT66), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(KEYINPUT66), .A3(new_n493), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n341), .A2(new_n347), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT67), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n501), .A2(new_n506), .A3(new_n502), .A4(new_n503), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n496), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n499), .A2(new_n503), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n495), .B1(new_n494), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n483), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n495), .A3(new_n494), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n482), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n476), .A2(new_n479), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n494), .A2(new_n517), .A3(new_n509), .ZN(new_n518));
  INV_X1    g332(.A(new_n494), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n505), .B2(new_n507), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n518), .B1(new_n520), .B2(new_n517), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n508), .B(new_n516), .C1(new_n521), .C2(new_n397), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n515), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n397), .ZN(new_n525));
  INV_X1    g339(.A(new_n508), .ZN(new_n526));
  INV_X1    g340(.A(new_n516), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT31), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n471), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n511), .A2(new_n482), .A3(new_n514), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n508), .B1(new_n521), .B2(new_n397), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n527), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n526), .B1(new_n495), .B2(new_n520), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT28), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n512), .A2(KEYINPUT70), .A3(new_n513), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n514), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n516), .A2(new_n532), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n541), .A3(new_n187), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n530), .A2(KEYINPUT32), .B1(G472), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n525), .A2(new_n523), .A3(new_n526), .A4(new_n527), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n511), .A2(new_n514), .ZN(new_n545));
  INV_X1    g359(.A(new_n482), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n523), .B1(new_n533), .B2(new_n527), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n470), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT32), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n469), .B1(new_n543), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT76), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n363), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n340), .A2(KEYINPUT76), .A3(new_n360), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n357), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n395), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT10), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n484), .A2(KEYINPUT10), .A3(new_n395), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n501), .A2(new_n502), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n402), .A2(new_n503), .A3(new_n400), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n562), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n359), .A2(new_n394), .A3(new_n362), .A4(new_n363), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n558), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT12), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n567), .A2(KEYINPUT12), .A3(new_n499), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT77), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G140), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n195), .A2(G227), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n576), .B(new_n564), .C1(new_n568), .C2(new_n569), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n564), .A2(new_n574), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT78), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n565), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n564), .A2(KEYINPUT78), .A3(new_n574), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n578), .A2(G469), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(G469), .A2(G902), .ZN(new_n587));
  INV_X1    g401(.A(G469), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n568), .A2(new_n569), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n579), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n574), .B1(new_n583), .B2(new_n564), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n588), .B(new_n187), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n289), .A2(new_n187), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G221), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT75), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n435), .A2(new_n553), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  INV_X1    g413(.A(new_n434), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n328), .A2(new_n330), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n328), .A2(new_n330), .A3(KEYINPUT96), .A4(new_n601), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n324), .A2(KEYINPUT33), .A3(new_n327), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n606), .A2(G478), .A3(new_n187), .A4(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n331), .A2(new_n332), .ZN(new_n611));
  INV_X1    g425(.A(new_n607), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n604), .B2(new_n605), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n613), .A2(KEYINPUT97), .A3(G478), .A4(new_n187), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT91), .B1(new_n286), .B2(new_n239), .ZN(new_n616));
  INV_X1    g430(.A(new_n239), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n280), .B(new_n617), .C1(new_n285), .C2(new_n277), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n600), .B(new_n615), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n529), .A2(new_n544), .A3(new_n547), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n187), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n593), .A2(new_n596), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n623), .A2(new_n530), .A3(new_n624), .A4(new_n469), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT98), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT34), .ZN(G6));
  NAND2_X1  g443(.A1(new_n282), .A2(new_n272), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n334), .A3(new_n239), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n434), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n623), .A2(new_n530), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n452), .A2(new_n453), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n439), .A2(KEYINPUT36), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n637), .B(new_n638), .Z(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n467), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n464), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n435), .A2(new_n597), .A3(new_n636), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT37), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G110), .ZN(G12));
  NAND3_X1  g458(.A1(new_n622), .A2(KEYINPUT32), .A3(new_n470), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n542), .A2(G472), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n552), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n426), .A2(new_n427), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n335), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n432), .A2(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n430), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n238), .B2(G475), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n630), .A2(new_n334), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n648), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n647), .A2(new_n597), .A3(new_n641), .A4(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n650), .A2(new_n655), .A3(new_n648), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n292), .ZN(G30));
  INV_X1    g474(.A(new_n334), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n281), .B2(new_n287), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n649), .B(KEYINPUT38), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n335), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n533), .A2(new_n527), .B1(new_n546), .B2(new_n535), .ZN(new_n666));
  OAI211_X1 g480(.A(KEYINPUT100), .B(G472), .C1(new_n666), .C2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n645), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n666), .A2(G472), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND2_X1  g486(.A1(G472), .A2(G902), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n669), .A2(new_n670), .A3(new_n552), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n552), .A2(new_n674), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT101), .B1(new_n676), .B2(new_n668), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n641), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n665), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n665), .A2(new_n678), .A3(KEYINPUT102), .A4(new_n679), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n652), .B(KEYINPUT39), .Z(new_n684));
  NOR2_X1   g498(.A1(new_n624), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n682), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT103), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n197), .ZN(G45));
  NAND4_X1  g505(.A1(new_n647), .A2(new_n597), .A3(new_n428), .A4(new_n641), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n615), .B(new_n652), .C1(new_n616), .C2(new_n618), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n192), .ZN(G48));
  NOR2_X1   g509(.A1(new_n590), .A2(new_n591), .ZN(new_n696));
  OAI21_X1  g510(.A(G469), .B1(new_n696), .B2(G902), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n596), .A3(new_n592), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n697), .A2(KEYINPUT104), .A3(new_n596), .A4(new_n592), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n620), .A2(new_n553), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n553), .A2(new_n706), .A3(new_n632), .A4(new_n702), .ZN(new_n707));
  INV_X1    g521(.A(new_n469), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n647), .A2(new_n632), .A3(new_n708), .A4(new_n702), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT105), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NOR2_X1   g526(.A1(new_n288), .A2(new_n334), .ZN(new_n713));
  INV_X1    g527(.A(new_n698), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n428), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT106), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n679), .B1(new_n543), .B2(new_n552), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n713), .A2(new_n716), .A3(new_n433), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NAND2_X1  g533(.A1(new_n505), .A2(new_n507), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n494), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n508), .B1(new_n721), .B2(new_n397), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n537), .B(new_n539), .C1(new_n722), .C2(new_n513), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n546), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n529), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT107), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n529), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n544), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n623), .B1(new_n729), .B2(new_n470), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n434), .B1(new_n700), .B2(new_n701), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n662), .A2(new_n730), .A3(new_n708), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n641), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n693), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n288), .A2(KEYINPUT108), .A3(new_n615), .A4(new_n652), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n716), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  NAND2_X1  g554(.A1(new_n736), .A2(new_n737), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT109), .B1(new_n649), .B2(new_n336), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n426), .A2(new_n743), .A3(new_n335), .A4(new_n427), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n597), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n552), .A2(KEYINPUT110), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n550), .A2(new_n747), .A3(new_n551), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n543), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n708), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n741), .A2(new_n745), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n745), .A2(new_n647), .A3(new_n708), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT42), .B1(new_n736), .B2(new_n737), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n752), .A2(KEYINPUT42), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND2_X1  g571(.A1(new_n655), .A2(KEYINPUT111), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n655), .A2(KEYINPUT111), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n309), .ZN(G36));
  NOR2_X1   g576(.A1(new_n616), .A2(new_n618), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT43), .B1(new_n763), .B2(KEYINPUT112), .ZN(new_n764));
  INV_X1    g578(.A(new_n615), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n288), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n763), .B(new_n615), .C1(KEYINPUT112), .C2(KEYINPUT43), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n636), .B(new_n679), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n578), .A2(new_n585), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT45), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(G469), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n587), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(G469), .C1(new_n771), .C2(G902), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n592), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n596), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n684), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n742), .A2(new_n744), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n768), .B2(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  XNOR2_X1  g599(.A(new_n777), .B(KEYINPUT47), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n693), .A2(new_n708), .A3(new_n647), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n222), .ZN(G42));
  NAND3_X1  g603(.A1(new_n708), .A2(new_n596), .A3(new_n335), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n288), .A2(new_n790), .A3(new_n765), .A4(new_n663), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n697), .A2(new_n592), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT49), .Z(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n675), .A3(new_n677), .A4(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n711), .A2(new_n703), .A3(new_n718), .A4(new_n732), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n756), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT118), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n756), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n658), .A2(new_n657), .B1(new_n692), .B2(new_n693), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n763), .A2(new_n661), .A3(new_n650), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n652), .B(KEYINPUT116), .Z(new_n805));
  NOR3_X1   g619(.A1(new_n624), .A2(new_n641), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n678), .A2(new_n804), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AND4_X1   g624(.A1(KEYINPUT52), .A2(new_n739), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n802), .B1(new_n738), .B2(new_n716), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(new_n812), .B2(new_n810), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n761), .ZN(new_n815));
  INV_X1    g629(.A(new_n734), .ZN(new_n816));
  AND4_X1   g630(.A1(KEYINPUT115), .A2(new_n741), .A3(new_n816), .A4(new_n745), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT115), .B1(new_n738), .B2(new_n745), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n619), .A2(KEYINPUT113), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n763), .A2(KEYINPUT114), .A3(new_n334), .A4(new_n600), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n281), .A2(new_n600), .A3(new_n334), .A4(new_n287), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n288), .A2(new_n825), .A3(new_n600), .A4(new_n615), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n820), .A2(new_n821), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n625), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n334), .B1(new_n282), .B2(new_n272), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n717), .A2(new_n654), .A3(new_n745), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n828), .A2(new_n598), .A3(new_n642), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n819), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n814), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n598), .A2(new_n828), .A3(new_n642), .A4(new_n830), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n741), .A2(new_n816), .A3(new_n745), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n738), .A2(KEYINPUT115), .A3(new_n745), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n761), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n836), .A2(new_n841), .A3(new_n756), .A4(new_n796), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n811), .A2(new_n813), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n835), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n833), .A2(new_n834), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n797), .A2(new_n819), .A3(new_n831), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(KEYINPUT53), .A3(new_n814), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n834), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n430), .B1(new_n766), .B2(new_n767), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n730), .A2(new_n708), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n335), .B(new_n663), .C1(KEYINPUT119), .C2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(new_n714), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n781), .A2(new_n714), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n816), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n857), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n678), .A2(new_n469), .A3(new_n859), .A4(new_n430), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n763), .A3(new_n765), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n858), .A2(new_n861), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n851), .A2(new_n853), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(new_n781), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n792), .A2(new_n596), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n786), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n786), .A2(KEYINPUT120), .A3(new_n871), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n869), .A2(new_n872), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n866), .B1(new_n865), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n195), .A2(G952), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n763), .A2(new_n765), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n863), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n851), .A2(new_n751), .A3(new_n860), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n885), .B2(KEYINPUT48), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(KEYINPUT48), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n888), .B2(new_n885), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n877), .A2(new_n879), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n868), .A2(new_n716), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n850), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT122), .Z(new_n894));
  OAI21_X1  g708(.A(new_n794), .B1(new_n892), .B2(new_n894), .ZN(G75));
  AOI21_X1  g709(.A(new_n187), .B1(new_n833), .B2(new_n844), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT56), .B1(new_n896), .B2(G210), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n368), .A2(new_n371), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n411), .A2(new_n407), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n898), .B(new_n899), .Z(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT55), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n897), .A2(new_n902), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n195), .A2(G952), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G51));
  INV_X1    g720(.A(KEYINPUT42), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n750), .B1(new_n736), .B2(new_n737), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(new_n745), .ZN(new_n909));
  AOI211_X1 g723(.A(KEYINPUT42), .B(new_n753), .C1(new_n736), .C2(new_n737), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n909), .A2(new_n795), .A3(KEYINPUT118), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n799), .B1(new_n756), .B2(new_n796), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n836), .B(new_n841), .C1(new_n811), .C2(new_n813), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n835), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT53), .B1(new_n847), .B2(new_n814), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT54), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(KEYINPUT123), .A3(new_n845), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n833), .A2(new_n844), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n587), .B(KEYINPUT57), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n696), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n896), .A2(G469), .A3(new_n771), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n905), .B1(new_n925), .B2(new_n926), .ZN(G54));
  NAND2_X1  g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n896), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n283), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n905), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n846), .B2(new_n849), .ZN(new_n938));
  INV_X1    g752(.A(new_n613), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n905), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n918), .A2(new_n613), .A3(new_n921), .A4(new_n937), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT60), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n919), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n454), .A2(new_n455), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n905), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n919), .A2(new_n639), .A3(new_n944), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n947), .A2(KEYINPUT61), .A3(new_n948), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  AOI21_X1  g768(.A(new_n195), .B1(new_n431), .B2(new_n337), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n828), .A2(new_n598), .A3(new_n642), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n795), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n955), .B1(new_n958), .B2(new_n195), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n899), .B1(G898), .B2(new_n195), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(G69));
  NAND2_X1  g775(.A1(new_n246), .A2(new_n249), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n521), .B(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(G900), .B1(new_n964), .B2(G227), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n195), .B(new_n965), .C1(G227), .C2(new_n964), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n688), .A2(new_n689), .A3(new_n812), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n788), .B1(new_n780), .B2(new_n783), .ZN(new_n970));
  INV_X1    g784(.A(new_n881), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n661), .B2(new_n288), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n972), .A2(new_n553), .A3(new_n685), .A4(new_n781), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(G953), .B1(new_n974), .B2(new_n963), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n778), .A2(new_n751), .A3(new_n804), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n812), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n756), .A2(new_n815), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(KEYINPUT125), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(KEYINPUT125), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n970), .B(new_n977), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(new_n963), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n966), .B1(new_n975), .B2(new_n982), .ZN(G72));
  XOR2_X1   g797(.A(new_n673), .B(KEYINPUT63), .Z(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT126), .Z(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n981), .B2(new_n958), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n533), .B(KEYINPUT127), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n516), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n848), .A2(new_n844), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n533), .A2(new_n527), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n989), .B(new_n984), .C1(new_n522), .C2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n948), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n969), .A2(new_n957), .A3(new_n970), .A4(new_n973), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n987), .B1(new_n993), .B2(new_n985), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n992), .B1(new_n527), .B2(new_n994), .ZN(G57));
endmodule


