

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U548 ( .A(KEYINPUT66), .B(n523), .ZN(n778) );
  NOR2_X1 U549 ( .A1(n851), .A2(n850), .ZN(n866) );
  XNOR2_X1 U550 ( .A(n972), .B(n673), .ZN(n674) );
  INV_X1 U551 ( .A(G290), .ZN(n673) );
  XNOR2_X1 U552 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U553 ( .A(KEYINPUT14), .B(n669), .Z(n513) );
  INV_X1 U554 ( .A(KEYINPUT30), .ZN(n819) );
  XNOR2_X1 U555 ( .A(n819), .B(KEYINPUT97), .ZN(n820) );
  XNOR2_X1 U556 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U557 ( .A(KEYINPUT29), .B(KEYINPUT96), .ZN(n813) );
  BUF_X1 U558 ( .A(n817), .Z(n829) );
  XNOR2_X1 U559 ( .A(n814), .B(n813), .ZN(n815) );
  OR2_X1 U560 ( .A1(n855), .A2(n854), .ZN(n856) );
  INV_X1 U561 ( .A(KEYINPUT84), .ZN(n687) );
  OR2_X1 U562 ( .A1(n779), .A2(G1384), .ZN(n780) );
  XNOR2_X1 U563 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U564 ( .A(G305), .B(G299), .ZN(n692) );
  XNOR2_X1 U565 ( .A(n693), .B(n692), .ZN(n763) );
  NOR2_X2 U566 ( .A1(G2105), .A2(n528), .ZN(n595) );
  AND2_X1 U567 ( .A1(n528), .A2(G2105), .ZN(n601) );
  INV_X1 U568 ( .A(KEYINPUT117), .ZN(n737) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n517), .Z(n680) );
  NOR2_X1 U570 ( .A1(G651), .A2(n636), .ZN(n683) );
  NAND2_X1 U571 ( .A1(n672), .A2(n671), .ZN(n972) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n675) );
  NAND2_X1 U573 ( .A1(n675), .A2(G85), .ZN(n515) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n636) );
  XNOR2_X1 U575 ( .A(KEYINPUT67), .B(G651), .ZN(n516) );
  NOR2_X1 U576 ( .A1(n636), .A2(n516), .ZN(n676) );
  NAND2_X1 U577 ( .A1(G72), .A2(n676), .ZN(n514) );
  NAND2_X1 U578 ( .A1(n515), .A2(n514), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n683), .A2(G47), .ZN(n519) );
  NOR2_X1 U580 ( .A1(G543), .A2(n516), .ZN(n517) );
  NAND2_X1 U581 ( .A1(G60), .A2(n680), .ZN(n518) );
  NAND2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n520) );
  OR2_X1 U583 ( .A1(n521), .A2(n520), .ZN(G290) );
  NOR2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X1 U585 ( .A(KEYINPUT17), .B(n522), .Z(n523) );
  NAND2_X1 U586 ( .A1(n778), .A2(G138), .ZN(n531) );
  INV_X1 U587 ( .A(KEYINPUT88), .ZN(n527) );
  INV_X1 U588 ( .A(G2104), .ZN(n528) );
  NAND2_X1 U589 ( .A1(G126), .A2(n601), .ZN(n525) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n599) );
  NAND2_X1 U591 ( .A1(G114), .A2(n599), .ZN(n524) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n595), .A2(G102), .ZN(n529) );
  AND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n779) );
  AND2_X1 U596 ( .A1(n531), .A2(n779), .ZN(G164) );
  NAND2_X1 U597 ( .A1(G112), .A2(n599), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(KEYINPUT112), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n595), .A2(G100), .ZN(n534) );
  NAND2_X1 U600 ( .A1(G136), .A2(n778), .ZN(n533) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U602 ( .A1(n601), .A2(G124), .ZN(n535) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(n535), .Z(n536) );
  NOR2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(KEYINPUT113), .B(n540), .ZN(G162) );
  NAND2_X1 U607 ( .A1(G101), .A2(n595), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(n541), .Z(n544) );
  NAND2_X1 U609 ( .A1(G113), .A2(n599), .ZN(n542) );
  XOR2_X1 U610 ( .A(KEYINPUT65), .B(n542), .Z(n543) );
  AND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n782) );
  NAND2_X1 U612 ( .A1(G125), .A2(n601), .ZN(n546) );
  NAND2_X1 U613 ( .A1(G137), .A2(n778), .ZN(n545) );
  AND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n783) );
  AND2_X1 U615 ( .A1(n782), .A2(n783), .ZN(G160) );
  NAND2_X1 U616 ( .A1(G99), .A2(n595), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n547), .B(KEYINPUT78), .ZN(n554) );
  NAND2_X1 U618 ( .A1(G111), .A2(n599), .ZN(n549) );
  NAND2_X1 U619 ( .A1(G135), .A2(n778), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n601), .A2(G123), .ZN(n550) );
  XOR2_X1 U622 ( .A(KEYINPUT18), .B(n550), .Z(n551) );
  NOR2_X1 U623 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U624 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U625 ( .A(KEYINPUT79), .B(n555), .Z(n954) );
  XOR2_X1 U626 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n563) );
  NAND2_X1 U627 ( .A1(n595), .A2(G95), .ZN(n557) );
  NAND2_X1 U628 ( .A1(G131), .A2(n778), .ZN(n556) );
  NAND2_X1 U629 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U630 ( .A1(G119), .A2(n601), .ZN(n559) );
  NAND2_X1 U631 ( .A1(G107), .A2(n599), .ZN(n558) );
  NAND2_X1 U632 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U633 ( .A1(n561), .A2(n560), .ZN(n880) );
  XNOR2_X1 U634 ( .A(n880), .B(KEYINPUT46), .ZN(n562) );
  XNOR2_X1 U635 ( .A(n563), .B(n562), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G130), .A2(n601), .ZN(n565) );
  NAND2_X1 U637 ( .A1(G118), .A2(n599), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U639 ( .A(KEYINPUT114), .B(n566), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n595), .A2(G106), .ZN(n568) );
  NAND2_X1 U641 ( .A1(G142), .A2(n778), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U643 ( .A(n569), .B(KEYINPUT45), .Z(n570) );
  NOR2_X1 U644 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U645 ( .A(n573), .B(n572), .Z(n574) );
  XNOR2_X1 U646 ( .A(n954), .B(n574), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n595), .A2(G103), .ZN(n576) );
  NAND2_X1 U648 ( .A1(G139), .A2(n778), .ZN(n575) );
  NAND2_X1 U649 ( .A1(n576), .A2(n575), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n599), .A2(G115), .ZN(n577) );
  XOR2_X1 U651 ( .A(KEYINPUT115), .B(n577), .Z(n579) );
  NAND2_X1 U652 ( .A1(n601), .A2(G127), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U654 ( .A(KEYINPUT47), .B(n580), .Z(n581) );
  NOR2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n942) );
  XNOR2_X1 U656 ( .A(G164), .B(n942), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U658 ( .A(n585), .B(G162), .Z(n594) );
  NAND2_X1 U659 ( .A1(G129), .A2(n601), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G117), .A2(n599), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n595), .A2(G105), .ZN(n588) );
  XOR2_X1 U663 ( .A(KEYINPUT38), .B(n588), .Z(n589) );
  NOR2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U665 ( .A1(G141), .A2(n778), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n875) );
  XOR2_X1 U667 ( .A(G160), .B(n875), .Z(n593) );
  XNOR2_X1 U668 ( .A(n594), .B(n593), .ZN(n608) );
  NAND2_X1 U669 ( .A1(n595), .A2(G104), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G140), .A2(n778), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U672 ( .A(KEYINPUT34), .B(n598), .ZN(n606) );
  NAND2_X1 U673 ( .A1(n599), .A2(G116), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT90), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G128), .A2(n601), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT35), .B(n604), .Z(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U679 ( .A(KEYINPUT36), .B(n607), .Z(n888) );
  XOR2_X1 U680 ( .A(n608), .B(n888), .Z(n609) );
  NOR2_X1 U681 ( .A1(G37), .A2(n609), .ZN(G395) );
  NAND2_X1 U682 ( .A1(n683), .A2(G52), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G64), .A2(n680), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n675), .A2(G90), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G77), .A2(n676), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U688 ( .A(KEYINPUT9), .B(n614), .Z(n615) );
  NOR2_X1 U689 ( .A1(n616), .A2(n615), .ZN(G171) );
  NAND2_X1 U690 ( .A1(G76), .A2(n676), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT74), .B(n617), .ZN(n621) );
  XOR2_X1 U692 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n619) );
  NAND2_X1 U693 ( .A1(G89), .A2(n675), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n622), .B(KEYINPUT5), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n683), .A2(G51), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G63), .A2(n680), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U700 ( .A(KEYINPUT6), .B(n625), .Z(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n628), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U703 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U704 ( .A1(n675), .A2(G88), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G62), .A2(n680), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G75), .A2(n676), .ZN(n631) );
  XNOR2_X1 U708 ( .A(KEYINPUT83), .B(n631), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n683), .A2(G50), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(G303) );
  NAND2_X1 U712 ( .A1(G87), .A2(n636), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n680), .A2(n639), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n683), .A2(G49), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(G288) );
  XOR2_X1 U718 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n643) );
  NAND2_X1 U719 ( .A1(G73), .A2(n676), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n643), .B(n642), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n675), .A2(G86), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G61), .A2(n680), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n683), .A2(G48), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U727 ( .A1(n675), .A2(G91), .ZN(n651) );
  NAND2_X1 U728 ( .A1(G78), .A2(n676), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U730 ( .A(KEYINPUT68), .B(n652), .Z(n656) );
  NAND2_X1 U731 ( .A1(n680), .A2(G65), .ZN(n654) );
  NAND2_X1 U732 ( .A1(n683), .A2(G53), .ZN(n653) );
  AND2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(G299) );
  NAND2_X1 U735 ( .A1(n683), .A2(G54), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G66), .A2(n680), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n675), .A2(G92), .ZN(n660) );
  NAND2_X1 U739 ( .A1(G79), .A2(n676), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U741 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U742 ( .A(n663), .B(KEYINPUT15), .Z(n975) );
  XOR2_X1 U743 ( .A(G286), .B(n975), .Z(n694) );
  NAND2_X1 U744 ( .A1(n675), .A2(G81), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n664), .B(KEYINPUT12), .ZN(n666) );
  NAND2_X1 U746 ( .A1(G68), .A2(n676), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n666), .A2(n665), .ZN(n668) );
  XOR2_X1 U748 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n667) );
  XNOR2_X1 U749 ( .A(n668), .B(n667), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G56), .A2(n680), .ZN(n669) );
  NOR2_X1 U751 ( .A1(n670), .A2(n513), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n683), .A2(G43), .ZN(n671) );
  XNOR2_X1 U753 ( .A(G288), .B(n674), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n675), .A2(G93), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G80), .A2(n676), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U757 ( .A(KEYINPUT80), .B(n679), .Z(n682) );
  NAND2_X1 U758 ( .A1(G67), .A2(n680), .ZN(n681) );
  NAND2_X1 U759 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U760 ( .A1(G55), .A2(n683), .ZN(n684) );
  XNOR2_X1 U761 ( .A(KEYINPUT81), .B(n684), .ZN(n685) );
  OR2_X1 U762 ( .A1(n686), .A2(n685), .ZN(n766) );
  XOR2_X1 U763 ( .A(n766), .B(KEYINPUT19), .Z(n688) );
  XOR2_X1 U764 ( .A(G303), .B(n691), .Z(n693) );
  XNOR2_X1 U765 ( .A(n694), .B(n763), .ZN(n695) );
  XOR2_X1 U766 ( .A(G171), .B(n695), .Z(n696) );
  NOR2_X1 U767 ( .A1(G37), .A2(n696), .ZN(G397) );
  XNOR2_X1 U768 ( .A(G1341), .B(G2454), .ZN(n697) );
  XNOR2_X1 U769 ( .A(n697), .B(G2430), .ZN(n698) );
  XNOR2_X1 U770 ( .A(n698), .B(G1348), .ZN(n704) );
  XOR2_X1 U771 ( .A(G2443), .B(G2427), .Z(n700) );
  XNOR2_X1 U772 ( .A(G2438), .B(G2446), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n700), .B(n699), .ZN(n702) );
  XOR2_X1 U774 ( .A(G2451), .B(G2435), .Z(n701) );
  XNOR2_X1 U775 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U776 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n705), .A2(G14), .ZN(n706) );
  XOR2_X1 U778 ( .A(KEYINPUT104), .B(n706), .Z(G401) );
  XNOR2_X1 U779 ( .A(KEYINPUT86), .B(G44), .ZN(n707) );
  XNOR2_X1 U780 ( .A(n707), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U781 ( .A(G82), .ZN(G220) );
  INV_X1 U782 ( .A(G132), .ZN(G219) );
  INV_X1 U783 ( .A(G57), .ZN(G237) );
  NOR2_X1 U784 ( .A1(G220), .A2(G219), .ZN(n708) );
  XOR2_X1 U785 ( .A(KEYINPUT22), .B(n708), .Z(n709) );
  NOR2_X1 U786 ( .A1(G218), .A2(n709), .ZN(n710) );
  XOR2_X1 U787 ( .A(KEYINPUT87), .B(n710), .Z(n711) );
  NAND2_X1 U788 ( .A1(G96), .A2(n711), .ZN(n915) );
  NAND2_X1 U789 ( .A1(n915), .A2(G2106), .ZN(n715) );
  NAND2_X1 U790 ( .A1(G69), .A2(G120), .ZN(n712) );
  NOR2_X1 U791 ( .A1(G237), .A2(n712), .ZN(n713) );
  NAND2_X1 U792 ( .A1(G108), .A2(n713), .ZN(n914) );
  NAND2_X1 U793 ( .A1(n914), .A2(G567), .ZN(n714) );
  NAND2_X1 U794 ( .A1(n715), .A2(n714), .ZN(n775) );
  INV_X1 U795 ( .A(n775), .ZN(G319) );
  XOR2_X1 U796 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n717) );
  XNOR2_X1 U797 ( .A(G2678), .B(KEYINPUT43), .ZN(n716) );
  XNOR2_X1 U798 ( .A(n717), .B(n716), .ZN(n721) );
  XOR2_X1 U799 ( .A(KEYINPUT42), .B(G2090), .Z(n719) );
  INV_X1 U800 ( .A(G2072), .ZN(n1001) );
  XOR2_X1 U801 ( .A(G2067), .B(n1001), .Z(n718) );
  XNOR2_X1 U802 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U803 ( .A(n721), .B(n720), .Z(n723) );
  XNOR2_X1 U804 ( .A(G2096), .B(G2100), .ZN(n722) );
  XNOR2_X1 U805 ( .A(n723), .B(n722), .ZN(n725) );
  XOR2_X1 U806 ( .A(G2078), .B(G2084), .Z(n724) );
  XNOR2_X1 U807 ( .A(n725), .B(n724), .ZN(G227) );
  XOR2_X1 U808 ( .A(KEYINPUT111), .B(G1976), .Z(n727) );
  INV_X1 U809 ( .A(G1971), .ZN(n982) );
  XOR2_X1 U810 ( .A(G1986), .B(n982), .Z(n726) );
  XNOR2_X1 U811 ( .A(n727), .B(n726), .ZN(n728) );
  XOR2_X1 U812 ( .A(n728), .B(KEYINPUT41), .Z(n730) );
  INV_X1 U813 ( .A(G1991), .ZN(n881) );
  XOR2_X1 U814 ( .A(G1996), .B(n881), .Z(n729) );
  XNOR2_X1 U815 ( .A(n730), .B(n729), .ZN(n734) );
  XOR2_X1 U816 ( .A(G1956), .B(G1961), .Z(n732) );
  XNOR2_X1 U817 ( .A(G1981), .B(G1966), .ZN(n731) );
  XNOR2_X1 U818 ( .A(n732), .B(n731), .ZN(n733) );
  XOR2_X1 U819 ( .A(n734), .B(n733), .Z(n736) );
  XNOR2_X1 U820 ( .A(G2474), .B(KEYINPUT110), .ZN(n735) );
  XNOR2_X1 U821 ( .A(n736), .B(n735), .ZN(G229) );
  NOR2_X1 U822 ( .A1(G395), .A2(G397), .ZN(n738) );
  XNOR2_X1 U823 ( .A(n738), .B(n737), .ZN(n743) );
  NOR2_X1 U824 ( .A1(G227), .A2(G229), .ZN(n739) );
  XOR2_X1 U825 ( .A(KEYINPUT49), .B(n739), .Z(n740) );
  NAND2_X1 U826 ( .A1(G319), .A2(n740), .ZN(n741) );
  NOR2_X1 U827 ( .A1(G401), .A2(n741), .ZN(n742) );
  NAND2_X1 U828 ( .A1(n743), .A2(n742), .ZN(G225) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  XNOR2_X1 U830 ( .A(G2096), .B(n954), .ZN(n744) );
  OR2_X1 U831 ( .A1(G2100), .A2(n744), .ZN(G156) );
  NAND2_X1 U832 ( .A1(G7), .A2(G661), .ZN(n745) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U834 ( .A(G223), .B(KEYINPUT69), .ZN(n909) );
  NAND2_X1 U835 ( .A1(n909), .A2(G567), .ZN(n746) );
  XOR2_X1 U836 ( .A(KEYINPUT11), .B(n746), .Z(G234) );
  XNOR2_X1 U837 ( .A(G860), .B(KEYINPUT71), .ZN(n751) );
  OR2_X1 U838 ( .A1(n972), .A2(n751), .ZN(G153) );
  XOR2_X1 U839 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U840 ( .A1(G868), .A2(G301), .ZN(n748) );
  INV_X1 U841 ( .A(n975), .ZN(n805) );
  INV_X1 U842 ( .A(G868), .ZN(n765) );
  NAND2_X1 U843 ( .A1(n805), .A2(n765), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n748), .A2(n747), .ZN(G284) );
  NOR2_X1 U845 ( .A1(G286), .A2(n765), .ZN(n750) );
  NOR2_X1 U846 ( .A1(G868), .A2(G299), .ZN(n749) );
  NOR2_X1 U847 ( .A1(n750), .A2(n749), .ZN(G297) );
  NAND2_X1 U848 ( .A1(G559), .A2(n751), .ZN(n752) );
  XOR2_X1 U849 ( .A(KEYINPUT75), .B(n752), .Z(n753) );
  NAND2_X1 U850 ( .A1(n753), .A2(n975), .ZN(n754) );
  XNOR2_X1 U851 ( .A(n754), .B(KEYINPUT76), .ZN(n755) );
  XNOR2_X1 U852 ( .A(KEYINPUT16), .B(n755), .ZN(G148) );
  NOR2_X1 U853 ( .A1(G559), .A2(n765), .ZN(n756) );
  NAND2_X1 U854 ( .A1(n975), .A2(n756), .ZN(n757) );
  XNOR2_X1 U855 ( .A(n757), .B(KEYINPUT77), .ZN(n759) );
  NOR2_X1 U856 ( .A1(n972), .A2(G868), .ZN(n758) );
  NOR2_X1 U857 ( .A1(n759), .A2(n758), .ZN(G282) );
  NAND2_X1 U858 ( .A1(n975), .A2(G559), .ZN(n762) );
  XNOR2_X1 U859 ( .A(n972), .B(n762), .ZN(n760) );
  NOR2_X1 U860 ( .A1(n760), .A2(G860), .ZN(n761) );
  XOR2_X1 U861 ( .A(n761), .B(n766), .Z(G145) );
  XOR2_X1 U862 ( .A(n763), .B(n762), .Z(n764) );
  NOR2_X1 U863 ( .A1(n765), .A2(n764), .ZN(n768) );
  NOR2_X1 U864 ( .A1(G868), .A2(n766), .ZN(n767) );
  NOR2_X1 U865 ( .A1(n768), .A2(n767), .ZN(G295) );
  NAND2_X1 U866 ( .A1(G2078), .A2(G2084), .ZN(n769) );
  XNOR2_X1 U867 ( .A(n769), .B(KEYINPUT85), .ZN(n770) );
  XNOR2_X1 U868 ( .A(n770), .B(KEYINPUT20), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n771), .A2(G2090), .ZN(n772) );
  XNOR2_X1 U870 ( .A(KEYINPUT21), .B(n772), .ZN(n773) );
  NAND2_X1 U871 ( .A1(n773), .A2(G2072), .ZN(G158) );
  NAND2_X1 U872 ( .A1(G483), .A2(G661), .ZN(n774) );
  NOR2_X1 U873 ( .A1(n775), .A2(n774), .ZN(n913) );
  NAND2_X1 U874 ( .A1(n913), .A2(G36), .ZN(G176) );
  INV_X1 U875 ( .A(G303), .ZN(G166) );
  XOR2_X1 U876 ( .A(G1981), .B(G305), .Z(n990) );
  INV_X1 U877 ( .A(KEYINPUT32), .ZN(n842) );
  XOR2_X1 U878 ( .A(KEYINPUT92), .B(G1961), .Z(n923) );
  INV_X1 U879 ( .A(G1384), .ZN(n776) );
  AND2_X1 U880 ( .A1(G138), .A2(n776), .ZN(n777) );
  NAND2_X1 U881 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U882 ( .A1(n781), .A2(n780), .ZN(n879) );
  INV_X1 U883 ( .A(n879), .ZN(n785) );
  AND2_X1 U884 ( .A1(n782), .A2(G40), .ZN(n784) );
  NAND2_X1 U885 ( .A1(n784), .A2(n783), .ZN(n878) );
  NOR2_X2 U886 ( .A1(n785), .A2(n878), .ZN(n790) );
  INV_X1 U887 ( .A(n790), .ZN(n817) );
  NAND2_X1 U888 ( .A1(n923), .A2(n829), .ZN(n787) );
  XNOR2_X1 U889 ( .A(G2078), .B(KEYINPUT25), .ZN(n1000) );
  NAND2_X1 U890 ( .A1(n790), .A2(n1000), .ZN(n786) );
  NAND2_X1 U891 ( .A1(n787), .A2(n786), .ZN(n823) );
  NAND2_X1 U892 ( .A1(n823), .A2(G171), .ZN(n816) );
  NOR2_X1 U893 ( .A1(n790), .A2(G1348), .ZN(n789) );
  NOR2_X1 U894 ( .A1(G2067), .A2(n829), .ZN(n788) );
  NOR2_X1 U895 ( .A1(n789), .A2(n788), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n805), .A2(n806), .ZN(n797) );
  NAND2_X1 U897 ( .A1(G1996), .A2(n790), .ZN(n791) );
  XNOR2_X1 U898 ( .A(n791), .B(KEYINPUT26), .ZN(n793) );
  NAND2_X1 U899 ( .A1(G1341), .A2(n829), .ZN(n792) );
  NAND2_X1 U900 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U901 ( .A(KEYINPUT94), .B(n794), .ZN(n795) );
  NOR2_X1 U902 ( .A1(n972), .A2(n795), .ZN(n796) );
  NAND2_X1 U903 ( .A1(n797), .A2(n796), .ZN(n804) );
  NOR2_X1 U904 ( .A1(n817), .A2(n1001), .ZN(n799) );
  XOR2_X1 U905 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n798) );
  XNOR2_X1 U906 ( .A(n799), .B(n798), .ZN(n801) );
  NAND2_X1 U907 ( .A1(n829), .A2(G1956), .ZN(n800) );
  NAND2_X1 U908 ( .A1(n801), .A2(n800), .ZN(n809) );
  NOR2_X1 U909 ( .A1(G299), .A2(n809), .ZN(n802) );
  XNOR2_X1 U910 ( .A(KEYINPUT95), .B(n802), .ZN(n803) );
  NAND2_X1 U911 ( .A1(n804), .A2(n803), .ZN(n808) );
  NOR2_X1 U912 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U913 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U914 ( .A1(G299), .A2(n809), .ZN(n810) );
  XOR2_X1 U915 ( .A(KEYINPUT28), .B(n810), .Z(n811) );
  NOR2_X1 U916 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U917 ( .A1(n816), .A2(n815), .ZN(n844) );
  NAND2_X1 U918 ( .A1(G8), .A2(n817), .ZN(n872) );
  NOR2_X1 U919 ( .A1(G1966), .A2(n872), .ZN(n849) );
  NOR2_X1 U920 ( .A1(G2084), .A2(n829), .ZN(n845) );
  NOR2_X1 U921 ( .A1(n849), .A2(n845), .ZN(n818) );
  NAND2_X1 U922 ( .A1(n818), .A2(G8), .ZN(n821) );
  NOR2_X1 U923 ( .A1(G168), .A2(n822), .ZN(n825) );
  NOR2_X1 U924 ( .A1(G171), .A2(n823), .ZN(n824) );
  NOR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(n827) );
  INV_X1 U926 ( .A(KEYINPUT31), .ZN(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n843) );
  INV_X1 U928 ( .A(G8), .ZN(n835) );
  NOR2_X1 U929 ( .A1(G1971), .A2(n872), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n828), .B(KEYINPUT98), .ZN(n831) );
  NOR2_X1 U931 ( .A1(n829), .A2(G2090), .ZN(n830) );
  NOR2_X1 U932 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U933 ( .A1(n832), .A2(G303), .ZN(n833) );
  XOR2_X1 U934 ( .A(KEYINPUT99), .B(n833), .Z(n834) );
  OR2_X1 U935 ( .A1(n835), .A2(n834), .ZN(n837) );
  AND2_X1 U936 ( .A1(n843), .A2(n837), .ZN(n836) );
  NAND2_X1 U937 ( .A1(n844), .A2(n836), .ZN(n840) );
  INV_X1 U938 ( .A(n837), .ZN(n838) );
  OR2_X1 U939 ( .A1(n838), .A2(G286), .ZN(n839) );
  NAND2_X1 U940 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n851) );
  NAND2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n847) );
  NAND2_X1 U943 ( .A1(G8), .A2(n845), .ZN(n846) );
  NAND2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U946 ( .A1(G1976), .A2(G288), .ZN(n858) );
  NOR2_X1 U947 ( .A1(G1971), .A2(G303), .ZN(n852) );
  NOR2_X1 U948 ( .A1(n858), .A2(n852), .ZN(n981) );
  XOR2_X1 U949 ( .A(n981), .B(KEYINPUT100), .Z(n853) );
  NOR2_X1 U950 ( .A1(n866), .A2(n853), .ZN(n855) );
  INV_X1 U951 ( .A(n872), .ZN(n868) );
  NAND2_X1 U952 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NAND2_X1 U953 ( .A1(n868), .A2(n980), .ZN(n854) );
  XOR2_X1 U954 ( .A(n856), .B(KEYINPUT64), .Z(n857) );
  NOR2_X1 U955 ( .A1(KEYINPUT33), .A2(n857), .ZN(n861) );
  NAND2_X1 U956 ( .A1(n858), .A2(KEYINPUT33), .ZN(n859) );
  NOR2_X1 U957 ( .A1(n859), .A2(n872), .ZN(n860) );
  NOR2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n990), .A2(n862), .ZN(n863) );
  XNOR2_X1 U960 ( .A(KEYINPUT101), .B(n863), .ZN(n897) );
  NAND2_X1 U961 ( .A1(G166), .A2(G8), .ZN(n864) );
  NOR2_X1 U962 ( .A1(G2090), .A2(n864), .ZN(n865) );
  NOR2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U965 ( .A(KEYINPUT102), .B(n869), .Z(n874) );
  NOR2_X1 U966 ( .A1(G1981), .A2(G305), .ZN(n870) );
  XOR2_X1 U967 ( .A(n870), .B(KEYINPUT24), .Z(n871) );
  OR2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n895) );
  XOR2_X1 U970 ( .A(KEYINPUT37), .B(G2067), .Z(n889) );
  OR2_X1 U971 ( .A1(n889), .A2(n888), .ZN(n947) );
  NOR2_X1 U972 ( .A1(G1996), .A2(n875), .ZN(n950) );
  NOR2_X1 U973 ( .A1(n880), .A2(n881), .ZN(n877) );
  AND2_X1 U974 ( .A1(G1996), .A2(n875), .ZN(n876) );
  OR2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n953) );
  NOR2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n899) );
  NAND2_X1 U977 ( .A1(n953), .A2(n899), .ZN(n900) );
  INV_X1 U978 ( .A(n900), .ZN(n885) );
  AND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT103), .B(n882), .Z(n952) );
  NOR2_X1 U981 ( .A1(G1986), .A2(G290), .ZN(n883) );
  NOR2_X1 U982 ( .A1(n952), .A2(n883), .ZN(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U984 ( .A1(n950), .A2(n886), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(KEYINPUT39), .ZN(n891) );
  NAND2_X1 U986 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(KEYINPUT91), .B(n890), .ZN(n961) );
  NAND2_X1 U988 ( .A1(n899), .A2(n961), .ZN(n901) );
  NAND2_X1 U989 ( .A1(n891), .A2(n901), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n947), .A2(n892), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n893), .A2(n899), .ZN(n905) );
  INV_X1 U992 ( .A(n905), .ZN(n894) );
  OR2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n896) );
  NOR2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n907) );
  XOR2_X1 U995 ( .A(G1986), .B(KEYINPUT89), .Z(n898) );
  XNOR2_X1 U996 ( .A(G290), .B(n898), .ZN(n977) );
  AND2_X1 U997 ( .A1(n977), .A2(n899), .ZN(n903) );
  NAND2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  OR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n904) );
  AND2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n908), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U1003 ( .A1(n909), .A2(G2106), .ZN(n910) );
  XOR2_X1 U1004 ( .A(KEYINPUT105), .B(n910), .Z(G217) );
  AND2_X1 U1005 ( .A1(G15), .A2(G2), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G661), .A2(n911), .ZN(G259) );
  NAND2_X1 U1007 ( .A1(G3), .A2(G1), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(G188) );
  XOR2_X1 U1009 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  XOR2_X1 U1010 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  INV_X1 U1012 ( .A(G120), .ZN(G236) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1015 ( .A(n916), .B(KEYINPUT107), .Z(G325) );
  INV_X1 U1016 ( .A(G325), .ZN(G261) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1018 ( .A(G1986), .B(G24), .ZN(n921) );
  XOR2_X1 U1019 ( .A(n982), .B(G22), .Z(n918) );
  XNOR2_X1 U1020 ( .A(G1976), .B(G23), .ZN(n917) );
  NOR2_X1 U1021 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(KEYINPUT127), .B(n919), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(KEYINPUT58), .B(n922), .ZN(n927) );
  XOR2_X1 U1025 ( .A(n923), .B(G5), .Z(n925) );
  XNOR2_X1 U1026 ( .A(G21), .B(G1966), .ZN(n924) );
  NOR2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n938) );
  XNOR2_X1 U1029 ( .A(G1341), .B(G19), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G20), .B(G1956), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n935) );
  XOR2_X1 U1032 ( .A(G4), .B(KEYINPUT126), .Z(n931) );
  XNOR2_X1 U1033 ( .A(G1348), .B(KEYINPUT59), .ZN(n930) );
  XNOR2_X1 U1034 ( .A(n931), .B(n930), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(G1981), .B(G6), .ZN(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(KEYINPUT60), .B(n936), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(KEYINPUT61), .B(n939), .ZN(n940) );
  INV_X1 U1041 ( .A(G16), .ZN(n971) );
  NAND2_X1 U1042 ( .A1(n940), .A2(n971), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n941), .A2(G11), .ZN(n970) );
  XOR2_X1 U1044 ( .A(G164), .B(G2078), .Z(n944) );
  XOR2_X1 U1045 ( .A(G2072), .B(n942), .Z(n943) );
  NOR2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(KEYINPUT120), .B(n945), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(n946), .B(KEYINPUT50), .ZN(n948) );
  NAND2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n964) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n951), .Z(n959) );
  OR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G160), .B(G2084), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(n962), .B(KEYINPUT119), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n965), .B(KEYINPUT52), .ZN(n966) );
  INV_X1 U1062 ( .A(KEYINPUT55), .ZN(n1020) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n1020), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(G29), .A2(n967), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT121), .B(n968), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n999) );
  XOR2_X1 U1067 ( .A(n971), .B(KEYINPUT56), .Z(n997) );
  XNOR2_X1 U1068 ( .A(n972), .B(G1341), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G299), .B(G1956), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n989) );
  XNOR2_X1 U1071 ( .A(G171), .B(G1961), .ZN(n979) );
  XOR2_X1 U1072 ( .A(G1348), .B(n975), .Z(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(G166), .A2(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1078 ( .A(KEYINPUT124), .B(n985), .Z(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1083 ( .A(KEYINPUT57), .B(n992), .Z(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(KEYINPUT125), .B(n995), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1023) );
  XNOR2_X1 U1088 ( .A(G27), .B(n1000), .ZN(n1012) );
  XOR2_X1 U1089 ( .A(KEYINPUT123), .B(n1001), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(n1002), .B(G33), .ZN(n1007) );
  XOR2_X1 U1091 ( .A(G32), .B(G1996), .Z(n1003) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(G28), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G26), .B(G2067), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G25), .B(G1991), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT122), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT53), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(G2084), .B(G34), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT54), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G35), .B(G2090), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1110 ( .A(G150), .ZN(G311) );
endmodule

