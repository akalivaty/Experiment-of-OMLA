//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(G50), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n209), .A2(new_n211), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n223), .A2(new_n224), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n207), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n217), .B(new_n231), .C1(new_n209), .C2(new_n211), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT67), .B(G50), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT71), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  AND2_X1   g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(new_n253), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n256), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G223), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G222), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n263), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n259), .B1(new_n269), .B2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n267), .B(new_n271), .C1(new_n268), .C2(new_n263), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n262), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G190), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n212), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G150), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n213), .A2(G33), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n203), .ZN(new_n285));
  INV_X1    g0085(.A(G50), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n213), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n279), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n277), .A2(new_n212), .A3(new_n278), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n213), .A2(G1), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n289), .A2(G50), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n286), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n274), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n273), .A2(new_n300), .B1(new_n297), .B2(KEYINPUT9), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT10), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n270), .A2(new_n272), .ZN(new_n303));
  INV_X1    g0103(.A(new_n262), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n305), .A2(G200), .B1(new_n306), .B2(new_n296), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n273), .A2(G190), .B1(new_n297), .B2(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(G20), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n313), .A2(new_n315), .B1(G20), .B2(G77), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n282), .B(KEYINPUT70), .ZN(new_n317));
  INV_X1    g0117(.A(new_n280), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n279), .B1(new_n268), .B2(new_n294), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n279), .A2(new_n294), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G77), .A3(new_n292), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n324), .A2(new_n251), .A3(new_n256), .ZN(new_n325));
  INV_X1    g0125(.A(new_n260), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(G244), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G232), .A2(G1698), .ZN(new_n328));
  INV_X1    g0128(.A(G1698), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G238), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n263), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n331), .B(new_n324), .C1(G107), .C2(new_n263), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n327), .A2(new_n332), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n323), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(G190), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(G200), .ZN(new_n341));
  AND4_X1   g0141(.A1(new_n322), .A2(new_n340), .A3(new_n320), .A4(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n305), .A2(G179), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n296), .B1(new_n273), .B2(G169), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AND4_X1   g0147(.A1(new_n250), .A2(new_n311), .A3(new_n343), .A4(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n346), .B1(new_n302), .B2(new_n310), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n250), .B1(new_n349), .B2(new_n343), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n282), .A2(new_n291), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n321), .A2(new_n352), .B1(new_n294), .B2(new_n282), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n201), .A2(new_n202), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n285), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n280), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT3), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(G33), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT7), .B(new_n213), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n367), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n213), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n263), .B2(G20), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n358), .B1(new_n371), .B2(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n289), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(new_n358), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n365), .A2(new_n366), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n359), .A2(KEYINPUT76), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n369), .A2(G20), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n202), .B1(new_n380), .B2(new_n370), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n375), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI211_X1 g0183(.A(KEYINPUT77), .B(new_n202), .C1(new_n380), .C2(new_n370), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n374), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n354), .B1(new_n373), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n329), .A2(G223), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT78), .B1(new_n367), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT78), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n263), .A2(new_n389), .A3(G223), .A4(new_n329), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n365), .A2(new_n366), .A3(G226), .A4(G1698), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n259), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n258), .B1(new_n260), .B2(new_n234), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n397), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n394), .B1(new_n390), .B2(new_n388), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(G179), .C1(new_n400), .C2(new_n259), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT18), .B1(new_n386), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n380), .A2(new_n370), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n358), .B1(new_n405), .B2(KEYINPUT77), .ZN(new_n406));
  INV_X1    g0206(.A(new_n384), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT16), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n368), .A2(new_n370), .ZN(new_n409));
  AOI21_X1  g0209(.A(G20), .B1(new_n365), .B2(new_n366), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT75), .B1(new_n410), .B2(KEYINPUT7), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n375), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n279), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n353), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n398), .A2(new_n401), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n403), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n300), .B1(new_n396), .B2(new_n397), .ZN(new_n420));
  INV_X1    g0220(.A(G190), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n399), .B(new_n421), .C1(new_n400), .C2(new_n259), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n353), .B(new_n423), .C1(new_n408), .C2(new_n414), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n423), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT73), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n318), .B2(new_n286), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n280), .A2(KEYINPUT73), .A3(G50), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n283), .A2(new_n268), .B1(new_n213), .B2(G68), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(KEYINPUT72), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n279), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT11), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n291), .A2(new_n202), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT12), .B1(new_n290), .B2(G68), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n290), .A2(KEYINPUT12), .A3(G68), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n321), .A2(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n435), .B2(new_n436), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n234), .A2(G1698), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n263), .B(new_n444), .C1(G226), .C2(G1698), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G97), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n324), .ZN(new_n448));
  INV_X1    g0248(.A(G238), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n258), .B1(new_n260), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT13), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n259), .B1(new_n445), .B2(new_n446), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT13), .B1(new_n454), .B2(new_n450), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(G190), .A3(new_n455), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n443), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT74), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT74), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n443), .A2(new_n457), .A3(new_n461), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n437), .A2(new_n442), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(new_n465), .A3(G169), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n453), .A2(G179), .A3(new_n455), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n456), .B2(G169), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n419), .A2(new_n428), .A3(new_n463), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n351), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n329), .A2(G264), .ZN(new_n473));
  NOR2_X1   g0273(.A1(G257), .A2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n365), .B(new_n366), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G303), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n359), .B2(new_n361), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n477), .A3(new_n324), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n254), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G270), .A3(new_n259), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n478), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n487), .A2(G169), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n255), .A2(G33), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n321), .A2(G116), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n290), .A2(G116), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G20), .B1(G33), .B2(G283), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n314), .A2(G97), .ZN(new_n494));
  INV_X1    g0294(.A(G116), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n493), .A2(new_n494), .B1(G20), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n279), .A2(KEYINPUT20), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT20), .B1(new_n279), .B2(new_n496), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n490), .B(new_n492), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n488), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n487), .A2(G200), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n504), .C1(new_n421), .C2(new_n487), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n487), .A2(KEYINPUT21), .A3(G169), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n478), .A2(G179), .A3(new_n482), .A4(new_n486), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n508), .A2(KEYINPUT80), .A3(new_n499), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT80), .B1(new_n508), .B2(new_n499), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n502), .B(new_n505), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G244), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G1698), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT4), .B1(new_n263), .B2(new_n514), .ZN(new_n515));
  AND4_X1   g0315(.A1(KEYINPUT4), .A2(new_n514), .A3(new_n365), .A4(new_n366), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n365), .A2(new_n366), .A3(G250), .A4(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n259), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n485), .A2(G257), .A3(new_n259), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n482), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n334), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n514), .A2(new_n365), .A3(new_n366), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n514), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n519), .A4(new_n518), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n523), .B1(new_n529), .B2(new_n324), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n337), .ZN(new_n531));
  INV_X1    g0331(.A(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n221), .A2(new_n532), .A3(KEYINPUT6), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(KEYINPUT79), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT79), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G107), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n533), .A2(new_n535), .A3(new_n537), .A4(new_n539), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n532), .B1(new_n380), .B2(new_n370), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n289), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n290), .A2(G97), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n321), .A2(new_n489), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n221), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n524), .B(new_n531), .C1(new_n547), .C2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G200), .B1(new_n521), .B2(new_n523), .ZN(new_n553));
  INV_X1    g0353(.A(new_n542), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n533), .A2(new_n535), .B1(new_n537), .B2(new_n539), .ZN(new_n555));
  OAI21_X1  g0355(.A(G20), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n280), .A2(G77), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n279), .B1(new_n558), .B2(new_n545), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n530), .A2(G190), .ZN(new_n560));
  INV_X1    g0360(.A(new_n551), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n553), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n213), .B1(new_n446), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n219), .A2(new_n221), .A3(new_n532), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n365), .A2(new_n366), .A3(new_n213), .A4(G68), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n563), .B1(new_n283), .B2(new_n221), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n279), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n289), .A2(new_n290), .A3(new_n313), .A4(new_n489), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n312), .A2(new_n294), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n254), .A2(new_n480), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n220), .B1(new_n255), .B2(G45), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n259), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n449), .A2(new_n329), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n513), .A2(G1698), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n365), .A2(new_n578), .A3(new_n366), .A4(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n314), .A2(new_n495), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n259), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n334), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n254), .A2(new_n480), .B1(new_n259), .B2(new_n575), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G238), .A2(G1698), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n513), .B2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n581), .B1(new_n587), .B2(new_n263), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n585), .B(new_n337), .C1(new_n588), .C2(new_n259), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n573), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(G200), .B1(new_n577), .B2(new_n583), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n321), .A2(G87), .A3(new_n489), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n569), .A2(new_n279), .B1(new_n294), .B2(new_n312), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n585), .B(G190), .C1(new_n588), .C2(new_n259), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n552), .A2(new_n562), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n485), .A2(G264), .A3(new_n259), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G250), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n222), .B2(G1698), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n263), .B1(G33), .B2(G294), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n482), .B(new_n598), .C1(new_n601), .C2(new_n259), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n602), .A2(G179), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n334), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n294), .A2(new_n532), .ZN(new_n605));
  XOR2_X1   g0405(.A(new_n605), .B(KEYINPUT25), .Z(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n550), .B2(new_n532), .ZN(new_n607));
  AND2_X1   g0407(.A1(KEYINPUT81), .A2(G87), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n365), .A2(new_n366), .A3(new_n608), .A4(new_n213), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT22), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n263), .A2(KEYINPUT22), .A3(new_n213), .A4(new_n608), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT23), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n213), .B2(G107), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n532), .A2(KEYINPUT23), .A3(G20), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n615), .B1(new_n581), .B2(new_n213), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g0417(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n618), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n611), .A2(new_n612), .A3(new_n616), .A4(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n289), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n603), .B(new_n604), .C1(new_n607), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n602), .A2(new_n300), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G190), .B2(new_n602), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n619), .A2(new_n621), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n279), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n605), .B(KEYINPUT25), .ZN(new_n628));
  INV_X1    g0428(.A(new_n550), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(G107), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n597), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n472), .A2(new_n512), .A3(new_n633), .ZN(G372));
  AND2_X1   g0434(.A1(new_n508), .A2(new_n499), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT21), .B1(new_n488), .B2(new_n499), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT84), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n508), .A2(new_n499), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n502), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n623), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n591), .A2(KEYINPUT83), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n585), .B1(new_n588), .B2(new_n259), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT83), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(G200), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n593), .A2(new_n594), .A3(new_n592), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n590), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n552), .A2(new_n631), .A3(new_n562), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n641), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n552), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n596), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT26), .B1(new_n655), .B2(new_n552), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n656), .A3(new_n590), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n472), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n470), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n339), .A2(new_n459), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n428), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n419), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n346), .B1(new_n662), .B2(new_n311), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n658), .A2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n255), .A2(new_n213), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n503), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n511), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n637), .A2(new_n640), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n671), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G330), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT85), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n670), .B1(new_n627), .B2(new_n630), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n632), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n623), .B2(new_n670), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n623), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n670), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n670), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(new_n686), .A3(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n208), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n565), .A2(G116), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n692), .A2(new_n255), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n692), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n696), .B(KEYINPUT86), .C1(new_n216), .C2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(KEYINPUT86), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  OAI21_X1  g0500(.A(new_n670), .B1(new_n651), .B2(new_n657), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n670), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT26), .B1(new_n648), .B2(new_n552), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n524), .A2(new_n531), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n559), .A2(new_n561), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n596), .A3(new_n653), .A4(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n705), .A2(new_n590), .A3(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n650), .B(new_n649), .C1(new_n687), .C2(new_n685), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT88), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT29), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n711), .B2(KEYINPUT29), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n703), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n602), .A2(new_n487), .A3(new_n337), .A4(new_n643), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n530), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n598), .B1(new_n601), .B2(new_n259), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n643), .ZN(new_n721));
  INV_X1    g0521(.A(new_n507), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n530), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n507), .A2(new_n720), .A3(new_n643), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n530), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n719), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n704), .B1(new_n728), .B2(KEYINPUT87), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT87), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n730), .B(new_n719), .C1(new_n724), .C2(new_n727), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n717), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n512), .A2(new_n633), .A3(new_n670), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n726), .B1(new_n725), .B2(new_n530), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n735), .B1(new_n530), .B2(new_n718), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n732), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n716), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n700), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(new_n678), .ZN(new_n743));
  INV_X1    g0543(.A(G13), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n255), .B1(new_n745), .B2(G45), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n697), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n676), .A2(new_n677), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n743), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n213), .A2(new_n300), .A3(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G87), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n213), .A2(new_n337), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n753), .B1(new_n757), .B2(new_n201), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n754), .A2(new_n421), .A3(new_n300), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n213), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n337), .A3(new_n300), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n263), .B1(new_n268), .B2(new_n759), .C1(new_n763), .C2(new_n202), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n755), .A2(new_n300), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n758), .B(new_n764), .C1(G50), .C2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n750), .A2(new_n421), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT91), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT91), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G107), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT90), .ZN(new_n774));
  OAI21_X1  g0574(.A(G20), .B1(new_n774), .B2(new_n421), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n766), .B(new_n772), .C1(new_n221), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(new_n761), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G159), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT33), .B(G317), .Z(new_n782));
  OAI221_X1 g0582(.A(new_n367), .B1(new_n759), .B2(new_n781), .C1(new_n763), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G329), .B2(new_n778), .ZN(new_n784));
  INV_X1    g0584(.A(G322), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n757), .A2(new_n785), .B1(new_n476), .B2(new_n751), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G326), .B2(new_n765), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n770), .A2(new_n789), .B1(new_n790), .B2(new_n776), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n777), .A2(new_n780), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n212), .B1(G20), .B2(new_n334), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n691), .A2(new_n367), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G355), .B1(new_n495), .B2(new_n691), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n245), .A2(new_n479), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n691), .A2(new_n263), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n216), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT89), .Z(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n793), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n747), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n803), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n794), .B(new_n805), .C1(new_n675), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n749), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT92), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NAND3_X1  g0610(.A1(new_n323), .A2(new_n335), .A3(new_n338), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n704), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n670), .B1(new_n320), .B2(new_n322), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n811), .B1(new_n342), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n701), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n816), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n818), .B(new_n670), .C1(new_n651), .C2(new_n657), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n740), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT96), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n822), .B(new_n747), .C1(new_n740), .C2(new_n820), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n793), .A2(new_n801), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n747), .B1(new_n268), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n771), .A2(G68), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n263), .B1(new_n751), .B2(new_n286), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n778), .B2(G132), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(new_n201), .C2(new_n776), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT94), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  INV_X1    g0632(.A(new_n759), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G150), .A2(new_n762), .B1(new_n833), .B2(G159), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(new_n765), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n834), .B1(new_n835), .B2(new_n836), .C1(new_n837), .C2(new_n757), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT34), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n831), .A2(new_n832), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n770), .A2(new_n219), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G311), .B2(new_n778), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT93), .Z(new_n843));
  AOI22_X1  g0643(.A1(G107), .A2(new_n752), .B1(new_n756), .B2(G294), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n476), .B2(new_n836), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n367), .B1(new_n495), .B2(new_n759), .C1(new_n763), .C2(new_n789), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n221), .B2(new_n776), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n840), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT95), .ZN(new_n850));
  INV_X1    g0650(.A(new_n793), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n825), .B1(new_n802), .B2(new_n818), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n823), .A2(new_n852), .ZN(G384));
  OAI21_X1  g0653(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n216), .A2(new_n854), .B1(G50), .B2(new_n202), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(G1), .A3(new_n744), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT97), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n495), .B(new_n215), .C1(new_n543), .C2(KEYINPUT35), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(KEYINPUT35), .B2(new_n543), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT36), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n403), .A2(new_n426), .A3(new_n418), .A4(new_n427), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n412), .A2(new_n375), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n374), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n354), .B1(new_n373), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n668), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n424), .B1(new_n386), .B2(new_n402), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n386), .B2(new_n668), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT98), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n372), .A2(KEYINPUT16), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n353), .B1(new_n414), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n398), .A2(new_n401), .A3(new_n668), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n870), .B1(new_n877), .B2(new_n424), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n872), .A2(new_n873), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT37), .B1(new_n415), .B2(new_n669), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n415), .A2(new_n417), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n424), .ZN(new_n882));
  INV_X1    g0682(.A(new_n876), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n424), .B1(new_n866), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT98), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT38), .B(new_n868), .C1(new_n879), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n415), .A2(new_n669), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n419), .B2(new_n428), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n881), .A2(new_n889), .A3(new_n424), .ZN(new_n891));
  INV_X1    g0691(.A(new_n869), .ZN(new_n892));
  AOI22_X1  g0692(.A1(KEYINPUT37), .A2(new_n891), .B1(new_n892), .B2(new_n880), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n888), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT39), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n887), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n873), .B1(new_n872), .B2(new_n878), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT98), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n899), .B2(new_n868), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n895), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n659), .A2(new_n670), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT99), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n419), .A2(new_n669), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n819), .A2(new_n813), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n464), .A2(new_n704), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n459), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n470), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n456), .A2(G169), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT14), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n467), .A3(new_n466), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n460), .B2(new_n462), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n912), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n868), .B1(new_n879), .B2(new_n886), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n888), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n887), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n907), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n906), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n472), .B(new_n703), .C1(new_n713), .C2(new_n714), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n663), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n887), .A2(new_n894), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n736), .A2(new_n730), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n728), .A2(KEYINPUT87), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT31), .A4(new_n704), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n732), .A2(new_n733), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n818), .A3(new_n917), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n928), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n922), .A2(new_n928), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n472), .A2(new_n933), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n677), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n927), .A2(new_n942), .B1(new_n255), .B2(new_n745), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT100), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n927), .A2(new_n942), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n862), .B1(new_n945), .B2(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n593), .A2(new_n592), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n704), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n649), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n590), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT43), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n652), .A2(new_n704), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n707), .A2(new_n704), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(new_n552), .A3(new_n562), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n689), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n961), .B(KEYINPUT101), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n652), .B1(new_n965), .B2(new_n685), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT102), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n704), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n954), .B(new_n957), .C1(new_n964), .C2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n964), .A2(new_n969), .A3(new_n956), .A4(new_n955), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n965), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n684), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n970), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n970), .B2(new_n972), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n692), .B(KEYINPUT41), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n689), .A2(new_n686), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n962), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT44), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n689), .A2(new_n686), .A3(new_n961), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT45), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n684), .ZN(new_n985));
  INV_X1    g0785(.A(new_n688), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n689), .B1(new_n683), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n743), .B(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n988), .A2(new_n716), .A3(new_n740), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n678), .B(new_n683), .C1(new_n981), .C2(new_n983), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n985), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n978), .B1(new_n991), .B2(new_n741), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n746), .B(KEYINPUT103), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n976), .B(new_n977), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n804), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n691), .B2(new_n313), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n798), .A2(new_n240), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n747), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n367), .B1(new_n771), .B2(G77), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT104), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(KEYINPUT104), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n775), .A2(G68), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n836), .A2(new_n837), .B1(new_n201), .B2(new_n751), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G159), .A2(new_n762), .B1(new_n833), .B2(G50), .ZN(new_n1005));
  INV_X1    g0805(.A(G150), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n757), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1004), .B(new_n1007), .C1(G137), .C2(new_n778), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n367), .B1(new_n763), .B2(new_n790), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n757), .A2(new_n476), .B1(new_n836), .B2(new_n781), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G283), .C2(new_n833), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n778), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n751), .A2(new_n495), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1013), .A2(new_n1014), .B1(KEYINPUT46), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT46), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n771), .A2(G97), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n775), .A2(G107), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1012), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1009), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT47), .Z(new_n1022));
  OAI221_X1 g0822(.A(new_n999), .B1(new_n806), .B2(new_n953), .C1(new_n1022), .C2(new_n851), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n995), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT105), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT105), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n995), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(G387));
  NOR2_X1   g0829(.A1(new_n989), .A2(new_n697), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n988), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1030), .B1(new_n741), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n683), .A2(new_n806), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n747), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n795), .A2(new_n694), .B1(new_n532), .B2(new_n691), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT106), .Z(new_n1036));
  NOR2_X1   g0836(.A1(new_n317), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g0838(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n693), .A3(new_n1039), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n691), .B(new_n263), .C1(new_n237), .C2(G45), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1034), .B1(new_n1042), .B2(new_n996), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n752), .A2(G77), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n757), .B2(new_n286), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n263), .B1(new_n202), .B2(new_n759), .C1(new_n763), .C2(new_n282), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(G150), .C2(new_n778), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n775), .A2(new_n313), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n765), .A2(G159), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT107), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1047), .A2(new_n1018), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G311), .A2(new_n762), .B1(new_n833), .B2(G303), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n1014), .B2(new_n757), .C1(new_n785), .C2(new_n836), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n789), .B2(new_n776), .C1(new_n790), .C2(new_n751), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT49), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n263), .B1(new_n778), .B2(G326), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n770), .B2(new_n495), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1051), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1043), .B1(new_n1062), .B2(new_n793), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1031), .A2(new_n994), .B1(new_n1033), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1032), .A2(new_n1064), .ZN(G393));
  NAND3_X1  g0865(.A1(new_n985), .A2(KEYINPUT108), .A3(new_n990), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n984), .A2(KEYINPUT108), .A3(new_n684), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n692), .B(new_n991), .C1(new_n1068), .C2(new_n989), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G150), .A2(new_n765), .B1(new_n756), .B2(G159), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT109), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n263), .B1(new_n763), .B2(new_n286), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G68), .B2(new_n752), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n837), .B2(new_n1013), .C1(new_n317), .C2(new_n759), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n776), .A2(new_n268), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n1072), .A2(new_n841), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(KEYINPUT110), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT110), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n263), .B1(new_n752), .B2(G283), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n772), .B(new_n1081), .C1(new_n785), .C2(new_n1013), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT112), .Z(new_n1083));
  AOI22_X1  g0883(.A1(G311), .A2(new_n756), .B1(new_n765), .B2(G317), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1084), .A2(new_n1086), .B1(G116), .B2(new_n775), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G303), .A2(new_n762), .B1(new_n833), .B2(G294), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1080), .A2(new_n1077), .B1(new_n1083), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n793), .B1(new_n1079), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n798), .A2(new_n248), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n804), .B1(new_n221), .B2(new_n208), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1034), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n803), .B2(new_n973), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1068), .B2(new_n994), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1069), .A2(new_n1097), .ZN(G390));
  NAND4_X1  g0898(.A1(new_n738), .A2(G330), .A3(new_n818), .A4(new_n917), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n903), .B(KEYINPUT99), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n812), .B1(new_n711), .B2(new_n815), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n918), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1100), .B1(new_n1104), .B2(new_n929), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n905), .B1(new_n908), .B2(new_n917), .ZN(new_n1106));
  OAI211_X1 g0906(.A(KEYINPUT113), .B(new_n1105), .C1(new_n902), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT113), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n921), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT39), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n929), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1106), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n929), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1099), .B1(new_n1113), .B2(new_n1103), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1104), .A2(new_n929), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n902), .B2(new_n1106), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n933), .A2(G330), .A3(new_n818), .A4(new_n917), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1107), .A2(new_n1115), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n994), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n775), .A2(G159), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1122), .B1(new_n835), .B2(new_n763), .C1(new_n759), .C2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT116), .Z(new_n1125));
  NAND2_X1  g0925(.A1(new_n778), .A2(G125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n367), .B1(new_n756), .B2(G132), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n765), .A2(G128), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n751), .A2(new_n1006), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT53), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n286), .B2(new_n770), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1125), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G107), .A2(new_n762), .B1(new_n833), .B2(G97), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n789), .B2(new_n836), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT117), .Z(new_n1136));
  NAND2_X1  g0936(.A1(new_n778), .A2(G294), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n826), .A2(new_n367), .A3(new_n753), .A4(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n776), .A2(new_n268), .B1(new_n495), .B2(new_n757), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(KEYINPUT118), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(KEYINPUT118), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n793), .B1(new_n1133), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n747), .B1(new_n282), .B2(new_n824), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n902), .C2(new_n802), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1121), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n738), .A2(G330), .A3(new_n818), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n918), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1118), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n933), .A2(G330), .A3(new_n818), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n918), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n908), .A2(new_n1151), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n933), .A2(G330), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n472), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n925), .A2(new_n663), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT114), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n925), .A2(new_n663), .A3(new_n1157), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT114), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1154), .A2(new_n1102), .A3(new_n1099), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n917), .A2(new_n818), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1156), .A2(new_n1163), .B1(new_n1149), .B2(new_n918), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1164), .B2(new_n909), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1161), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1159), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1147), .A2(new_n1148), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT115), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1120), .A2(KEYINPUT115), .A3(new_n1167), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1120), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1167), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n697), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1146), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(G378));
  NAND2_X1  g0977(.A1(new_n296), .A2(new_n669), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT55), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n349), .B(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1183), .A2(new_n1184), .A3(KEYINPUT120), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT120), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1187), .A2(new_n802), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n263), .A2(G41), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n312), .B2(new_n759), .C1(new_n763), .C2(new_n221), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1044), .B1(new_n836), .B2(new_n495), .C1(new_n532), .C2(new_n757), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(G283), .C2(new_n778), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n771), .A2(G58), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1003), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1189), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n286), .C1(G33), .C2(G41), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n762), .A2(G132), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n835), .B2(new_n759), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G128), .B2(new_n756), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1123), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n752), .A2(new_n1203), .B1(new_n765), .B2(G125), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n1006), .C2(new_n776), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n771), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n778), .C2(G124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(new_n1195), .B2(new_n1194), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n793), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n747), .B1(new_n286), .B2(new_n824), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1188), .A2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(KEYINPUT40), .B(new_n934), .C1(new_n921), .C2(new_n887), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1187), .B(G330), .C1(new_n1216), .C2(new_n936), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n677), .B1(new_n937), .B2(new_n938), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT121), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n924), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1221), .B(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1223), .B2(new_n994), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT115), .B1(new_n1120), .B2(new_n1167), .ZN(new_n1225));
  AND4_X1   g1025(.A1(KEYINPUT115), .A2(new_n1147), .A3(new_n1148), .A4(new_n1167), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1160), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1223), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1158), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(KEYINPUT57), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n692), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1224), .B1(new_n1228), .B2(new_n1233), .ZN(G375));
  NAND2_X1  g1034(.A1(new_n918), .A2(new_n801), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n793), .A2(G68), .A3(new_n801), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n367), .B1(new_n532), .B2(new_n759), .C1(new_n763), .C2(new_n495), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G303), .B2(new_n778), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n771), .A2(G77), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n757), .A2(new_n789), .B1(new_n221), .B2(new_n751), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G294), .B2(new_n765), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1048), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n778), .A2(G128), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n263), .B1(new_n763), .B2(new_n1123), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G132), .B2(new_n765), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G159), .A2(new_n752), .B1(new_n756), .B2(G137), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1193), .A2(new_n1243), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n775), .A2(G50), .B1(G150), .B2(new_n833), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT122), .Z(new_n1249));
  OAI21_X1  g1049(.A(new_n1242), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n747), .B(new_n1236), .C1(new_n1250), .C2(new_n793), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1165), .A2(new_n994), .B1(new_n1235), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1174), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n1254), .B2(new_n978), .ZN(G381));
  INV_X1    g1055(.A(G375), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1032), .A2(new_n809), .A3(new_n1064), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(G390), .A2(new_n1257), .A3(G384), .A4(G381), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n1028), .A3(new_n1176), .A4(new_n1258), .ZN(G407));
  INV_X1    g1059(.A(G213), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(G343), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1176), .A2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(G375), .C2(new_n1262), .ZN(G409));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1024), .A2(new_n1069), .A3(new_n1097), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(G390), .A2(new_n995), .A3(new_n1023), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G393), .B(new_n809), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(G390), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1266), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1272), .A2(new_n995), .A3(new_n1023), .A4(G390), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1269), .A2(new_n1271), .A3(KEYINPUT125), .A4(new_n1273), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G378), .B(new_n1224), .C1(new_n1228), .C2(new_n1233), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n924), .B1(new_n1220), .B2(KEYINPUT121), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1229), .A2(new_n1283), .A3(new_n978), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1230), .A2(new_n994), .A3(new_n1231), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1188), .B2(new_n1214), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1176), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1261), .B1(new_n1280), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G384), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1253), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n692), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1254), .B2(KEYINPUT60), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1252), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1289), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1167), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(new_n1290), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G384), .B(new_n1252), .C1(new_n1297), .C2(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1261), .A2(KEYINPUT123), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1295), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1261), .A2(G2897), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1300), .B(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1279), .B1(new_n1288), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1304), .B1(new_n1288), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n1261), .B(new_n1305), .C1(new_n1280), .C2(new_n1287), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1304), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1278), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1306), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1312), .B(new_n1279), .C1(new_n1288), .C2(new_n1302), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1274), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1309), .B2(KEYINPUT63), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1264), .B1(new_n1311), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1288), .A2(new_n1306), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1274), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1303), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1312), .A3(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1323), .A2(new_n1303), .A3(new_n1307), .ZN(new_n1324));
  OAI211_X1 g1124(.A(KEYINPUT126), .B(new_n1322), .C1(new_n1324), .C2(new_n1278), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1317), .A2(new_n1325), .ZN(G405));
  NAND2_X1  g1126(.A1(G375), .A2(new_n1176), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1280), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1327), .A2(KEYINPUT127), .A3(new_n1280), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1306), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1330), .A2(new_n1305), .A3(new_n1331), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1278), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1335), .B(new_n1336), .ZN(G402));
endmodule


