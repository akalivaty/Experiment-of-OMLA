

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U546 ( .A1(G651), .A2(n576), .ZN(n791) );
  AND2_X1 U547 ( .A1(n745), .A2(n912), .ZN(n509) );
  OR2_X1 U548 ( .A1(n744), .A2(n743), .ZN(n510) );
  NOR2_X1 U549 ( .A1(n690), .A2(n961), .ZN(n639) );
  XNOR2_X1 U550 ( .A(KEYINPUT100), .B(KEYINPUT30), .ZN(n684) );
  XNOR2_X1 U551 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U552 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U553 ( .A1(G1966), .A2(n733), .ZN(n708) );
  NAND2_X1 U554 ( .A1(n625), .A2(n624), .ZN(n690) );
  NAND2_X1 U555 ( .A1(n792), .A2(G56), .ZN(n634) );
  NOR2_X2 U556 ( .A1(G2105), .A2(n515), .ZN(n872) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n517), .Z(n873) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n752) );
  NOR2_X1 U559 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U560 ( .A(G2105), .ZN(n516) );
  NOR2_X2 U561 ( .A1(n516), .A2(G2104), .ZN(n868) );
  NAND2_X1 U562 ( .A1(G126), .A2(n868), .ZN(n511) );
  XNOR2_X1 U563 ( .A(n511), .B(KEYINPUT88), .ZN(n514) );
  INV_X1 U564 ( .A(G2104), .ZN(n515) );
  NAND2_X1 U565 ( .A1(G102), .A2(n872), .ZN(n512) );
  XOR2_X1 U566 ( .A(KEYINPUT89), .B(n512), .Z(n513) );
  NAND2_X1 U567 ( .A1(n514), .A2(n513), .ZN(n521) );
  NOR2_X1 U568 ( .A1(n516), .A2(n515), .ZN(n869) );
  NAND2_X1 U569 ( .A1(G114), .A2(n869), .ZN(n519) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  NAND2_X1 U571 ( .A1(G138), .A2(n873), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U573 ( .A1(n521), .A2(n520), .ZN(G164) );
  NAND2_X1 U574 ( .A1(G101), .A2(n872), .ZN(n522) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(n522), .Z(n525) );
  NAND2_X1 U576 ( .A1(G125), .A2(n868), .ZN(n523) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n523), .Z(n524) );
  NAND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n873), .A2(G137), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n869), .A2(G113), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n576) );
  INV_X1 U583 ( .A(G651), .ZN(n530) );
  NOR2_X1 U584 ( .A1(n576), .A2(n530), .ZN(n786) );
  NAND2_X1 U585 ( .A1(n786), .A2(G72), .ZN(n533) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n531) );
  XNOR2_X1 U587 ( .A(n531), .B(KEYINPUT64), .ZN(n787) );
  NAND2_X1 U588 ( .A1(G85), .A2(n787), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n791), .A2(G47), .ZN(n537) );
  NOR2_X1 U591 ( .A1(G543), .A2(n530), .ZN(n534) );
  XOR2_X1 U592 ( .A(KEYINPUT66), .B(n534), .Z(n535) );
  XNOR2_X2 U593 ( .A(KEYINPUT1), .B(n535), .ZN(n792) );
  NAND2_X1 U594 ( .A1(G60), .A2(n792), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n537), .A2(n536), .ZN(n538) );
  OR2_X1 U596 ( .A1(n539), .A2(n538), .ZN(G290) );
  NAND2_X1 U597 ( .A1(G73), .A2(n786), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n540), .B(KEYINPUT2), .ZN(n547) );
  NAND2_X1 U599 ( .A1(n791), .A2(G48), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G86), .A2(n787), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n792), .A2(G61), .ZN(n543) );
  XOR2_X1 U603 ( .A(KEYINPUT82), .B(n543), .Z(n544) );
  NOR2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(G305) );
  NAND2_X1 U606 ( .A1(n791), .A2(G52), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G64), .A2(n792), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n786), .A2(G77), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT67), .B(n550), .Z(n552) );
  NAND2_X1 U611 ( .A1(G90), .A2(n787), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U614 ( .A1(n555), .A2(n554), .ZN(G171) );
  NAND2_X1 U615 ( .A1(G89), .A2(n787), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G76), .A2(n786), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n559), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G63), .A2(n792), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT76), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G51), .A2(n791), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U627 ( .A1(n786), .A2(G75), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G88), .A2(n787), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U630 ( .A(KEYINPUT84), .B(n569), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G62), .A2(n792), .ZN(n570) );
  XNOR2_X1 U632 ( .A(KEYINPUT83), .B(n570), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n791), .A2(G50), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(G303) );
  XNOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .ZN(n575) );
  XNOR2_X1 U637 ( .A(n575), .B(KEYINPUT77), .ZN(G286) );
  NAND2_X1 U638 ( .A1(G87), .A2(n576), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U641 ( .A1(n792), .A2(n579), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G49), .A2(n791), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT81), .B(n580), .Z(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(G288) );
  NOR2_X2 U645 ( .A1(G164), .A2(G1384), .ZN(n624) );
  NAND2_X1 U646 ( .A1(G160), .A2(G40), .ZN(n623) );
  NOR2_X1 U647 ( .A1(n624), .A2(n623), .ZN(n745) );
  NAND2_X1 U648 ( .A1(G117), .A2(n869), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G141), .A2(n873), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n872), .A2(G105), .ZN(n585) );
  XOR2_X1 U652 ( .A(KEYINPUT38), .B(n585), .Z(n586) );
  NOR2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n868), .A2(G129), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n880) );
  NOR2_X1 U656 ( .A1(n880), .A2(G1996), .ZN(n590) );
  XNOR2_X1 U657 ( .A(n590), .B(KEYINPUT104), .ZN(n994) );
  XNOR2_X1 U658 ( .A(n745), .B(KEYINPUT92), .ZN(n599) );
  NAND2_X1 U659 ( .A1(G1996), .A2(n880), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G107), .A2(n869), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G131), .A2(n873), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G119), .A2(n868), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G95), .A2(n872), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n882) );
  NAND2_X1 U667 ( .A1(G1991), .A2(n882), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n981) );
  NAND2_X1 U669 ( .A1(n599), .A2(n981), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT93), .ZN(n746) );
  NOR2_X1 U671 ( .A1(G1991), .A2(n882), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT105), .B(n601), .Z(n985) );
  NOR2_X1 U673 ( .A1(G1986), .A2(G290), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n985), .A2(n602), .ZN(n603) );
  NOR2_X1 U675 ( .A1(n746), .A2(n603), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n994), .A2(n604), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT39), .ZN(n617) );
  NAND2_X1 U678 ( .A1(G104), .A2(n872), .ZN(n607) );
  NAND2_X1 U679 ( .A1(G140), .A2(n873), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U681 ( .A(KEYINPUT34), .B(n608), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n869), .A2(G116), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT90), .ZN(n611) );
  NAND2_X1 U684 ( .A1(G128), .A2(n868), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U686 ( .A(n612), .B(KEYINPUT35), .Z(n613) );
  NOR2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U688 ( .A(KEYINPUT36), .B(n615), .Z(n616) );
  XNOR2_X1 U689 ( .A(KEYINPUT91), .B(n616), .ZN(n891) );
  XNOR2_X1 U690 ( .A(G2067), .B(KEYINPUT37), .ZN(n618) );
  NOR2_X1 U691 ( .A1(n891), .A2(n618), .ZN(n989) );
  NAND2_X1 U692 ( .A1(n989), .A2(n745), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n617), .A2(n622), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n891), .A2(n618), .ZN(n982) );
  NAND2_X1 U695 ( .A1(n619), .A2(n982), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n745), .A2(n620), .ZN(n621) );
  XOR2_X1 U697 ( .A(KEYINPUT106), .B(n621), .Z(n751) );
  INV_X1 U698 ( .A(n622), .ZN(n749) );
  INV_X1 U699 ( .A(n623), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G8), .A2(n690), .ZN(n733) );
  NOR2_X1 U701 ( .A1(G1981), .A2(G305), .ZN(n626) );
  XOR2_X1 U702 ( .A(n626), .B(KEYINPUT24), .Z(n627) );
  NOR2_X1 U703 ( .A1(n733), .A2(n627), .ZN(n744) );
  NAND2_X1 U704 ( .A1(G81), .A2(n787), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT12), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G68), .A2(n786), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n631), .B(KEYINPUT13), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G43), .A2(n791), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n636) );
  XOR2_X1 U711 ( .A(n634), .B(KEYINPUT14), .Z(n635) );
  NOR2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X2 U713 ( .A(KEYINPUT72), .B(n637), .Z(n919) );
  XOR2_X1 U714 ( .A(KEYINPUT96), .B(G1996), .Z(n961) );
  XNOR2_X1 U715 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n638) );
  XNOR2_X1 U716 ( .A(n639), .B(n638), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n690), .A2(G1341), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U719 ( .A1(n919), .A2(n642), .ZN(n657) );
  NAND2_X1 U720 ( .A1(G92), .A2(n787), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G66), .A2(n792), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U723 ( .A(KEYINPUT74), .B(n645), .ZN(n649) );
  NAND2_X1 U724 ( .A1(G79), .A2(n786), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G54), .A2(n791), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U728 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(n904) );
  NAND2_X1 U730 ( .A1(n657), .A2(n904), .ZN(n655) );
  NOR2_X1 U731 ( .A1(G2067), .A2(n690), .ZN(n653) );
  INV_X1 U732 ( .A(n690), .ZN(n678) );
  NOR2_X1 U733 ( .A1(n678), .A2(G1348), .ZN(n652) );
  NOR2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT98), .ZN(n659) );
  OR2_X1 U737 ( .A1(n904), .A2(n657), .ZN(n658) );
  AND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n791), .A2(G53), .ZN(n661) );
  NAND2_X1 U740 ( .A1(G91), .A2(n787), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n786), .A2(G78), .ZN(n662) );
  XOR2_X1 U743 ( .A(KEYINPUT68), .B(n662), .Z(n663) );
  NOR2_X1 U744 ( .A1(n664), .A2(n663), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G65), .A2(n792), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n910) );
  NAND2_X1 U747 ( .A1(n678), .A2(G2072), .ZN(n667) );
  XOR2_X1 U748 ( .A(KEYINPUT27), .B(n667), .Z(n669) );
  XOR2_X1 U749 ( .A(G1956), .B(KEYINPUT95), .Z(n937) );
  NAND2_X1 U750 ( .A1(n937), .A2(n690), .ZN(n668) );
  NAND2_X1 U751 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U752 ( .A1(n910), .A2(n673), .ZN(n670) );
  NOR2_X1 U753 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U754 ( .A(KEYINPUT99), .B(n672), .ZN(n676) );
  AND2_X1 U755 ( .A1(n910), .A2(n673), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT28), .B(n674), .Z(n675) );
  AND2_X1 U757 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U758 ( .A(n677), .B(KEYINPUT29), .ZN(n706) );
  OR2_X1 U759 ( .A1(n678), .A2(G1961), .ZN(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT25), .B(G2078), .ZN(n970) );
  NAND2_X1 U761 ( .A1(n678), .A2(n970), .ZN(n679) );
  NAND2_X1 U762 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G171), .A2(n682), .ZN(n681) );
  XNOR2_X1 U764 ( .A(KEYINPUT94), .B(n681), .ZN(n704) );
  NAND2_X1 U765 ( .A1(n706), .A2(n704), .ZN(n695) );
  NOR2_X1 U766 ( .A1(G171), .A2(n682), .ZN(n688) );
  NOR2_X1 U767 ( .A1(G2084), .A2(n690), .ZN(n711) );
  NOR2_X1 U768 ( .A1(n708), .A2(n711), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G8), .A2(n683), .ZN(n685) );
  NOR2_X1 U770 ( .A1(G168), .A2(n686), .ZN(n687) );
  XOR2_X1 U771 ( .A(KEYINPUT31), .B(n689), .Z(n707) );
  NOR2_X1 U772 ( .A1(G1971), .A2(n733), .ZN(n692) );
  NOR2_X1 U773 ( .A1(G2090), .A2(n690), .ZN(n691) );
  NOR2_X1 U774 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U775 ( .A1(n693), .A2(G303), .ZN(n696) );
  AND2_X1 U776 ( .A1(n707), .A2(n696), .ZN(n694) );
  NAND2_X1 U777 ( .A1(n695), .A2(n694), .ZN(n700) );
  INV_X1 U778 ( .A(n696), .ZN(n697) );
  OR2_X1 U779 ( .A1(n697), .A2(G286), .ZN(n698) );
  AND2_X1 U780 ( .A1(G8), .A2(n698), .ZN(n699) );
  NAND2_X1 U781 ( .A1(n700), .A2(n699), .ZN(n702) );
  XOR2_X1 U782 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n701) );
  XNOR2_X1 U783 ( .A(n702), .B(n701), .ZN(n721) );
  INV_X1 U784 ( .A(n708), .ZN(n703) );
  AND2_X1 U785 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U786 ( .A1(n706), .A2(n705), .ZN(n710) );
  OR2_X1 U787 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U788 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U789 ( .A1(G8), .A2(n711), .ZN(n712) );
  NAND2_X1 U790 ( .A1(n713), .A2(n712), .ZN(n723) );
  NAND2_X1 U791 ( .A1(n721), .A2(n723), .ZN(n716) );
  NOR2_X1 U792 ( .A1(G2090), .A2(G303), .ZN(n714) );
  NAND2_X1 U793 ( .A1(G8), .A2(n714), .ZN(n715) );
  NAND2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n718) );
  INV_X1 U795 ( .A(KEYINPUT103), .ZN(n717) );
  XNOR2_X1 U796 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U797 ( .A1(n719), .A2(n733), .ZN(n742) );
  NAND2_X1 U798 ( .A1(G288), .A2(G1976), .ZN(n720) );
  XNOR2_X1 U799 ( .A(n720), .B(KEYINPUT102), .ZN(n909) );
  AND2_X1 U800 ( .A1(n721), .A2(n909), .ZN(n728) );
  INV_X1 U801 ( .A(n733), .ZN(n722) );
  AND2_X1 U802 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U803 ( .A1(G1976), .A2(G288), .ZN(n907) );
  NAND2_X1 U804 ( .A1(n907), .A2(KEYINPUT33), .ZN(n724) );
  NOR2_X1 U805 ( .A1(n724), .A2(n733), .ZN(n737) );
  INV_X1 U806 ( .A(n737), .ZN(n725) );
  AND2_X1 U807 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U808 ( .A1(n728), .A2(n727), .ZN(n739) );
  INV_X1 U809 ( .A(KEYINPUT33), .ZN(n735) );
  INV_X1 U810 ( .A(n909), .ZN(n731) );
  NOR2_X1 U811 ( .A1(G1971), .A2(G303), .ZN(n729) );
  NOR2_X1 U812 ( .A1(n907), .A2(n729), .ZN(n730) );
  OR2_X1 U813 ( .A1(n731), .A2(n730), .ZN(n732) );
  OR2_X1 U814 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U815 ( .A1(n735), .A2(n734), .ZN(n736) );
  OR2_X1 U816 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U817 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U818 ( .A(G1981), .B(G305), .Z(n921) );
  NAND2_X1 U819 ( .A1(n740), .A2(n921), .ZN(n741) );
  NAND2_X1 U820 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U821 ( .A(G1986), .B(G290), .ZN(n912) );
  NOR2_X1 U822 ( .A1(n746), .A2(n509), .ZN(n747) );
  NAND2_X1 U823 ( .A1(n510), .A2(n747), .ZN(n748) );
  NOR2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U826 ( .A(n753), .B(n752), .ZN(G329) );
  XOR2_X1 U827 ( .A(G2443), .B(G2446), .Z(n755) );
  XNOR2_X1 U828 ( .A(G2427), .B(G2451), .ZN(n754) );
  XNOR2_X1 U829 ( .A(n755), .B(n754), .ZN(n761) );
  XOR2_X1 U830 ( .A(G2430), .B(G2454), .Z(n757) );
  XNOR2_X1 U831 ( .A(G1341), .B(G1348), .ZN(n756) );
  XNOR2_X1 U832 ( .A(n757), .B(n756), .ZN(n759) );
  XOR2_X1 U833 ( .A(G2435), .B(G2438), .Z(n758) );
  XNOR2_X1 U834 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U835 ( .A(n761), .B(n760), .Z(n762) );
  AND2_X1 U836 ( .A1(G14), .A2(n762), .ZN(G401) );
  AND2_X1 U837 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U838 ( .A(G860), .ZN(n770) );
  OR2_X1 U839 ( .A1(n770), .A2(n919), .ZN(G153) );
  INV_X1 U840 ( .A(G57), .ZN(G237) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  XOR2_X1 U842 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n764) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n763) );
  XNOR2_X1 U844 ( .A(n764), .B(n763), .ZN(G223) );
  INV_X1 U845 ( .A(G223), .ZN(n826) );
  NAND2_X1 U846 ( .A1(n826), .A2(G567), .ZN(n765) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n765), .Z(G234) );
  XNOR2_X1 U848 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U849 ( .A1(G868), .A2(G301), .ZN(n767) );
  OR2_X1 U850 ( .A1(n904), .A2(G868), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n767), .A2(n766), .ZN(G284) );
  XOR2_X1 U852 ( .A(n910), .B(KEYINPUT69), .Z(G299) );
  NAND2_X1 U853 ( .A1(G286), .A2(G868), .ZN(n769) );
  INV_X1 U854 ( .A(G868), .ZN(n807) );
  NAND2_X1 U855 ( .A1(G299), .A2(n807), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n770), .A2(G559), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n771), .A2(n904), .ZN(n772) );
  XNOR2_X1 U859 ( .A(n772), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U860 ( .A1(n904), .A2(G868), .ZN(n773) );
  XNOR2_X1 U861 ( .A(KEYINPUT78), .B(n773), .ZN(n774) );
  NOR2_X1 U862 ( .A1(G559), .A2(n774), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n919), .A2(G868), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(G282) );
  NAND2_X1 U865 ( .A1(G111), .A2(n869), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G135), .A2(n873), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n868), .A2(G123), .ZN(n779) );
  XOR2_X1 U869 ( .A(KEYINPUT18), .B(n779), .Z(n780) );
  NOR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n872), .A2(G99), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n986) );
  XOR2_X1 U873 ( .A(n986), .B(G2096), .Z(n785) );
  XNOR2_X1 U874 ( .A(G2100), .B(KEYINPUT79), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(G156) );
  NAND2_X1 U876 ( .A1(n786), .A2(G80), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G93), .A2(n787), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U879 ( .A(KEYINPUT80), .B(n790), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n791), .A2(G55), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G67), .A2(n792), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n808) );
  NAND2_X1 U884 ( .A1(n904), .A2(G559), .ZN(n805) );
  XNOR2_X1 U885 ( .A(n919), .B(n805), .ZN(n797) );
  NOR2_X1 U886 ( .A1(G860), .A2(n797), .ZN(n798) );
  XOR2_X1 U887 ( .A(n808), .B(n798), .Z(G145) );
  INV_X1 U888 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U889 ( .A(KEYINPUT19), .B(G288), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n799), .B(G299), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n800), .B(n808), .ZN(n802) );
  XNOR2_X1 U892 ( .A(n919), .B(G166), .ZN(n801) );
  XNOR2_X1 U893 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U894 ( .A(n803), .B(G305), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n804), .B(G290), .ZN(n894) );
  XNOR2_X1 U896 ( .A(n894), .B(n805), .ZN(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n810) );
  NOR2_X1 U898 ( .A1(G868), .A2(n808), .ZN(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XNOR2_X1 U901 ( .A(n811), .B(KEYINPUT85), .ZN(n812) );
  XNOR2_X1 U902 ( .A(n812), .B(KEYINPUT20), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(G2090), .ZN(n814) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U907 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U910 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U911 ( .A1(G96), .A2(n818), .ZN(n832) );
  NAND2_X1 U912 ( .A1(n832), .A2(G2106), .ZN(n823) );
  NAND2_X1 U913 ( .A1(G120), .A2(G108), .ZN(n819) );
  NOR2_X1 U914 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(G69), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n821), .B(KEYINPUT86), .ZN(n831) );
  NAND2_X1 U917 ( .A1(n831), .A2(G567), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n834) );
  NAND2_X1 U919 ( .A1(G483), .A2(G661), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n834), .A2(n824), .ZN(n825) );
  XOR2_X1 U921 ( .A(KEYINPUT87), .B(n825), .Z(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n826), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n827) );
  XOR2_X1 U925 ( .A(KEYINPUT108), .B(n827), .Z(n828) );
  NAND2_X1 U926 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U928 ( .A1(n830), .A2(n829), .ZN(G188) );
  XOR2_X1 U929 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n833), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U935 ( .A(G261), .ZN(G325) );
  INV_X1 U936 ( .A(n834), .ZN(G319) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n836) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n838) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U942 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U943 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1986), .B(G1976), .Z(n844) );
  XNOR2_X1 U947 ( .A(G1956), .B(G1971), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U949 ( .A(n845), .B(G2474), .Z(n847) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1981), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U952 ( .A(KEYINPUT41), .B(G1991), .Z(n849) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1961), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U955 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G112), .A2(n869), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n852), .B(KEYINPUT110), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G124), .A2(n868), .ZN(n853) );
  XNOR2_X1 U959 ( .A(n853), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U960 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G100), .A2(n872), .ZN(n857) );
  NAND2_X1 U962 ( .A1(G136), .A2(n873), .ZN(n856) );
  NAND2_X1 U963 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U964 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G103), .A2(n872), .ZN(n861) );
  NAND2_X1 U966 ( .A1(G139), .A2(n873), .ZN(n860) );
  NAND2_X1 U967 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n869), .A2(G115), .ZN(n862) );
  XNOR2_X1 U969 ( .A(n862), .B(KEYINPUT112), .ZN(n864) );
  NAND2_X1 U970 ( .A1(G127), .A2(n868), .ZN(n863) );
  NAND2_X1 U971 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U972 ( .A(KEYINPUT47), .B(n865), .Z(n866) );
  NOR2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n997) );
  NAND2_X1 U974 ( .A1(G130), .A2(n868), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G118), .A2(n869), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G106), .A2(n872), .ZN(n875) );
  NAND2_X1 U978 ( .A1(G142), .A2(n873), .ZN(n874) );
  NAND2_X1 U979 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  NOR2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n997), .B(n879), .ZN(n890) );
  XNOR2_X1 U983 ( .A(G162), .B(n880), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n881), .B(n986), .ZN(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n882), .B(KEYINPUT111), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U988 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U989 ( .A(G160), .B(G164), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n892) );
  XOR2_X1 U992 ( .A(n892), .B(n891), .Z(n893) );
  NOR2_X1 U993 ( .A1(G37), .A2(n893), .ZN(G395) );
  XOR2_X1 U994 ( .A(n894), .B(G286), .Z(n896) );
  XNOR2_X1 U995 ( .A(n904), .B(G171), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U997 ( .A1(G37), .A2(n897), .ZN(G397) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n898), .B(KEYINPUT49), .ZN(n899) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n899), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n900), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(KEYINPUT113), .B(n901), .ZN(n903) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n902) );
  NAND2_X1 U1004 ( .A1(n903), .A2(n902), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1007 ( .A(G171), .B(G1961), .Z(n906) );
  XOR2_X1 U1008 ( .A(n904), .B(G1348), .Z(n905) );
  NOR2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n918) );
  XOR2_X1 U1010 ( .A(n907), .B(KEYINPUT120), .Z(n908) );
  NAND2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(G166), .B(G1971), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(G1956), .B(n910), .ZN(n911) );
  NOR2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n927) );
  XNOR2_X1 U1018 ( .A(G1341), .B(n919), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n920), .B(KEYINPUT121), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(G1966), .B(G168), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n923), .B(KEYINPUT57), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1025 ( .A(KEYINPUT122), .B(n928), .Z(n930) );
  XNOR2_X1 U1026 ( .A(KEYINPUT56), .B(G16), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n1012) );
  XNOR2_X1 U1028 ( .A(G5), .B(G1961), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(KEYINPUT123), .ZN(n945) );
  XNOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(G4), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G20), .B(n937), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT124), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1039 ( .A(KEYINPUT60), .B(n941), .Z(n943) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n954) );
  XOR2_X1 U1043 ( .A(G1971), .B(G22), .Z(n948) );
  XOR2_X1 U1044 ( .A(G24), .B(KEYINPUT126), .Z(n946) );
  XNOR2_X1 U1045 ( .A(n946), .B(G1986), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1047 ( .A(KEYINPUT125), .B(G1976), .Z(n949) );
  XNOR2_X1 U1048 ( .A(G23), .B(n949), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1050 ( .A(KEYINPUT58), .B(n952), .Z(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(KEYINPUT61), .B(n955), .ZN(n957) );
  INV_X1 U1053 ( .A(G16), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n958), .A2(G11), .ZN(n1010) );
  XOR2_X1 U1056 ( .A(KEYINPUT118), .B(G34), .Z(n960) );
  XNOR2_X1 U1057 ( .A(G2084), .B(KEYINPUT54), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(n960), .B(n959), .ZN(n977) );
  XNOR2_X1 U1059 ( .A(G2090), .B(G35), .ZN(n975) );
  XNOR2_X1 U1060 ( .A(n961), .B(G32), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G26), .ZN(n963) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n962) );
  NOR2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1064 ( .A1(G28), .A2(n964), .ZN(n967) );
  XOR2_X1 U1065 ( .A(G25), .B(G1991), .Z(n965) );
  XNOR2_X1 U1066 ( .A(KEYINPUT117), .B(n965), .ZN(n966) );
  NOR2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1069 ( .A(G27), .B(n970), .Z(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(KEYINPUT119), .B(n978), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(G29), .A2(n979), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(n980), .B(KEYINPUT55), .ZN(n1008) );
  INV_X1 U1077 ( .A(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n992) );
  XOR2_X1 U1079 ( .A(G2084), .B(G160), .Z(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(KEYINPUT115), .B(n990), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n1004) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n995), .Z(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT116), .B(n996), .Z(n1002) );
  XOR2_X1 U1089 ( .A(G2072), .B(n997), .Z(n999) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1000), .Z(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT52), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(G29), .A2(n1006), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1013), .Z(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

