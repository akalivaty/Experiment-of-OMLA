

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(G2105), .A2(n531), .ZN(n896) );
  AND2_X1 U558 ( .A1(n742), .A2(n741), .ZN(n525) );
  AND2_X1 U559 ( .A1(n746), .A2(n724), .ZN(n725) );
  INV_X1 U560 ( .A(G8), .ZN(n704) );
  OR2_X1 U561 ( .A1(n766), .A2(n704), .ZN(n705) );
  NOR2_X1 U562 ( .A1(n765), .A2(n764), .ZN(n768) );
  INV_X1 U563 ( .A(KEYINPUT102), .ZN(n788) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  OR2_X1 U565 ( .A1(n698), .A2(n697), .ZN(n792) );
  INV_X1 U566 ( .A(KEYINPUT87), .ZN(n527) );
  NOR2_X1 U567 ( .A1(G651), .A2(n657), .ZN(n665) );
  XNOR2_X1 U568 ( .A(n528), .B(n527), .ZN(n529) );
  NOR2_X1 U569 ( .A1(n535), .A2(n534), .ZN(G164) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U571 ( .A1(n891), .A2(G114), .ZN(n530) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n526), .Z(n895) );
  NAND2_X1 U573 ( .A1(n895), .A2(G138), .ZN(n528) );
  NAND2_X1 U574 ( .A1(n530), .A2(n529), .ZN(n535) );
  INV_X1 U575 ( .A(G2104), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G102), .A2(n896), .ZN(n533) );
  AND2_X1 U577 ( .A1(n531), .A2(G2105), .ZN(n892) );
  NAND2_X1 U578 ( .A1(G126), .A2(n892), .ZN(n532) );
  NAND2_X1 U579 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U580 ( .A(G2427), .B(G2435), .Z(n537) );
  XNOR2_X1 U581 ( .A(G2454), .B(G2443), .ZN(n536) );
  XNOR2_X1 U582 ( .A(n537), .B(n536), .ZN(n544) );
  XOR2_X1 U583 ( .A(G2451), .B(KEYINPUT105), .Z(n539) );
  XNOR2_X1 U584 ( .A(G2430), .B(G2438), .ZN(n538) );
  XNOR2_X1 U585 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U586 ( .A(n540), .B(G2446), .Z(n542) );
  XNOR2_X1 U587 ( .A(G1341), .B(G1348), .ZN(n541) );
  XNOR2_X1 U588 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U589 ( .A(n544), .B(n543), .ZN(n545) );
  AND2_X1 U590 ( .A1(n545), .A2(G14), .ZN(G401) );
  AND2_X1 U591 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U592 ( .A1(G123), .A2(n892), .ZN(n546) );
  XNOR2_X1 U593 ( .A(n546), .B(KEYINPUT18), .ZN(n553) );
  NAND2_X1 U594 ( .A1(G135), .A2(n895), .ZN(n548) );
  NAND2_X1 U595 ( .A1(G111), .A2(n891), .ZN(n547) );
  NAND2_X1 U596 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U597 ( .A1(G99), .A2(n896), .ZN(n549) );
  XNOR2_X1 U598 ( .A(KEYINPUT77), .B(n549), .ZN(n550) );
  NOR2_X1 U599 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U600 ( .A1(n553), .A2(n552), .ZN(n977) );
  XNOR2_X1 U601 ( .A(G2096), .B(n977), .ZN(n554) );
  OR2_X1 U602 ( .A1(G2100), .A2(n554), .ZN(G156) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  XOR2_X1 U606 ( .A(KEYINPUT0), .B(G543), .Z(n657) );
  NAND2_X1 U607 ( .A1(n665), .A2(G52), .ZN(n558) );
  INV_X1 U608 ( .A(G651), .ZN(n559) );
  NOR2_X1 U609 ( .A1(G543), .A2(n559), .ZN(n555) );
  XOR2_X1 U610 ( .A(KEYINPUT1), .B(n555), .Z(n556) );
  XNOR2_X1 U611 ( .A(KEYINPUT66), .B(n556), .ZN(n666) );
  NAND2_X1 U612 ( .A1(G64), .A2(n666), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n564) );
  NOR2_X1 U614 ( .A1(G651), .A2(G543), .ZN(n661) );
  NAND2_X1 U615 ( .A1(G90), .A2(n661), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n657), .A2(n559), .ZN(n662) );
  NAND2_X1 U617 ( .A1(G77), .A2(n662), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U621 ( .A(KEYINPUT67), .B(n565), .Z(G171) );
  NAND2_X1 U622 ( .A1(G137), .A2(n895), .ZN(n566) );
  XOR2_X1 U623 ( .A(n566), .B(KEYINPUT65), .Z(n570) );
  XOR2_X1 U624 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n568) );
  NAND2_X1 U625 ( .A1(G101), .A2(n896), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n568), .B(n567), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n698) );
  NAND2_X1 U628 ( .A1(G113), .A2(n891), .ZN(n572) );
  NAND2_X1 U629 ( .A1(G125), .A2(n892), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n696) );
  NOR2_X1 U631 ( .A1(n698), .A2(n696), .ZN(G160) );
  NAND2_X1 U632 ( .A1(G78), .A2(n662), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT68), .ZN(n580) );
  NAND2_X1 U634 ( .A1(n661), .A2(G91), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G65), .A2(n666), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G53), .A2(n665), .ZN(n576) );
  XNOR2_X1 U638 ( .A(KEYINPUT69), .B(n576), .ZN(n577) );
  NOR2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(G299) );
  NAND2_X1 U641 ( .A1(G89), .A2(n661), .ZN(n581) );
  XNOR2_X1 U642 ( .A(n581), .B(KEYINPUT4), .ZN(n582) );
  XNOR2_X1 U643 ( .A(n582), .B(KEYINPUT72), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G76), .A2(n662), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U646 ( .A(KEYINPUT5), .B(n585), .ZN(n592) );
  XNOR2_X1 U647 ( .A(KEYINPUT6), .B(KEYINPUT74), .ZN(n590) );
  NAND2_X1 U648 ( .A1(G63), .A2(n666), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n665), .A2(G51), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT73), .B(n586), .Z(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U652 ( .A(n590), .B(n589), .Z(n591) );
  NAND2_X1 U653 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U654 ( .A(KEYINPUT7), .B(n593), .ZN(G168) );
  XOR2_X1 U655 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n594) );
  XNOR2_X1 U657 ( .A(n594), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U658 ( .A(G223), .ZN(n843) );
  NAND2_X1 U659 ( .A1(n843), .A2(G567), .ZN(n595) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n595), .Z(G234) );
  XOR2_X1 U661 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n597) );
  NAND2_X1 U662 ( .A1(G56), .A2(n666), .ZN(n596) );
  XNOR2_X1 U663 ( .A(n597), .B(n596), .ZN(n604) );
  NAND2_X1 U664 ( .A1(G81), .A2(n661), .ZN(n598) );
  XOR2_X1 U665 ( .A(KEYINPUT12), .B(n598), .Z(n599) );
  XNOR2_X1 U666 ( .A(n599), .B(KEYINPUT71), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G68), .A2(n662), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U669 ( .A(KEYINPUT13), .B(n602), .Z(n603) );
  NOR2_X1 U670 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U671 ( .A1(n665), .A2(G43), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n606), .A2(n605), .ZN(n920) );
  INV_X1 U673 ( .A(G860), .ZN(n619) );
  OR2_X1 U674 ( .A1(n920), .A2(n619), .ZN(G153) );
  INV_X1 U675 ( .A(G171), .ZN(G301) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n615) );
  NAND2_X1 U677 ( .A1(G79), .A2(n662), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G54), .A2(n665), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n661), .A2(G92), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G66), .A2(n666), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n613), .B(KEYINPUT15), .ZN(n928) );
  INV_X1 U685 ( .A(n928), .ZN(n908) );
  OR2_X1 U686 ( .A1(n908), .A2(G868), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(G284) );
  XNOR2_X1 U688 ( .A(KEYINPUT75), .B(G868), .ZN(n616) );
  NOR2_X1 U689 ( .A1(G286), .A2(n616), .ZN(n618) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(G297) );
  NAND2_X1 U692 ( .A1(G559), .A2(n619), .ZN(n620) );
  XNOR2_X1 U693 ( .A(KEYINPUT76), .B(n620), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n621), .A2(n908), .ZN(n622) );
  XNOR2_X1 U695 ( .A(KEYINPUT16), .B(n622), .ZN(G148) );
  NOR2_X1 U696 ( .A1(G868), .A2(n920), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G868), .A2(n908), .ZN(n623) );
  NOR2_X1 U698 ( .A1(G559), .A2(n623), .ZN(n624) );
  NOR2_X1 U699 ( .A1(n625), .A2(n624), .ZN(G282) );
  NAND2_X1 U700 ( .A1(G559), .A2(n908), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(n920), .ZN(n677) );
  XNOR2_X1 U702 ( .A(KEYINPUT78), .B(n677), .ZN(n627) );
  NOR2_X1 U703 ( .A1(G860), .A2(n627), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT83), .ZN(n639) );
  NAND2_X1 U705 ( .A1(G55), .A2(n665), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(KEYINPUT82), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n662), .A2(G80), .ZN(n630) );
  XOR2_X1 U708 ( .A(KEYINPUT79), .B(n630), .Z(n632) );
  NAND2_X1 U709 ( .A1(n661), .A2(G93), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U711 ( .A(KEYINPUT80), .B(n633), .Z(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G67), .A2(n666), .ZN(n636) );
  XNOR2_X1 U714 ( .A(KEYINPUT81), .B(n636), .ZN(n637) );
  NOR2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n679) );
  XOR2_X1 U716 ( .A(n639), .B(n679), .Z(G145) );
  NAND2_X1 U717 ( .A1(n661), .A2(G86), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G61), .A2(n666), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n662), .A2(G73), .ZN(n642) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n665), .A2(G48), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(G305) );
  AND2_X1 U725 ( .A1(G60), .A2(n666), .ZN(n650) );
  NAND2_X1 U726 ( .A1(G85), .A2(n661), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G72), .A2(n662), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n665), .A2(G47), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n652), .A2(n651), .ZN(G290) );
  NAND2_X1 U732 ( .A1(G49), .A2(n665), .ZN(n654) );
  NAND2_X1 U733 ( .A1(G74), .A2(G651), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U735 ( .A1(n666), .A2(n655), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT84), .ZN(n659) );
  NAND2_X1 U737 ( .A1(G87), .A2(n657), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U739 ( .A(KEYINPUT85), .B(n660), .Z(G288) );
  NAND2_X1 U740 ( .A1(G88), .A2(n661), .ZN(n664) );
  NAND2_X1 U741 ( .A1(G75), .A2(n662), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n665), .A2(G50), .ZN(n668) );
  NAND2_X1 U744 ( .A1(G62), .A2(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U746 ( .A1(n670), .A2(n669), .ZN(G166) );
  XOR2_X1 U747 ( .A(G290), .B(G288), .Z(n671) );
  XNOR2_X1 U748 ( .A(G305), .B(n671), .ZN(n674) );
  XOR2_X1 U749 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n672) );
  XNOR2_X1 U750 ( .A(G299), .B(n672), .ZN(n673) );
  XOR2_X1 U751 ( .A(n674), .B(n673), .Z(n676) );
  XNOR2_X1 U752 ( .A(G166), .B(n679), .ZN(n675) );
  XNOR2_X1 U753 ( .A(n676), .B(n675), .ZN(n912) );
  XNOR2_X1 U754 ( .A(n677), .B(n912), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n678), .A2(G868), .ZN(n681) );
  OR2_X1 U756 ( .A1(G868), .A2(n679), .ZN(n680) );
  NAND2_X1 U757 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U762 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U766 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U767 ( .A1(G96), .A2(n688), .ZN(n847) );
  NAND2_X1 U768 ( .A1(n847), .A2(G2106), .ZN(n692) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n689) );
  NOR2_X1 U770 ( .A1(G237), .A2(n689), .ZN(n690) );
  NAND2_X1 U771 ( .A1(G108), .A2(n690), .ZN(n848) );
  NAND2_X1 U772 ( .A1(n848), .A2(G567), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n692), .A2(n691), .ZN(n849) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U775 ( .A1(n849), .A2(n693), .ZN(n846) );
  NAND2_X1 U776 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  NOR2_X1 U778 ( .A1(G288), .A2(G1976), .ZN(n694) );
  XNOR2_X1 U779 ( .A(n694), .B(KEYINPUT100), .ZN(n921) );
  INV_X1 U780 ( .A(G40), .ZN(n695) );
  OR2_X1 U781 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U782 ( .A(n792), .B(KEYINPUT91), .ZN(n699) );
  NOR2_X1 U783 ( .A1(G164), .A2(G1384), .ZN(n793) );
  NAND2_X2 U784 ( .A1(n699), .A2(n793), .ZN(n731) );
  NAND2_X1 U785 ( .A1(G8), .A2(n731), .ZN(n700) );
  XOR2_X1 U786 ( .A(KEYINPUT92), .B(n700), .Z(n779) );
  NAND2_X1 U787 ( .A1(n921), .A2(n779), .ZN(n703) );
  XNOR2_X1 U788 ( .A(KEYINPUT101), .B(G1981), .ZN(n701) );
  XNOR2_X1 U789 ( .A(n701), .B(G305), .ZN(n940) );
  AND2_X1 U790 ( .A1(n940), .A2(KEYINPUT33), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n782) );
  INV_X1 U792 ( .A(n779), .ZN(n787) );
  NOR2_X1 U793 ( .A1(n787), .A2(G1966), .ZN(n765) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n731), .ZN(n766) );
  OR2_X1 U795 ( .A1(n765), .A2(n705), .ZN(n706) );
  XNOR2_X1 U796 ( .A(KEYINPUT30), .B(n706), .ZN(n707) );
  NOR2_X1 U797 ( .A1(G168), .A2(n707), .ZN(n711) );
  INV_X1 U798 ( .A(G1961), .ZN(n1019) );
  NAND2_X1 U799 ( .A1(n1019), .A2(n731), .ZN(n709) );
  XOR2_X1 U800 ( .A(KEYINPUT93), .B(n731), .Z(n722) );
  INV_X1 U801 ( .A(n722), .ZN(n727) );
  XNOR2_X1 U802 ( .A(KEYINPUT25), .B(G2078), .ZN(n955) );
  NAND2_X1 U803 ( .A1(n727), .A2(n955), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n753) );
  NOR2_X1 U805 ( .A1(G171), .A2(n753), .ZN(n710) );
  NOR2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U807 ( .A(KEYINPUT31), .B(n712), .Z(n762) );
  NOR2_X1 U808 ( .A1(G2090), .A2(n731), .ZN(n714) );
  NOR2_X1 U809 ( .A1(n787), .A2(G1971), .ZN(n713) );
  NOR2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U811 ( .A(KEYINPUT99), .B(n715), .Z(n716) );
  NAND2_X1 U812 ( .A1(n716), .A2(G303), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n762), .A2(n717), .ZN(n719) );
  INV_X1 U814 ( .A(n717), .ZN(n718) );
  OR2_X1 U815 ( .A1(n718), .A2(G286), .ZN(n754) );
  NAND2_X1 U816 ( .A1(n719), .A2(n754), .ZN(n757) );
  INV_X1 U817 ( .A(KEYINPUT27), .ZN(n721) );
  NAND2_X1 U818 ( .A1(n727), .A2(G2072), .ZN(n720) );
  XNOR2_X1 U819 ( .A(n721), .B(n720), .ZN(n746) );
  NAND2_X1 U820 ( .A1(G1956), .A2(n722), .ZN(n745) );
  INV_X1 U821 ( .A(n745), .ZN(n723) );
  NOR2_X1 U822 ( .A1(G299), .A2(n723), .ZN(n724) );
  XNOR2_X1 U823 ( .A(n725), .B(KEYINPUT96), .ZN(n726) );
  INV_X1 U824 ( .A(n726), .ZN(n743) );
  NAND2_X1 U825 ( .A1(n731), .A2(G1348), .ZN(n739) );
  NAND2_X1 U826 ( .A1(G2067), .A2(n727), .ZN(n728) );
  XNOR2_X1 U827 ( .A(n728), .B(KEYINPUT95), .ZN(n737) );
  INV_X1 U828 ( .A(n731), .ZN(n729) );
  NAND2_X1 U829 ( .A1(G1996), .A2(n729), .ZN(n730) );
  XNOR2_X1 U830 ( .A(KEYINPUT26), .B(n730), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n731), .A2(G1341), .ZN(n732) );
  XOR2_X1 U832 ( .A(KEYINPUT94), .B(n732), .Z(n733) );
  NOR2_X1 U833 ( .A1(n920), .A2(n733), .ZN(n734) );
  NAND2_X1 U834 ( .A1(n735), .A2(n734), .ZN(n740) );
  AND2_X1 U835 ( .A1(n928), .A2(n740), .ZN(n736) );
  NOR2_X1 U836 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U837 ( .A1(n739), .A2(n738), .ZN(n742) );
  OR2_X1 U838 ( .A1(n928), .A2(n740), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n743), .A2(n525), .ZN(n744) );
  XNOR2_X1 U840 ( .A(KEYINPUT97), .B(n744), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U842 ( .A1(G299), .A2(n747), .ZN(n748) );
  XOR2_X1 U843 ( .A(KEYINPUT28), .B(n748), .Z(n749) );
  NOR2_X1 U844 ( .A1(n750), .A2(n749), .ZN(n752) );
  XNOR2_X1 U845 ( .A(KEYINPUT98), .B(KEYINPUT29), .ZN(n751) );
  XNOR2_X1 U846 ( .A(n752), .B(n751), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G171), .A2(n753), .ZN(n760) );
  AND2_X1 U848 ( .A1(n760), .A2(n754), .ZN(n755) );
  NAND2_X1 U849 ( .A1(n761), .A2(n755), .ZN(n756) );
  NAND2_X1 U850 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n758), .A2(G8), .ZN(n759) );
  XNOR2_X1 U852 ( .A(n759), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n761), .A2(n760), .ZN(n763) );
  AND2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U855 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n785) );
  NOR2_X1 U858 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n771), .A2(n921), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n785), .A2(n772), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NAND2_X1 U862 ( .A1(n940), .A2(n932), .ZN(n773) );
  NOR2_X1 U863 ( .A1(KEYINPUT33), .A2(n773), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n778) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U866 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n791) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G8), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n789) );
  XNOR2_X1 U874 ( .A(n789), .B(n788), .ZN(n790) );
  NOR2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n806) );
  NOR2_X1 U876 ( .A1(n793), .A2(n792), .ZN(n838) );
  NAND2_X1 U877 ( .A1(G116), .A2(n891), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G128), .A2(n892), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U880 ( .A(KEYINPUT35), .B(n796), .Z(n803) );
  NAND2_X1 U881 ( .A1(n895), .A2(G140), .ZN(n797) );
  XNOR2_X1 U882 ( .A(KEYINPUT89), .B(n797), .ZN(n800) );
  NAND2_X1 U883 ( .A1(n896), .A2(G104), .ZN(n798) );
  XOR2_X1 U884 ( .A(KEYINPUT88), .B(n798), .Z(n799) );
  NOR2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U886 ( .A(KEYINPUT34), .B(n801), .Z(n802) );
  NOR2_X1 U887 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U888 ( .A(KEYINPUT36), .B(n804), .ZN(n888) );
  XNOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U890 ( .A1(n888), .A2(n826), .ZN(n979) );
  NAND2_X1 U891 ( .A1(n838), .A2(n979), .ZN(n835) );
  INV_X1 U892 ( .A(n835), .ZN(n805) );
  NOR2_X1 U893 ( .A1(n806), .A2(n805), .ZN(n825) );
  NAND2_X1 U894 ( .A1(G141), .A2(n895), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G129), .A2(n892), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n896), .A2(G105), .ZN(n809) );
  XOR2_X1 U898 ( .A(KEYINPUT38), .B(n809), .Z(n810) );
  NOR2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n891), .A2(G117), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n904) );
  NAND2_X1 U902 ( .A1(G1996), .A2(n904), .ZN(n814) );
  XOR2_X1 U903 ( .A(KEYINPUT90), .B(n814), .Z(n822) );
  NAND2_X1 U904 ( .A1(G131), .A2(n895), .ZN(n816) );
  NAND2_X1 U905 ( .A1(G95), .A2(n896), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n820) );
  NAND2_X1 U907 ( .A1(G107), .A2(n891), .ZN(n818) );
  NAND2_X1 U908 ( .A1(G119), .A2(n892), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n887) );
  INV_X1 U911 ( .A(G1991), .ZN(n828) );
  NOR2_X1 U912 ( .A1(n887), .A2(n828), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n974) );
  XOR2_X1 U914 ( .A(G1986), .B(G290), .Z(n927) );
  NAND2_X1 U915 ( .A1(n974), .A2(n927), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n838), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n841) );
  NAND2_X1 U918 ( .A1(n888), .A2(n826), .ZN(n983) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n904), .ZN(n827) );
  XOR2_X1 U920 ( .A(KEYINPUT103), .B(n827), .Z(n971) );
  INV_X1 U921 ( .A(n974), .ZN(n831) );
  NOR2_X1 U922 ( .A1(G1986), .A2(G290), .ZN(n829) );
  AND2_X1 U923 ( .A1(n828), .A2(n887), .ZN(n976) );
  NOR2_X1 U924 ( .A1(n829), .A2(n976), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U926 ( .A1(n971), .A2(n832), .ZN(n833) );
  XNOR2_X1 U927 ( .A(KEYINPUT104), .B(n833), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n834), .B(KEYINPUT39), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n983), .A2(n837), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U933 ( .A(n842), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U936 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U938 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(G69), .ZN(G235) );
  NOR2_X1 U943 ( .A1(n848), .A2(n847), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  INV_X1 U945 ( .A(n849), .ZN(G319) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n851) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1956), .B(G1961), .Z(n859) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1966), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U958 ( .A(n860), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U959 ( .A(G1976), .B(G1971), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U961 ( .A(G2474), .B(G1981), .Z(n864) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U965 ( .A1(n892), .A2(G124), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G136), .A2(n895), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U969 ( .A(KEYINPUT106), .B(n870), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G112), .A2(n891), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G100), .A2(n896), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(G162) );
  XOR2_X1 U974 ( .A(KEYINPUT107), .B(KEYINPUT46), .Z(n876) );
  XNOR2_X1 U975 ( .A(G160), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n886) );
  NAND2_X1 U977 ( .A1(G139), .A2(n895), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G103), .A2(n896), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G115), .A2(n891), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G127), .A2(n892), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n987) );
  XNOR2_X1 U985 ( .A(G164), .B(n987), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n884), .B(G162), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n906) );
  NAND2_X1 U990 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G130), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U993 ( .A1(G142), .A2(n895), .ZN(n898) );
  NAND2_X1 U994 ( .A1(G106), .A2(n896), .ZN(n897) );
  NAND2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U996 ( .A(n899), .B(KEYINPUT45), .Z(n900) );
  NOR2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(n977), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(n920), .B(G286), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(G171), .B(n908), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1005 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n914) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n915), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(KEYINPUT108), .B(n917), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1016 ( .A(KEYINPUT56), .B(G16), .ZN(n946) );
  XNOR2_X1 U1017 ( .A(n920), .B(G1341), .ZN(n938) );
  XOR2_X1 U1018 ( .A(n921), .B(KEYINPUT118), .Z(n923) );
  XNOR2_X1 U1019 ( .A(G1961), .B(G171), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n935) );
  XNOR2_X1 U1021 ( .A(G303), .B(G1971), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G299), .B(G1956), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n931) );
  XOR2_X1 U1025 ( .A(G1348), .B(n928), .Z(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT117), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(KEYINPUT119), .B(n936), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(KEYINPUT120), .B(n939), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G168), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(KEYINPUT57), .B(n942), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n1001) );
  XNOR2_X1 U1038 ( .A(KEYINPUT114), .B(KEYINPUT55), .ZN(n966) );
  XNOR2_X1 U1039 ( .A(G1991), .B(G25), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n954) );
  XOR2_X1 U1042 ( .A(G2067), .B(G26), .Z(n949) );
  NAND2_X1 U1043 ( .A1(n949), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(KEYINPUT112), .B(G1996), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G32), .B(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1048 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n959), .B(KEYINPUT113), .ZN(n964) );
  XNOR2_X1 U1052 ( .A(G2084), .B(G34), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT54), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(n966), .B(n965), .ZN(n968) );
  XOR2_X1 U1058 ( .A(G29), .B(KEYINPUT115), .Z(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n969), .B(KEYINPUT116), .ZN(n999) );
  INV_X1 U1061 ( .A(G29), .ZN(n997) );
  XOR2_X1 U1062 ( .A(G2090), .B(G162), .Z(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1064 ( .A(KEYINPUT51), .B(n972), .Z(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n985) );
  XOR2_X1 U1066 ( .A(G160), .B(G2084), .Z(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n980) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1070 ( .A(KEYINPUT109), .B(n981), .Z(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(KEYINPUT110), .B(n986), .ZN(n992) );
  XOR2_X1 U1074 ( .A(G2072), .B(n987), .Z(n989) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(KEYINPUT50), .B(n990), .ZN(n991) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1079 ( .A(n993), .B(KEYINPUT52), .Z(n994) );
  XNOR2_X1 U1080 ( .A(KEYINPUT111), .B(n994), .ZN(n995) );
  NOR2_X1 U1081 ( .A1(KEYINPUT55), .A2(n995), .ZN(n996) );
  NOR2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1083 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1084 ( .A1(n1001), .A2(n1000), .ZN(n1033) );
  XNOR2_X1 U1085 ( .A(G16), .B(KEYINPUT121), .ZN(n1030) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n1028) );
  XOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .Z(n1002) );
  XNOR2_X1 U1088 ( .A(G4), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(G6), .B(G1981), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1009), .B(KEYINPUT123), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(n1011), .B(n1010), .ZN(n1026) );
  XOR2_X1 U1098 ( .A(G1976), .B(G23), .Z(n1014) );
  XOR2_X1 U1099 ( .A(G24), .B(KEYINPUT126), .Z(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(G1986), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT125), .B(G1971), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(G22), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1018), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1019), .B(G5), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT124), .B(G1966), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(G21), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1028), .B(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(G11), .ZN(n1032) );
  NOR2_X1 U1115 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1116 ( .A(n1034), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

