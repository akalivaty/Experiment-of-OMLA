

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n332), .B(n331), .ZN(n556) );
  XNOR2_X2 U324 ( .A(n292), .B(n303), .ZN(n384) );
  XOR2_X2 U325 ( .A(G78GAT), .B(G148GAT), .Z(n292) );
  XOR2_X1 U326 ( .A(n387), .B(KEYINPUT70), .Z(n291) );
  XOR2_X1 U327 ( .A(KEYINPUT41), .B(n449), .Z(n542) );
  INV_X1 U328 ( .A(G204GAT), .ZN(n450) );
  NOR2_X1 U329 ( .A1(n536), .A2(n552), .ZN(n582) );
  XNOR2_X1 U330 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(G1353GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n334) );
  XOR2_X1 U333 ( .A(KEYINPUT91), .B(G204GAT), .Z(n294) );
  XOR2_X1 U334 ( .A(G50GAT), .B(G162GAT), .Z(n402) );
  XOR2_X1 U335 ( .A(G22GAT), .B(G155GAT), .Z(n345) );
  XNOR2_X1 U336 ( .A(n402), .B(n345), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n307) );
  XOR2_X1 U338 ( .A(KEYINPUT22), .B(G211GAT), .Z(n296) );
  XNOR2_X1 U339 ( .A(KEYINPUT23), .B(KEYINPUT86), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n298) );
  XNOR2_X1 U342 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U345 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n302) );
  XNOR2_X1 U346 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n435) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n435), .B(n384), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U351 ( .A(n307), .B(n306), .Z(n309) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n308) );
  XOR2_X1 U353 ( .A(n309), .B(n308), .Z(n313) );
  XOR2_X1 U354 ( .A(KEYINPUT21), .B(G218GAT), .Z(n311) );
  XNOR2_X1 U355 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U357 ( .A(G197GAT), .B(n312), .Z(n335) );
  XNOR2_X1 U358 ( .A(n313), .B(n335), .ZN(n553) );
  XOR2_X1 U359 ( .A(KEYINPUT83), .B(G71GAT), .Z(n315) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U362 ( .A(n316), .B(G134GAT), .Z(n318) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G127GAT), .Z(n346) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(n346), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n324) );
  XOR2_X1 U366 ( .A(G120GAT), .B(KEYINPUT81), .Z(n320) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n439) );
  XOR2_X1 U369 ( .A(G176GAT), .B(n439), .Z(n322) );
  NAND2_X1 U370 ( .A1(G227GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U372 ( .A(n324), .B(n323), .Z(n332) );
  XOR2_X1 U373 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n326) );
  XNOR2_X1 U374 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U376 ( .A(G169GAT), .B(n327), .Z(n342) );
  XOR2_X1 U377 ( .A(G183GAT), .B(KEYINPUT82), .Z(n329) );
  XNOR2_X1 U378 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n342), .B(n330), .ZN(n331) );
  NAND2_X1 U381 ( .A1(n553), .A2(n556), .ZN(n333) );
  XNOR2_X1 U382 ( .A(n334), .B(n333), .ZN(n536) );
  XOR2_X1 U383 ( .A(G36GAT), .B(G190GAT), .Z(n400) );
  XOR2_X1 U384 ( .A(n400), .B(n335), .Z(n337) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U387 ( .A(G8GAT), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n338), .B(G211GAT), .ZN(n361) );
  XOR2_X1 U389 ( .A(n339), .B(n361), .Z(n344) );
  XOR2_X1 U390 ( .A(G64GAT), .B(G92GAT), .Z(n341) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(G204GAT), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n394) );
  XNOR2_X1 U393 ( .A(n342), .B(n394), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n514) );
  XOR2_X1 U395 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n418) );
  XOR2_X1 U396 ( .A(G64GAT), .B(n345), .Z(n348) );
  XNOR2_X1 U397 ( .A(n346), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U399 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n350) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U402 ( .A(n352), .B(n351), .Z(n354) );
  XOR2_X1 U403 ( .A(G1GAT), .B(KEYINPUT67), .Z(n375) );
  XNOR2_X1 U404 ( .A(n375), .B(KEYINPUT76), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U406 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n356) );
  XNOR2_X1 U407 ( .A(KEYINPUT14), .B(KEYINPUT77), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U409 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U410 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n360) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G57GAT), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n393) );
  XNOR2_X1 U413 ( .A(n361), .B(n393), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n578) );
  XNOR2_X1 U415 ( .A(KEYINPUT112), .B(n578), .ZN(n564) );
  XOR2_X1 U416 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n365) );
  XNOR2_X1 U417 ( .A(G8GAT), .B(KEYINPUT64), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n379) );
  XOR2_X1 U419 ( .A(G197GAT), .B(G22GAT), .Z(n367) );
  XNOR2_X1 U420 ( .A(G50GAT), .B(G36GAT), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U422 ( .A(G15GAT), .B(G113GAT), .Z(n369) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(G141GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U426 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n373) );
  NAND2_X1 U427 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U432 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n381) );
  XNOR2_X1 U433 ( .A(G43GAT), .B(G29GAT), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U435 ( .A(KEYINPUT7), .B(n382), .ZN(n399) );
  XOR2_X1 U436 ( .A(n383), .B(n399), .Z(n539) );
  XOR2_X1 U437 ( .A(n384), .B(KEYINPUT73), .Z(n386) );
  NAND2_X1 U438 ( .A1(G230GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U440 ( .A(G99GAT), .B(G85GAT), .Z(n401) );
  XNOR2_X1 U441 ( .A(G120GAT), .B(n401), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n291), .B(n388), .ZN(n392) );
  XOR2_X1 U443 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n390) );
  XNOR2_X1 U444 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U446 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n396), .B(n395), .ZN(n449) );
  NOR2_X1 U449 ( .A1(n539), .A2(n542), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n397), .B(KEYINPUT46), .ZN(n398) );
  NOR2_X1 U451 ( .A1(n564), .A2(n398), .ZN(n416) );
  INV_X1 U452 ( .A(n399), .ZN(n415) );
  XOR2_X1 U453 ( .A(n401), .B(n400), .Z(n404) );
  XOR2_X1 U454 ( .A(G134GAT), .B(KEYINPUT75), .Z(n438) );
  XNOR2_X1 U455 ( .A(n402), .B(n438), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U457 ( .A(KEYINPUT74), .B(G92GAT), .Z(n406) );
  NAND2_X1 U458 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U460 ( .A(n408), .B(n407), .Z(n413) );
  XOR2_X1 U461 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n410) );
  XNOR2_X1 U462 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U464 ( .A(G106GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U465 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U466 ( .A(n415), .B(n414), .Z(n569) );
  INV_X1 U467 ( .A(n569), .ZN(n550) );
  NAND2_X1 U468 ( .A1(n416), .A2(n550), .ZN(n417) );
  XNOR2_X1 U469 ( .A(n418), .B(n417), .ZN(n424) );
  INV_X1 U470 ( .A(n539), .ZN(n575) );
  XNOR2_X1 U471 ( .A(KEYINPUT36), .B(n550), .ZN(n584) );
  INV_X1 U472 ( .A(n578), .ZN(n546) );
  NOR2_X1 U473 ( .A1(n584), .A2(n546), .ZN(n419) );
  XOR2_X1 U474 ( .A(KEYINPUT45), .B(n419), .Z(n420) );
  NOR2_X1 U475 ( .A1(n575), .A2(n420), .ZN(n421) );
  NAND2_X1 U476 ( .A1(n449), .A2(n421), .ZN(n422) );
  XOR2_X1 U477 ( .A(KEYINPUT114), .B(n422), .Z(n423) );
  NOR2_X1 U478 ( .A1(n424), .A2(n423), .ZN(n425) );
  XNOR2_X1 U479 ( .A(KEYINPUT48), .B(n425), .ZN(n523) );
  NOR2_X1 U480 ( .A1(n514), .A2(n523), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n426), .B(KEYINPUT54), .ZN(n448) );
  XOR2_X1 U482 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n447) );
  XOR2_X1 U485 ( .A(G85GAT), .B(G155GAT), .Z(n430) );
  XNOR2_X1 U486 ( .A(G127GAT), .B(G148GAT), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n432) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(G57GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U491 ( .A(n434), .B(n433), .Z(n445) );
  XOR2_X1 U492 ( .A(n435), .B(KEYINPUT94), .Z(n437) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U495 ( .A(n438), .B(G162GAT), .Z(n441) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n511) );
  NAND2_X1 U501 ( .A1(n448), .A2(n511), .ZN(n552) );
  INV_X1 U502 ( .A(n449), .ZN(n454) );
  NAND2_X1 U503 ( .A1(n582), .A2(n454), .ZN(n453) );
  XOR2_X1 U504 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n451) );
  NOR2_X1 U505 ( .A1(n454), .A2(n539), .ZN(n485) );
  XNOR2_X1 U506 ( .A(n514), .B(KEYINPUT27), .ZN(n462) );
  NOR2_X1 U507 ( .A1(n536), .A2(n462), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT98), .B(n455), .Z(n459) );
  NOR2_X1 U509 ( .A1(n556), .A2(n514), .ZN(n456) );
  NOR2_X1 U510 ( .A1(n553), .A2(n456), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT25), .B(n457), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U513 ( .A1(n511), .A2(n460), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n461), .B(KEYINPUT99), .ZN(n465) );
  XNOR2_X1 U515 ( .A(n553), .B(KEYINPUT28), .ZN(n476) );
  NOR2_X1 U516 ( .A1(n511), .A2(n462), .ZN(n521) );
  NAND2_X1 U517 ( .A1(n556), .A2(n521), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n476), .A2(n463), .ZN(n464) );
  NOR2_X1 U519 ( .A1(n465), .A2(n464), .ZN(n480) );
  NAND2_X1 U520 ( .A1(n550), .A2(n578), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT80), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT16), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n480), .A2(n468), .ZN(n499) );
  NAND2_X1 U524 ( .A1(n485), .A2(n499), .ZN(n477) );
  NOR2_X1 U525 ( .A1(n511), .A2(n477), .ZN(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U528 ( .A(G1GAT), .B(n471), .Z(G1324GAT) );
  NOR2_X1 U529 ( .A1(n514), .A2(n477), .ZN(n472) );
  XOR2_X1 U530 ( .A(G8GAT), .B(n472), .Z(G1325GAT) );
  NOR2_X1 U531 ( .A1(n556), .A2(n477), .ZN(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U534 ( .A(G15GAT), .B(n475), .Z(G1326GAT) );
  INV_X1 U535 ( .A(n476), .ZN(n524) );
  NOR2_X1 U536 ( .A1(n524), .A2(n477), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT102), .B(n478), .Z(n479) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(n479), .ZN(G1327GAT) );
  INV_X1 U539 ( .A(KEYINPUT104), .ZN(n488) );
  INV_X1 U540 ( .A(KEYINPUT37), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n584), .A2(n480), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n546), .A2(n481), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT103), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n510) );
  AND2_X1 U545 ( .A1(n510), .A2(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT38), .B(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n496) );
  NOR2_X1 U548 ( .A1(n511), .A2(n496), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n514), .A2(n496), .ZN(n491) );
  XOR2_X1 U552 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n493) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n495) );
  NOR2_X1 U556 ( .A1(n556), .A2(n496), .ZN(n494) );
  XOR2_X1 U557 ( .A(n495), .B(n494), .Z(G1330GAT) );
  NOR2_X1 U558 ( .A1(n524), .A2(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  NOR2_X1 U561 ( .A1(n575), .A2(n542), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n509), .A2(n499), .ZN(n504) );
  NOR2_X1 U563 ( .A1(n511), .A2(n504), .ZN(n500) );
  XOR2_X1 U564 ( .A(n500), .B(KEYINPUT42), .Z(n501) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n504), .ZN(n502) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n556), .A2(n504), .ZN(n503) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n503), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n504), .A2(n524), .ZN(n508) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n506) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT108), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n517) );
  NOR2_X1 U576 ( .A1(n511), .A2(n517), .ZN(n512) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n512), .Z(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT110), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n517), .ZN(n515) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n556), .A2(n517), .ZN(n516) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n524), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  XOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT115), .Z(n527) );
  INV_X1 U588 ( .A(n521), .ZN(n522) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n524), .A2(n538), .ZN(n525) );
  NOR2_X1 U591 ( .A1(n556), .A2(n525), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n532), .A2(n575), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n529) );
  INV_X1 U595 ( .A(n542), .ZN(n561) );
  NAND2_X1 U596 ( .A1(n532), .A2(n561), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  NAND2_X1 U598 ( .A1(n564), .A2(n532), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U602 ( .A1(n532), .A2(n569), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n535), .ZN(G1343GAT) );
  INV_X1 U605 ( .A(n536), .ZN(n537) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n539), .A2(n549), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n542), .A2(n549), .ZN(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n549), .ZN(n547) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(n547), .Z(n548) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT55), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n570) );
  NAND2_X1 U622 ( .A1(n570), .A2(n575), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n559) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(n560), .Z(n563) );
  NAND2_X1 U628 ( .A1(n570), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  XOR2_X1 U630 ( .A(G183GAT), .B(KEYINPUT121), .Z(n566) );
  NAND2_X1 U631 ( .A1(n570), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT123), .B(n568), .Z(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1351GAT) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT59), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(n574), .Z(n577) );
  NAND2_X1 U641 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NAND2_X1 U643 ( .A1(n582), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n586) );
  INV_X1 U648 ( .A(n582), .ZN(n583) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

