//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT94), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G8gat), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  AOI21_X1  g013(.A(G1gat), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n210), .A2(new_n215), .A3(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT92), .ZN(new_n226));
  NOR3_X1   g025(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT92), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G29gat), .A2(G36gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n221), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n221), .A2(new_n232), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n230), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT93), .B(KEYINPUT15), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n220), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT96), .B1(new_n219), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n210), .A2(new_n215), .A3(new_n212), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n215), .B1(new_n210), .B2(new_n212), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n230), .B1(new_n227), .B2(new_n228), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n225), .A2(KEYINPUT92), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n232), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n221), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n220), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT93), .B(KEYINPUT15), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(new_n221), .A3(new_n232), .A4(new_n235), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n243), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n240), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n243), .A2(KEYINPUT96), .A3(new_n253), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT95), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT13), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(KEYINPUT17), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT17), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n248), .A2(new_n252), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n243), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n219), .A2(new_n239), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n264), .A2(new_n265), .A3(new_n258), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n260), .B1(new_n266), .B2(KEYINPUT18), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT18), .ZN(new_n268));
  NOR4_X1   g067(.A1(new_n264), .A2(new_n265), .A3(new_n268), .A4(new_n258), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n206), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n264), .ZN(new_n271));
  INV_X1    g070(.A(new_n258), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n254), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  INV_X1    g073(.A(new_n269), .ZN(new_n275));
  INV_X1    g074(.A(new_n206), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(new_n260), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT87), .ZN(new_n279));
  XOR2_X1   g078(.A(G141gat), .B(G148gat), .Z(new_n280));
  INV_X1    g079(.A(G155gat), .ZN(new_n281));
  INV_X1    g080(.A(G162gat), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT2), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G155gat), .B(G162gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n285), .A3(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291));
  INV_X1    g090(.A(G211gat), .ZN(new_n292));
  INV_X1    g091(.A(G218gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n297));
  INV_X1    g096(.A(G204gat), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n300));
  AOI21_X1  g099(.A(G204gat), .B1(new_n300), .B2(new_n295), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n294), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G211gat), .B(G218gat), .Z(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n298), .B1(new_n296), .B2(new_n297), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(G204gat), .A3(new_n295), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n294), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n289), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n290), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT85), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n287), .A2(new_n317), .A3(new_n288), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n312), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT74), .B1(new_n304), .B2(new_n309), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT85), .B(new_n290), .C1(new_n311), .C2(new_n313), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n316), .A2(new_n323), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT86), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n310), .B(new_n320), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n324), .B1(new_n329), .B2(new_n319), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n316), .A4(new_n326), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n287), .A2(KEYINPUT77), .A3(new_n288), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT77), .B1(new_n287), .B2(new_n288), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n304), .A2(KEYINPUT82), .A3(new_n309), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n308), .B1(new_n307), .B2(new_n294), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g140(.A(KEYINPUT83), .B(new_n336), .C1(new_n341), .C2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT3), .B1(new_n337), .B2(new_n340), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n334), .A2(new_n335), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n346), .A3(new_n323), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n324), .B(KEYINPUT81), .Z(new_n349));
  AND3_X1   g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n347), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n333), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G22gat), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n333), .B(new_n354), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n353), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n353), .B2(new_n355), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n279), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n349), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT84), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n354), .B1(new_n366), .B2(new_n333), .ZN(new_n367));
  INV_X1    g166(.A(new_n355), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n355), .A3(new_n358), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(KEYINPUT87), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT68), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  INV_X1    g173(.A(G120gat), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT1), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G113gat), .A2(G120gat), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n372), .A2(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n373), .B2(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(new_n372), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(KEYINPUT68), .A3(new_n377), .A4(new_n376), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n290), .A3(new_n318), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n287), .A3(new_n288), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n382), .C1(new_n334), .C2(new_n335), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n390), .A3(KEYINPUT79), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(new_n393), .A3(KEYINPUT4), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n386), .A2(new_n391), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n289), .A2(new_n381), .A3(new_n379), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n385), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT78), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n400));
  AOI211_X1 g199(.A(new_n400), .B(new_n385), .C1(new_n387), .C2(new_n396), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n389), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT4), .B(new_n382), .C1(new_n334), .C2(new_n335), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n385), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT5), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n395), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G1gat), .B(G29gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n408), .B2(new_n413), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n413), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n419), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  AND2_X1   g224(.A1(G226gat), .A2(G233gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(KEYINPUT29), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n429), .A2(KEYINPUT23), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(KEYINPUT23), .ZN(new_n431));
  INV_X1    g230(.A(G169gat), .ZN(new_n432));
  INV_X1    g231(.A(G176gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT24), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(G183gat), .A3(G190gat), .ZN(new_n439));
  INV_X1    g238(.A(G183gat), .ZN(new_n440));
  INV_X1    g239(.A(G190gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(new_n442), .B2(new_n438), .ZN(new_n443));
  XOR2_X1   g242(.A(KEYINPUT65), .B(G183gat), .Z(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(G190gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n445), .A3(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n441), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT64), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n436), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n449), .B2(KEYINPUT25), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n434), .A2(KEYINPUT26), .A3(new_n429), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n442), .B(new_n451), .C1(KEYINPUT26), .C2(new_n429), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT27), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G183gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n440), .A2(KEYINPUT27), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT28), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(G190gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n453), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n460));
  AOI21_X1  g259(.A(G190gat), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n459), .B(new_n461), .C1(new_n444), .C2(new_n453), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n458), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n452), .B1(new_n463), .B2(KEYINPUT67), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n450), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT75), .B(new_n450), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n428), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n464), .A2(new_n465), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n426), .A3(new_n450), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n470), .A2(new_n473), .A3(new_n329), .ZN(new_n474));
  INV_X1    g273(.A(new_n329), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n468), .A2(new_n426), .A3(new_n469), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n466), .A2(new_n427), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n425), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT30), .B(new_n425), .C1(new_n474), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n468), .A2(new_n469), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n427), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n475), .A3(new_n472), .ZN(new_n485));
  INV_X1    g284(.A(new_n425), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n476), .A2(new_n477), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n475), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n481), .A2(KEYINPUT76), .A3(new_n482), .A4(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n482), .A2(KEYINPUT76), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n361), .A2(new_n371), .B1(new_n422), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT69), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(new_n450), .C1(new_n464), .C2(new_n465), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n382), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G227gat), .ZN(new_n497));
  INV_X1    g296(.A(G233gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n471), .A2(new_n494), .A3(new_n383), .A4(new_n450), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT32), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G15gat), .B(G43gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G71gat), .B(G99gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n502), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT33), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n501), .A2(KEYINPUT32), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n497), .B2(new_n498), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT34), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT34), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n516), .B(new_n519), .C1(new_n497), .C2(new_n498), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n510), .A2(new_n518), .A3(new_n520), .A4(new_n514), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT36), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT36), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT88), .B1(new_n492), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n422), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n359), .A2(new_n360), .A3(new_n279), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT87), .B1(new_n369), .B2(new_n370), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533));
  INV_X1    g332(.A(new_n526), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n524), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n391), .A2(new_n384), .A3(new_n394), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n398), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n538), .B(KEYINPUT39), .C1(new_n398), .C2(new_n397), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n412), .B(KEYINPUT90), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(new_n541), .C1(KEYINPUT39), .C2(new_n538), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT40), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n408), .A2(new_n544), .A3(new_n540), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n408), .B2(new_n540), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n542), .A2(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n543), .B2(new_n542), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n489), .A2(new_n549), .A3(new_n490), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n489), .B2(new_n490), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n359), .A2(new_n360), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n417), .B1(new_n545), .B2(new_n546), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n414), .A3(new_n479), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n425), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n488), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n476), .A2(new_n477), .A3(new_n475), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT37), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n475), .B1(new_n484), .B2(new_n472), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT38), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n556), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n485), .B1(new_n487), .B2(new_n475), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n560), .B1(new_n557), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT38), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n554), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n528), .A2(new_n536), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n522), .A2(new_n523), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n554), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n552), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT35), .B1(new_n555), .B2(new_n414), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n550), .A4(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n369), .A2(new_n370), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT35), .B1(new_n580), .B2(new_n529), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n278), .B1(new_n572), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(G57gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(KEYINPUT97), .ZN(new_n586));
  AND2_X1   g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(G57gat), .A3(G64gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n587), .B2(KEYINPUT9), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT98), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n585), .A2(KEYINPUT97), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(G64gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  XNOR2_X1  g396(.A(G71gat), .B(G78gat), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n586), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(G57gat), .B2(G64gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n598), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(G127gat), .Z(new_n610));
  OAI21_X1  g409(.A(new_n219), .B1(new_n606), .B2(new_n605), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n281), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  OR2_X1    g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n261), .A2(new_n263), .ZN(new_n620));
  NAND2_X1  g419(.A1(G85gat), .A2(G92gat), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT8), .ZN(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n624), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G99gat), .ZN(new_n631));
  INV_X1    g430(.A(G106gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n625), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT100), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n636), .A3(new_n625), .ZN(new_n637));
  NOR2_X1   g436(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n621), .ZN(new_n639));
  NAND2_X1  g438(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n630), .A2(new_n635), .A3(new_n637), .A4(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n626), .A3(new_n629), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n644), .A2(new_n638), .A3(new_n621), .ZN(new_n645));
  OAI211_X1 g444(.A(KEYINPUT100), .B(new_n634), .C1(new_n643), .C2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n620), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n642), .A2(new_n646), .ZN(new_n649));
  AND2_X1   g448(.A1(G232gat), .A2(G233gat), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n253), .A2(new_n649), .B1(KEYINPUT41), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G190gat), .B(G218gat), .Z(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n650), .A2(KEYINPUT41), .ZN(new_n656));
  XNOR2_X1  g455(.A(G134gat), .B(G162gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n654), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n654), .B2(new_n655), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n619), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n603), .B1(new_n593), .B2(new_n599), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n649), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n665), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT102), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n647), .A2(new_n605), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n649), .A2(new_n665), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n671), .A2(KEYINPUT102), .A3(new_n672), .A4(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n666), .A2(KEYINPUT10), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(KEYINPUT103), .B(new_n664), .C1(new_n670), .C2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(new_n672), .A3(new_n669), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n674), .A3(new_n673), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT103), .B1(new_n681), .B2(new_n664), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n664), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n666), .B2(new_n667), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(G120gat), .B(G148gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT104), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  NOR2_X1   g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n681), .A2(new_n664), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n690), .B1(new_n694), .B2(new_n686), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n663), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n583), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n422), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(G1gat), .Z(G1324gat));
  NAND2_X1  g499(.A1(new_n572), .A2(new_n582), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n270), .A2(new_n277), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n575), .A2(new_n550), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT16), .B(G8gat), .Z(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n697), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n708), .A2(KEYINPUT105), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n211), .B1(new_n706), .B2(new_n697), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n708), .B1(new_n714), .B2(new_n709), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n710), .B1(new_n713), .B2(new_n715), .ZN(G1325gat));
  OAI21_X1  g515(.A(G15gat), .B1(new_n698), .B2(new_n535), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n573), .A2(G15gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n698), .B2(new_n718), .ZN(G1326gat));
  NOR2_X1   g518(.A1(new_n530), .A2(new_n531), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n583), .A2(new_n721), .A3(new_n697), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  INV_X1    g523(.A(new_n422), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n619), .A2(new_n696), .ZN(new_n726));
  INV_X1    g525(.A(new_n662), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n583), .A2(new_n223), .A3(new_n725), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT45), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n662), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n701), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n492), .A2(new_n527), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n571), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n582), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT44), .B1(new_n737), .B2(new_n727), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n726), .A2(new_n702), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT106), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n734), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n725), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n731), .B1(new_n743), .B2(new_n223), .ZN(G1328gat));
  NOR4_X1   g543(.A1(new_n703), .A2(G36gat), .A3(new_n705), .A4(new_n728), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT46), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n742), .A2(new_n704), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n224), .B2(new_n747), .ZN(G1329gat));
  XNOR2_X1  g547(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n734), .A2(new_n738), .A3(new_n535), .A4(new_n741), .ZN(new_n751));
  INV_X1    g550(.A(G43gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n729), .A2(new_n752), .A3(new_n578), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n703), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI221_X1 g555(.A(new_n749), .B1(new_n703), .B2(new_n754), .C1(new_n751), .C2(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1330gat));
  NOR2_X1   g557(.A1(new_n728), .A2(G50gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n583), .A2(new_n721), .A3(new_n759), .ZN(new_n760));
  NOR4_X1   g559(.A1(new_n734), .A2(new_n738), .A3(new_n579), .A4(new_n741), .ZN(new_n761));
  INV_X1    g560(.A(G50gat), .ZN(new_n762));
  OAI211_X1 g561(.A(KEYINPUT48), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n701), .A2(new_n733), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n571), .A2(new_n735), .B1(new_n577), .B2(new_n581), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n732), .B1(new_n765), .B2(new_n662), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n764), .A2(new_n766), .A3(new_n721), .A4(new_n740), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n767), .A2(new_n768), .A3(G50gat), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(G50gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n583), .A2(new_n772), .A3(new_n721), .A4(new_n759), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n769), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n763), .B1(new_n775), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g575(.A(new_n696), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n663), .A2(new_n702), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n737), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n422), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(new_n585), .ZN(G1332gat));
  NOR2_X1   g580(.A1(new_n779), .A2(new_n705), .ZN(new_n782));
  NOR2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  AND2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n782), .B2(new_n783), .ZN(G1333gat));
  OR3_X1    g585(.A1(new_n779), .A2(KEYINPUT111), .A3(new_n573), .ZN(new_n787));
  INV_X1    g586(.A(G71gat), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT111), .B1(new_n779), .B2(new_n573), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n737), .A2(G71gat), .A3(new_n527), .A4(new_n778), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT110), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n790), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1334gat));
  NOR2_X1   g596(.A1(new_n779), .A2(new_n720), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g598(.A1(new_n619), .A2(new_n702), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n696), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n734), .A2(new_n738), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n422), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n737), .A2(new_n727), .A3(new_n800), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n809), .A2(new_n627), .A3(new_n725), .A4(new_n696), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n810), .ZN(G1336gat));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR4_X1   g612(.A1(new_n734), .A2(new_n738), .A3(new_n705), .A4(new_n801), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n628), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n704), .A2(new_n628), .A3(new_n696), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT112), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n807), .B2(new_n808), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n813), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n809), .A2(new_n817), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n812), .C1(new_n628), .C2(new_n814), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n803), .B2(new_n535), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n631), .A3(new_n578), .A4(new_n696), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1338gat));
  NAND2_X1  g625(.A1(new_n802), .A2(new_n721), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n579), .A2(G106gat), .A3(new_n777), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n827), .A2(G106gat), .B1(new_n809), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n632), .B1(new_n802), .B2(new_n554), .ZN(new_n831));
  INV_X1    g630(.A(new_n808), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n805), .A2(new_n806), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n828), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n830), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(new_n835), .ZN(G1339gat));
  INV_X1    g635(.A(new_n619), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n681), .B2(new_n664), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n677), .A2(new_n839), .A3(new_n682), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n690), .B1(new_n693), .B2(KEYINPUT54), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT103), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n693), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n670), .A2(new_n675), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n684), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n847), .A3(new_n676), .ZN(new_n848));
  INV_X1    g647(.A(new_n841), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT55), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n842), .A2(new_n702), .A3(new_n692), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n272), .B1(new_n271), .B2(new_n254), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n259), .B1(new_n255), .B2(new_n256), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n205), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n277), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n696), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n727), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n727), .A3(new_n856), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n850), .A2(new_n692), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n837), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n619), .A2(new_n278), .A3(new_n662), .A4(new_n777), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n422), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n704), .A2(new_n580), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n702), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n864), .A2(new_n721), .ZN(new_n870));
  AND4_X1   g669(.A1(new_n725), .A2(new_n870), .A3(new_n578), .A4(new_n705), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n278), .A2(new_n374), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n868), .B2(new_n696), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n777), .A2(new_n375), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n871), .B2(new_n875), .ZN(G1341gat));
  NOR3_X1   g675(.A1(new_n867), .A2(G127gat), .A3(new_n837), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n871), .A2(new_n619), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(G127gat), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT114), .Z(G1342gat));
  OR3_X1    g679(.A1(new_n867), .A2(G134gat), .A3(new_n662), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n871), .A2(new_n727), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G134gat), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  INV_X1    g687(.A(new_n863), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n855), .B1(new_n692), .B2(new_n695), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n841), .B1(new_n683), .B2(new_n847), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n891), .A2(KEYINPUT55), .B1(new_n683), .B2(new_n691), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n848), .A2(new_n849), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n278), .B1(new_n893), .B2(new_n838), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT115), .B1(new_n895), .B2(new_n727), .ZN(new_n896));
  INV_X1    g695(.A(new_n861), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n702), .B1(new_n891), .B2(KEYINPUT55), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n857), .B1(new_n898), .B2(new_n860), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n662), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n889), .B1(new_n902), .B2(new_n837), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n720), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT116), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n899), .A2(new_n662), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n861), .B1(new_n909), .B2(KEYINPUT115), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n619), .B1(new_n910), .B2(new_n901), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n908), .B(new_n905), .C1(new_n911), .C2(new_n889), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n579), .B1(new_n862), .B2(new_n863), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n904), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n704), .A2(new_n527), .A3(new_n422), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n702), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G141gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n862), .A2(new_n863), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n527), .A2(new_n579), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n725), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n278), .A2(G141gat), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n922), .A2(new_n704), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n888), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n922), .A2(KEYINPUT117), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n920), .A2(new_n921), .A3(new_n929), .A4(new_n725), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n705), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n888), .B1(new_n931), .B2(new_n924), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n932), .B1(new_n918), .B2(G141gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n887), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n932), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n925), .B1(new_n918), .B2(G141gat), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n936), .B(KEYINPUT118), .C1(new_n888), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(G1344gat));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT120), .B1(new_n913), .B2(KEYINPUT57), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n904), .B1(new_n864), .B2(new_n720), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n913), .A2(KEYINPUT57), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n944), .B2(KEYINPUT120), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n917), .A2(new_n696), .ZN(new_n946));
  OAI21_X1  g745(.A(G148gat), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n916), .A2(new_n696), .A3(new_n917), .ZN(new_n950));
  INV_X1    g749(.A(G148gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(KEYINPUT59), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n947), .A2(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n931), .A2(G148gat), .A3(new_n777), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n940), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n954), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n950), .A2(new_n952), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n942), .B2(new_n943), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n696), .B(new_n917), .C1(new_n959), .C2(new_n941), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n948), .B1(new_n960), .B2(G148gat), .ZN(new_n961));
  OAI211_X1 g760(.A(KEYINPUT121), .B(new_n956), .C1(new_n957), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n955), .A2(new_n962), .ZN(G1345gat));
  AND2_X1   g762(.A1(new_n916), .A2(new_n917), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(G155gat), .A3(new_n619), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n928), .A2(new_n705), .A3(new_n930), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n619), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n966), .A3(new_n619), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n281), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n965), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n965), .B(KEYINPUT123), .C1(new_n968), .C2(new_n970), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1346gat));
  AOI21_X1  g774(.A(G162gat), .B1(new_n967), .B2(new_n727), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n662), .A2(new_n282), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n964), .B2(new_n977), .ZN(G1347gat));
  NOR3_X1   g777(.A1(new_n705), .A2(new_n725), .A3(new_n580), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n920), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(G169gat), .B1(new_n981), .B2(new_n702), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n705), .A2(new_n725), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n870), .A2(new_n578), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n278), .A2(new_n432), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1348gat));
  NAND3_X1  g785(.A1(new_n981), .A2(new_n433), .A3(new_n696), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n984), .A2(new_n696), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n988), .B2(new_n433), .ZN(G1349gat));
  NOR3_X1   g788(.A1(new_n980), .A2(new_n456), .A3(new_n837), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n984), .A2(new_n619), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n990), .B1(new_n991), .B2(new_n444), .ZN(new_n992));
  XOR2_X1   g791(.A(new_n992), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g792(.A(new_n441), .B1(new_n984), .B2(new_n727), .ZN(new_n994));
  XOR2_X1   g793(.A(new_n994), .B(KEYINPUT61), .Z(new_n995));
  NAND3_X1  g794(.A1(new_n981), .A2(new_n441), .A3(new_n727), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1351gat));
  NAND2_X1  g796(.A1(new_n983), .A2(new_n535), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n999), .B1(new_n959), .B2(new_n941), .ZN(new_n1000));
  OAI21_X1  g799(.A(G197gat), .B1(new_n1000), .B2(new_n278), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n998), .A2(new_n914), .ZN(new_n1002));
  INV_X1    g801(.A(G197gat), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1002), .A2(new_n1003), .A3(new_n702), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT124), .ZN(G1352gat));
  XNOR2_X1  g805(.A(KEYINPUT125), .B(G204gat), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n777), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1010));
  OAI21_X1  g809(.A(new_n1007), .B1(new_n1000), .B2(new_n777), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1353gat));
  OAI211_X1 g811(.A(new_n619), .B(new_n999), .C1(new_n959), .C2(new_n941), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g814(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g815(.A(G211gat), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1017));
  OAI21_X1  g816(.A(KEYINPUT63), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OR2_X1    g817(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT63), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n1019), .A2(new_n1020), .A3(G211gat), .A4(new_n1015), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1002), .A2(new_n292), .A3(new_n619), .ZN(new_n1022));
  XOR2_X1   g821(.A(new_n1022), .B(KEYINPUT126), .Z(new_n1023));
  NAND3_X1  g822(.A1(new_n1018), .A2(new_n1021), .A3(new_n1023), .ZN(G1354gat));
  OAI21_X1  g823(.A(G218gat), .B1(new_n1000), .B2(new_n662), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1002), .A2(new_n293), .A3(new_n727), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1025), .A2(new_n1026), .ZN(G1355gat));
endmodule


