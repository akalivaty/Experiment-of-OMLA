

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X2 U550 ( .A(KEYINPUT17), .B(n527), .Z(n678) );
  NOR2_X1 U551 ( .A1(n531), .A2(n530), .ZN(G160) );
  NAND2_X1 U552 ( .A1(n814), .A2(n813), .ZN(n516) );
  NOR2_X1 U553 ( .A1(n763), .A2(n754), .ZN(n517) );
  NOR2_X1 U554 ( .A1(n752), .A2(n763), .ZN(n518) );
  NOR2_X1 U555 ( .A1(n808), .A2(n807), .ZN(n519) );
  XOR2_X1 U556 ( .A(n749), .B(KEYINPUT107), .Z(n520) );
  XNOR2_X1 U557 ( .A(KEYINPUT30), .B(KEYINPUT102), .ZN(n687) );
  XNOR2_X1 U558 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U559 ( .A1(n694), .A2(n693), .ZN(n695) );
  INV_X1 U560 ( .A(KEYINPUT105), .ZN(n726) );
  NAND2_X1 U561 ( .A1(G160), .A2(n685), .ZN(n728) );
  NAND2_X1 U562 ( .A1(G8), .A2(n728), .ZN(n763) );
  NOR2_X1 U563 ( .A1(G651), .A2(n648), .ZN(n643) );
  INV_X1 U564 ( .A(G2105), .ZN(n526) );
  AND2_X1 U565 ( .A1(G2104), .A2(n526), .ZN(n521) );
  XNOR2_X2 U566 ( .A(n521), .B(KEYINPUT64), .ZN(n878) );
  NAND2_X1 U567 ( .A1(n878), .A2(G101), .ZN(n522) );
  XOR2_X1 U568 ( .A(KEYINPUT23), .B(n522), .Z(n525) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U570 ( .A1(G113), .A2(n873), .ZN(n523) );
  XOR2_X1 U571 ( .A(KEYINPUT65), .B(n523), .Z(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n526), .ZN(n875) );
  NAND2_X1 U574 ( .A1(G125), .A2(n875), .ZN(n529) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  NAND2_X1 U576 ( .A1(G137), .A2(n678), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n529), .A2(n528), .ZN(n530) );
  INV_X1 U578 ( .A(G651), .ZN(n536) );
  NOR2_X1 U579 ( .A1(G543), .A2(n536), .ZN(n532) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n532), .Z(n647) );
  NAND2_X1 U581 ( .A1(G64), .A2(n647), .ZN(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n648) );
  NAND2_X1 U583 ( .A1(G52), .A2(n643), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n541) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U586 ( .A1(n637), .A2(G90), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT67), .B(n535), .Z(n538) );
  NOR2_X1 U588 ( .A1(n648), .A2(n536), .ZN(n638) );
  NAND2_X1 U589 ( .A1(n638), .A2(G77), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U592 ( .A1(n541), .A2(n540), .ZN(G171) );
  INV_X1 U593 ( .A(G132), .ZN(G219) );
  INV_X1 U594 ( .A(G82), .ZN(G220) );
  NAND2_X1 U595 ( .A1(G94), .A2(G452), .ZN(n542) );
  XOR2_X1 U596 ( .A(KEYINPUT68), .B(n542), .Z(G173) );
  NAND2_X1 U597 ( .A1(G7), .A2(G661), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n543), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U599 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n545) );
  XNOR2_X1 U600 ( .A(G223), .B(KEYINPUT71), .ZN(n821) );
  NAND2_X1 U601 ( .A1(G567), .A2(n821), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n545), .B(n544), .ZN(G234) );
  XOR2_X1 U603 ( .A(KEYINPUT12), .B(KEYINPUT75), .Z(n547) );
  NAND2_X1 U604 ( .A1(G81), .A2(n637), .ZN(n546) );
  XNOR2_X1 U605 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U606 ( .A(KEYINPUT74), .B(n548), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n638), .A2(G68), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT13), .B(n551), .Z(n555) );
  NAND2_X1 U610 ( .A1(G56), .A2(n647), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n552), .B(KEYINPUT14), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n553), .B(KEYINPUT73), .ZN(n554) );
  NOR2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U614 ( .A(n556), .B(KEYINPUT76), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G43), .A2(n643), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n966) );
  INV_X1 U617 ( .A(G860), .ZN(n607) );
  OR2_X1 U618 ( .A1(n966), .A2(n607), .ZN(G153) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  NAND2_X1 U620 ( .A1(G868), .A2(G301), .ZN(n568) );
  NAND2_X1 U621 ( .A1(n643), .A2(G54), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G92), .A2(n637), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G79), .A2(n638), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G66), .A2(n647), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT77), .B(n561), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT15), .B(n566), .Z(n961) );
  INV_X1 U630 ( .A(G868), .ZN(n586) );
  NAND2_X1 U631 ( .A1(n961), .A2(n586), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(G284) );
  NAND2_X1 U633 ( .A1(G65), .A2(n647), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G53), .A2(n643), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G91), .A2(n637), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G78), .A2(n638), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n971) );
  XNOR2_X1 U640 ( .A(n971), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U641 ( .A1(G63), .A2(n647), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G51), .A2(n643), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(KEYINPUT6), .B(n577), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n637), .A2(G89), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n578), .B(KEYINPUT4), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G76), .A2(n638), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U649 ( .A(n581), .B(KEYINPUT5), .Z(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT7), .B(n584), .Z(n585) );
  XNOR2_X1 U652 ( .A(KEYINPUT78), .B(n585), .ZN(G168) );
  XOR2_X1 U653 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U654 ( .A1(G299), .A2(n586), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G868), .A2(G286), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U657 ( .A(KEYINPUT79), .B(n589), .Z(G297) );
  NAND2_X1 U658 ( .A1(n607), .A2(G559), .ZN(n590) );
  INV_X1 U659 ( .A(n961), .ZN(n605) );
  NAND2_X1 U660 ( .A1(n590), .A2(n605), .ZN(n591) );
  XNOR2_X1 U661 ( .A(n591), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U662 ( .A1(G868), .A2(n966), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G868), .A2(n605), .ZN(n592) );
  NOR2_X1 U664 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U666 ( .A1(G111), .A2(n873), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G99), .A2(n878), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n875), .A2(G123), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT18), .B(n597), .Z(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n678), .A2(G135), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n922) );
  XOR2_X1 U674 ( .A(G2096), .B(KEYINPUT80), .Z(n602) );
  XNOR2_X1 U675 ( .A(n922), .B(n602), .ZN(n604) );
  INV_X1 U676 ( .A(G2100), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(G156) );
  NAND2_X1 U678 ( .A1(G559), .A2(n605), .ZN(n606) );
  XOR2_X1 U679 ( .A(n966), .B(n606), .Z(n657) );
  NAND2_X1 U680 ( .A1(n607), .A2(n657), .ZN(n616) );
  NAND2_X1 U681 ( .A1(n643), .A2(G55), .ZN(n608) );
  XOR2_X1 U682 ( .A(KEYINPUT81), .B(n608), .Z(n610) );
  NAND2_X1 U683 ( .A1(n647), .A2(G67), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U685 ( .A(KEYINPUT82), .B(n611), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G93), .A2(n637), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G80), .A2(n638), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n659) );
  XOR2_X1 U690 ( .A(n616), .B(n659), .Z(G145) );
  NAND2_X1 U691 ( .A1(n637), .A2(G86), .ZN(n617) );
  XOR2_X1 U692 ( .A(KEYINPUT83), .B(n617), .Z(n619) );
  NAND2_X1 U693 ( .A1(n647), .A2(G61), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U695 ( .A(KEYINPUT84), .B(n620), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n638), .A2(G73), .ZN(n621) );
  XOR2_X1 U697 ( .A(KEYINPUT2), .B(n621), .Z(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n643), .A2(G48), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT85), .B(n626), .Z(G305) );
  NAND2_X1 U702 ( .A1(G60), .A2(n647), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G47), .A2(n643), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G85), .A2(n637), .ZN(n629) );
  XOR2_X1 U706 ( .A(KEYINPUT66), .B(n629), .Z(n630) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n638), .A2(G72), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U710 ( .A1(G62), .A2(n647), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G50), .A2(n643), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U713 ( .A(KEYINPUT86), .B(n636), .ZN(n642) );
  NAND2_X1 U714 ( .A1(G88), .A2(n637), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G75), .A2(n638), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n642), .A2(n641), .ZN(G166) );
  NAND2_X1 U718 ( .A1(G49), .A2(n643), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n650), .A2(n649), .ZN(G288) );
  XNOR2_X1 U724 ( .A(n659), .B(G305), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n652) );
  XNOR2_X1 U726 ( .A(G290), .B(G166), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U728 ( .A(n653), .B(G288), .Z(n654) );
  XNOR2_X1 U729 ( .A(G299), .B(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n889) );
  XNOR2_X1 U731 ( .A(n657), .B(n889), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n658), .A2(G868), .ZN(n661) );
  OR2_X1 U733 ( .A1(G868), .A2(n659), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n661), .A2(n660), .ZN(G295) );
  XOR2_X1 U735 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n663) );
  NAND2_X1 U736 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n664), .A2(G2090), .ZN(n665) );
  XOR2_X1 U739 ( .A(KEYINPUT89), .B(n665), .Z(n666) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XOR2_X1 U742 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G108), .A2(G120), .ZN(n668) );
  NOR2_X1 U745 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(G69), .A2(n669), .ZN(n911) );
  NAND2_X1 U747 ( .A1(n911), .A2(G567), .ZN(n675) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U750 ( .A1(G218), .A2(n671), .ZN(n672) );
  XNOR2_X1 U751 ( .A(KEYINPUT90), .B(n672), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n673), .A2(G96), .ZN(n910) );
  NAND2_X1 U753 ( .A1(n910), .A2(G2106), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n675), .A2(n674), .ZN(n825) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n676) );
  XOR2_X1 U756 ( .A(KEYINPUT91), .B(n676), .Z(n677) );
  NOR2_X1 U757 ( .A1(n825), .A2(n677), .ZN(n824) );
  NAND2_X1 U758 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(G138), .A2(n678), .ZN(n680) );
  NAND2_X1 U760 ( .A1(G102), .A2(n878), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U762 ( .A1(G114), .A2(n873), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G126), .A2(n875), .ZN(n681) );
  NAND2_X1 U764 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U765 ( .A1(n684), .A2(n683), .ZN(G164) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n767) );
  AND2_X1 U768 ( .A1(n767), .A2(G40), .ZN(n685) );
  NOR2_X1 U769 ( .A1(G1966), .A2(n763), .ZN(n738) );
  NOR2_X1 U770 ( .A1(G2084), .A2(n728), .ZN(n739) );
  NOR2_X1 U771 ( .A1(n738), .A2(n739), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G8), .A2(n686), .ZN(n688) );
  NOR2_X1 U773 ( .A1(n689), .A2(G168), .ZN(n694) );
  XOR2_X1 U774 ( .A(G2078), .B(KEYINPUT25), .Z(n946) );
  NOR2_X1 U775 ( .A1(n946), .A2(n728), .ZN(n691) );
  INV_X1 U776 ( .A(n728), .ZN(n708) );
  NOR2_X1 U777 ( .A1(n708), .A2(G1961), .ZN(n690) );
  NOR2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U779 ( .A(KEYINPUT99), .B(n692), .ZN(n721) );
  NOR2_X1 U780 ( .A1(G171), .A2(n721), .ZN(n693) );
  XNOR2_X1 U781 ( .A(KEYINPUT31), .B(n695), .ZN(n696) );
  XNOR2_X1 U782 ( .A(n696), .B(KEYINPUT103), .ZN(n725) );
  NAND2_X1 U783 ( .A1(G1956), .A2(n728), .ZN(n697) );
  XNOR2_X1 U784 ( .A(KEYINPUT101), .B(n697), .ZN(n701) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(KEYINPUT100), .Z(n699) );
  NAND2_X1 U786 ( .A1(n708), .A2(G2072), .ZN(n698) );
  XOR2_X1 U787 ( .A(n699), .B(n698), .Z(n700) );
  NOR2_X1 U788 ( .A1(n701), .A2(n700), .ZN(n703) );
  NOR2_X1 U789 ( .A1(n971), .A2(n703), .ZN(n702) );
  XOR2_X1 U790 ( .A(n702), .B(KEYINPUT28), .Z(n719) );
  NAND2_X1 U791 ( .A1(n971), .A2(n703), .ZN(n717) );
  AND2_X1 U792 ( .A1(n708), .A2(G1996), .ZN(n704) );
  XOR2_X1 U793 ( .A(n704), .B(KEYINPUT26), .Z(n706) );
  NAND2_X1 U794 ( .A1(n728), .A2(G1341), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U796 ( .A1(n966), .A2(n707), .ZN(n712) );
  NAND2_X1 U797 ( .A1(G1348), .A2(n728), .ZN(n710) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n708), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n713) );
  NOR2_X1 U800 ( .A1(n961), .A2(n713), .ZN(n711) );
  OR2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n961), .A2(n713), .ZN(n714) );
  NAND2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U806 ( .A(KEYINPUT29), .B(n720), .Z(n723) );
  NAND2_X1 U807 ( .A1(G171), .A2(n721), .ZN(n722) );
  NAND2_X1 U808 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U809 ( .A1(n725), .A2(n724), .ZN(n736) );
  NAND2_X1 U810 ( .A1(n736), .A2(G286), .ZN(n727) );
  XNOR2_X1 U811 ( .A(n727), .B(n726), .ZN(n733) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n763), .ZN(n730) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U814 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U815 ( .A1(G303), .A2(n731), .ZN(n732) );
  NAND2_X1 U816 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U817 ( .A1(n734), .A2(G8), .ZN(n735) );
  XNOR2_X1 U818 ( .A(n735), .B(KEYINPUT32), .ZN(n744) );
  INV_X1 U819 ( .A(n736), .ZN(n737) );
  NOR2_X1 U820 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U821 ( .A1(G8), .A2(n739), .ZN(n740) );
  NAND2_X1 U822 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U823 ( .A(KEYINPUT104), .B(n742), .ZN(n743) );
  NAND2_X1 U824 ( .A1(n744), .A2(n743), .ZN(n751) );
  NOR2_X1 U825 ( .A1(G2090), .A2(G303), .ZN(n745) );
  NAND2_X1 U826 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U827 ( .A1(n751), .A2(n746), .ZN(n747) );
  XNOR2_X1 U828 ( .A(n747), .B(KEYINPUT106), .ZN(n748) );
  NAND2_X1 U829 ( .A1(n748), .A2(n763), .ZN(n749) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U832 ( .A1(n753), .A2(n750), .ZN(n970) );
  NAND2_X1 U833 ( .A1(n751), .A2(n970), .ZN(n757) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n969) );
  INV_X1 U835 ( .A(n969), .ZN(n752) );
  NAND2_X1 U836 ( .A1(n753), .A2(KEYINPUT33), .ZN(n754) );
  XOR2_X1 U837 ( .A(G1981), .B(G305), .Z(n977) );
  INV_X1 U838 ( .A(n977), .ZN(n755) );
  NOR2_X1 U839 ( .A1(n517), .A2(n755), .ZN(n758) );
  AND2_X1 U840 ( .A1(n518), .A2(n758), .ZN(n756) );
  AND2_X1 U841 ( .A1(n757), .A2(n756), .ZN(n760) );
  AND2_X1 U842 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U843 ( .A1(n760), .A2(n759), .ZN(n765) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XOR2_X1 U845 ( .A(n761), .B(KEYINPUT24), .Z(n762) );
  OR2_X1 U846 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U847 ( .A1(n765), .A2(n764), .ZN(n808) );
  NAND2_X1 U848 ( .A1(G160), .A2(G40), .ZN(n766) );
  NOR2_X1 U849 ( .A1(n767), .A2(n766), .ZN(n817) );
  NAND2_X1 U850 ( .A1(G140), .A2(n678), .ZN(n769) );
  NAND2_X1 U851 ( .A1(G104), .A2(n878), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U853 ( .A(KEYINPUT34), .B(n770), .ZN(n776) );
  NAND2_X1 U854 ( .A1(n873), .A2(G116), .ZN(n771) );
  XOR2_X1 U855 ( .A(KEYINPUT93), .B(n771), .Z(n773) );
  NAND2_X1 U856 ( .A1(n875), .A2(G128), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U858 ( .A(n774), .B(KEYINPUT35), .Z(n775) );
  NOR2_X1 U859 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U860 ( .A(KEYINPUT95), .B(n777), .Z(n779) );
  XOR2_X1 U861 ( .A(KEYINPUT36), .B(KEYINPUT94), .Z(n778) );
  XOR2_X1 U862 ( .A(n779), .B(n778), .Z(n863) );
  XOR2_X1 U863 ( .A(G2067), .B(KEYINPUT37), .Z(n780) );
  XOR2_X1 U864 ( .A(KEYINPUT92), .B(n780), .Z(n816) );
  NOR2_X1 U865 ( .A1(n863), .A2(n816), .ZN(n914) );
  NAND2_X1 U866 ( .A1(n817), .A2(n914), .ZN(n781) );
  XNOR2_X1 U867 ( .A(n781), .B(KEYINPUT96), .ZN(n809) );
  INV_X1 U868 ( .A(n809), .ZN(n806) );
  NAND2_X1 U869 ( .A1(G117), .A2(n873), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G129), .A2(n875), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n878), .A2(G105), .ZN(n784) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n678), .A2(G141), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n861) );
  NOR2_X1 U877 ( .A1(G1996), .A2(n861), .ZN(n929) );
  INV_X1 U878 ( .A(n817), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n861), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G119), .A2(n875), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G131), .A2(n678), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G107), .A2(n873), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G95), .A2(n878), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  OR2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n862) );
  NAND2_X1 U887 ( .A1(G1991), .A2(n862), .ZN(n795) );
  XOR2_X1 U888 ( .A(KEYINPUT97), .B(n795), .Z(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U890 ( .A(KEYINPUT98), .B(n798), .Z(n931) );
  NOR2_X1 U891 ( .A1(n799), .A2(n931), .ZN(n811) );
  NOR2_X1 U892 ( .A1(G1991), .A2(n862), .ZN(n925) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U894 ( .A1(n925), .A2(n800), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n811), .A2(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n929), .A2(n802), .ZN(n803) );
  XNOR2_X1 U897 ( .A(KEYINPUT39), .B(n803), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n804), .A2(n817), .ZN(n805) );
  OR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n814) );
  INV_X1 U900 ( .A(n814), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n520), .A2(n519), .ZN(n815) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n963) );
  NAND2_X1 U903 ( .A1(n963), .A2(n817), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n812) );
  OR2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n815), .A2(n516), .ZN(n819) );
  AND2_X1 U907 ( .A1(n863), .A2(n816), .ZN(n915) );
  NAND2_X1 U908 ( .A1(n915), .A2(n817), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U910 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U913 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U916 ( .A(n825), .ZN(G319) );
  XNOR2_X1 U917 ( .A(G1961), .B(KEYINPUT41), .ZN(n835) );
  XOR2_X1 U918 ( .A(G1956), .B(G1966), .Z(n827) );
  XNOR2_X1 U919 ( .A(G1981), .B(G1976), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U921 ( .A(G1971), .B(G1986), .Z(n829) );
  XNOR2_X1 U922 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U924 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U925 ( .A(G2474), .B(KEYINPUT112), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n835), .B(n834), .ZN(G229) );
  XOR2_X1 U928 ( .A(KEYINPUT111), .B(G2090), .Z(n837) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2084), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U931 ( .A(n838), .B(G2096), .Z(n840) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2072), .ZN(n839) );
  XNOR2_X1 U933 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U934 ( .A(G2678), .B(KEYINPUT43), .Z(n842) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2100), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U937 ( .A(n844), .B(n843), .Z(G227) );
  NAND2_X1 U938 ( .A1(G112), .A2(n873), .ZN(n846) );
  NAND2_X1 U939 ( .A1(G100), .A2(n878), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n846), .A2(n845), .ZN(n852) );
  NAND2_X1 U941 ( .A1(n875), .A2(G124), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U943 ( .A1(G136), .A2(n678), .ZN(n848) );
  NAND2_X1 U944 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U945 ( .A(KEYINPUT113), .B(n850), .Z(n851) );
  NOR2_X1 U946 ( .A1(n852), .A2(n851), .ZN(G162) );
  NAND2_X1 U947 ( .A1(G139), .A2(n678), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G103), .A2(n878), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U950 ( .A1(G115), .A2(n873), .ZN(n856) );
  NAND2_X1 U951 ( .A1(G127), .A2(n875), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U953 ( .A(KEYINPUT47), .B(n857), .Z(n858) );
  NOR2_X1 U954 ( .A1(n859), .A2(n858), .ZN(n916) );
  XOR2_X1 U955 ( .A(G160), .B(n916), .Z(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n867) );
  XNOR2_X1 U957 ( .A(n862), .B(G162), .ZN(n865) );
  XNOR2_X1 U958 ( .A(G164), .B(n863), .ZN(n864) );
  XNOR2_X1 U959 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U960 ( .A(n867), .B(n866), .ZN(n872) );
  XOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n869) );
  XNOR2_X1 U962 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U964 ( .A(n922), .B(n870), .ZN(n871) );
  XNOR2_X1 U965 ( .A(n872), .B(n871), .ZN(n887) );
  NAND2_X1 U966 ( .A1(n873), .A2(G118), .ZN(n874) );
  XNOR2_X1 U967 ( .A(n874), .B(KEYINPUT114), .ZN(n877) );
  NAND2_X1 U968 ( .A1(G130), .A2(n875), .ZN(n876) );
  NAND2_X1 U969 ( .A1(n877), .A2(n876), .ZN(n885) );
  NAND2_X1 U970 ( .A1(G106), .A2(n878), .ZN(n879) );
  XOR2_X1 U971 ( .A(KEYINPUT115), .B(n879), .Z(n881) );
  NAND2_X1 U972 ( .A1(n678), .A2(G142), .ZN(n880) );
  NAND2_X1 U973 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U974 ( .A(KEYINPUT116), .B(n882), .Z(n883) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n883), .ZN(n884) );
  NOR2_X1 U976 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U977 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U978 ( .A1(G37), .A2(n888), .ZN(G395) );
  XNOR2_X1 U979 ( .A(n889), .B(n966), .ZN(n890) );
  XNOR2_X1 U980 ( .A(n890), .B(G286), .ZN(n892) );
  XOR2_X1 U981 ( .A(n961), .B(G171), .Z(n891) );
  XNOR2_X1 U982 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U983 ( .A1(G37), .A2(n893), .ZN(G397) );
  XNOR2_X1 U984 ( .A(G2451), .B(G2443), .ZN(n903) );
  XOR2_X1 U985 ( .A(G2446), .B(G2454), .Z(n895) );
  XNOR2_X1 U986 ( .A(KEYINPUT109), .B(G2435), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U988 ( .A(KEYINPUT108), .B(G2438), .Z(n897) );
  XNOR2_X1 U989 ( .A(G1341), .B(G1348), .ZN(n896) );
  XNOR2_X1 U990 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U991 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U992 ( .A(G2430), .B(G2427), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U994 ( .A(n903), .B(n902), .ZN(n904) );
  NAND2_X1 U995 ( .A1(n904), .A2(G14), .ZN(n913) );
  NAND2_X1 U996 ( .A1(G319), .A2(n913), .ZN(n907) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n905) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U999 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(n909), .A2(n908), .ZN(G225) );
  XNOR2_X1 U1002 ( .A(KEYINPUT119), .B(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(G120), .ZN(G236) );
  INV_X1 U1005 ( .A(G108), .ZN(G238) );
  INV_X1 U1006 ( .A(G96), .ZN(G221) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n912), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U1010 ( .A(G325), .ZN(G261) );
  INV_X1 U1011 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1012 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1017) );
  INV_X1 U1013 ( .A(KEYINPUT55), .ZN(n937) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n927) );
  XOR2_X1 U1015 ( .A(G2072), .B(n916), .Z(n918) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT50), .B(n919), .Z(n921) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n934) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n930), .Z(n932) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n935), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1031 ( .A1(n938), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1032 ( .A(KEYINPUT121), .B(G2067), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(n939), .B(G26), .ZN(n950) );
  XNOR2_X1 U1034 ( .A(G1996), .B(G32), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n945) );
  XOR2_X1 U1037 ( .A(G1991), .B(G25), .Z(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(G28), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT120), .B(n943), .Z(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G27), .B(n946), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n951), .B(KEYINPUT53), .ZN(n954) );
  XOR2_X1 U1045 ( .A(G2084), .B(G34), .Z(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(n952), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G35), .B(G2090), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(n957), .Z(n958) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n958), .ZN(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT122), .B(n959), .Z(n960) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n960), .ZN(n1013) );
  XNOR2_X1 U1054 ( .A(G16), .B(KEYINPUT56), .ZN(n985) );
  XNOR2_X1 U1055 ( .A(G171), .B(G1961), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(G1348), .B(n961), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G1341), .B(n966), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n983) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n975) );
  XNOR2_X1 U1062 ( .A(G1956), .B(n971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n976), .B(KEYINPUT123), .ZN(n981) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1069 ( .A(KEYINPUT57), .B(n979), .Z(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n1011) );
  INV_X1 U1073 ( .A(G16), .ZN(n1009) );
  XOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .Z(n986) );
  XNOR2_X1 U1075 ( .A(G4), .B(n986), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G6), .B(G1981), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G1341), .B(G19), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G1956), .B(G20), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n993), .B(KEYINPUT125), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n994), .ZN(n1004) );
  XNOR2_X1 U1084 ( .A(G1961), .B(KEYINPUT124), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(G5), .ZN(n1002) );
  XNOR2_X1 U1086 ( .A(G1976), .B(G23), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n999) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(KEYINPUT58), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G21), .B(G1966), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(n1017), .B(n1016), .ZN(G150) );
  INV_X1 U1102 ( .A(G150), .ZN(G311) );
endmodule

