

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n390), .B(n294), .ZN(n295) );
  XNOR2_X1 U324 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U325 ( .A(KEYINPUT29), .B(n293), .ZN(n294) );
  XNOR2_X1 U326 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n406) );
  NOR2_X1 U327 ( .A1(n513), .A2(n425), .ZN(n564) );
  XNOR2_X1 U328 ( .A(n407), .B(n406), .ZN(n524) );
  XNOR2_X1 U329 ( .A(n301), .B(n300), .ZN(n303) );
  INV_X1 U330 ( .A(G183GAT), .ZN(n451) );
  XOR2_X1 U331 ( .A(n446), .B(n445), .Z(n517) );
  XOR2_X1 U332 ( .A(n462), .B(KEYINPUT28), .Z(n526) );
  XNOR2_X1 U333 ( .A(n451), .B(KEYINPUT120), .ZN(n452) );
  XNOR2_X1 U334 ( .A(n453), .B(n452), .ZN(G1350GAT) );
  XOR2_X1 U335 ( .A(G43GAT), .B(KEYINPUT8), .Z(n292) );
  XNOR2_X1 U336 ( .A(KEYINPUT66), .B(KEYINPUT7), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n390) );
  NAND2_X1 U338 ( .A1(G229GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U339 ( .A(G15GAT), .B(G22GAT), .Z(n363) );
  XNOR2_X1 U340 ( .A(n295), .B(n363), .ZN(n301) );
  XOR2_X1 U341 ( .A(KEYINPUT30), .B(G197GAT), .Z(n297) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G141GAT), .ZN(n296) );
  XOR2_X1 U343 ( .A(n297), .B(n296), .Z(n299) );
  XNOR2_X1 U344 ( .A(G50GAT), .B(G29GAT), .ZN(n298) );
  XOR2_X1 U345 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  XOR2_X1 U346 ( .A(G113GAT), .B(G1GAT), .Z(n341) );
  XNOR2_X1 U347 ( .A(n413), .B(n341), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n566) );
  XOR2_X1 U349 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n305) );
  XNOR2_X1 U350 ( .A(KEYINPUT23), .B(KEYINPUT85), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n307) );
  XNOR2_X1 U353 ( .A(G22GAT), .B(KEYINPUT84), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(n309), .B(n308), .Z(n319) );
  XOR2_X1 U356 ( .A(G148GAT), .B(G106GAT), .Z(n311) );
  XNOR2_X1 U357 ( .A(G204GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(KEYINPUT67), .B(n312), .Z(n356) );
  XOR2_X1 U360 ( .A(G50GAT), .B(G162GAT), .Z(n380) );
  XOR2_X1 U361 ( .A(G211GAT), .B(KEYINPUT21), .Z(n314) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n421) );
  XOR2_X1 U364 ( .A(n380), .B(n421), .Z(n316) );
  NAND2_X1 U365 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n356), .B(n317), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U369 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n321) );
  XNOR2_X1 U370 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(n322), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n323), .B(n324), .ZN(n462) );
  INV_X1 U374 ( .A(n324), .ZN(n331) );
  XOR2_X1 U375 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n326) );
  XNOR2_X1 U376 ( .A(G162GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(n327), .B(KEYINPUT90), .Z(n329) );
  XOR2_X1 U379 ( .A(G120GAT), .B(G57GAT), .Z(n349) );
  XNOR2_X1 U380 ( .A(G148GAT), .B(n349), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n345) );
  XOR2_X1 U383 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n333) );
  XNOR2_X1 U384 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U386 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n335) );
  XNOR2_X1 U387 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(n337), .B(n336), .Z(n343) );
  XOR2_X1 U390 ( .A(G29GAT), .B(G134GAT), .Z(n379) );
  XOR2_X1 U391 ( .A(KEYINPUT0), .B(G127GAT), .Z(n438) );
  XOR2_X1 U392 ( .A(n379), .B(n438), .Z(n339) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n469) );
  XNOR2_X1 U398 ( .A(KEYINPUT95), .B(n469), .ZN(n513) );
  XOR2_X1 U399 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n351) );
  XOR2_X1 U400 ( .A(KEYINPUT69), .B(G92GAT), .Z(n347) );
  XNOR2_X1 U401 ( .A(G99GAT), .B(KEYINPUT68), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U403 ( .A(G85GAT), .B(n348), .Z(n398) );
  XNOR2_X1 U404 ( .A(n349), .B(n398), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U406 ( .A(G71GAT), .B(KEYINPUT13), .Z(n362) );
  XOR2_X1 U407 ( .A(KEYINPUT32), .B(n362), .Z(n353) );
  NAND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XOR2_X1 U409 ( .A(n353), .B(n352), .Z(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n358) );
  XOR2_X1 U411 ( .A(G176GAT), .B(G64GAT), .Z(n410) );
  XNOR2_X1 U412 ( .A(n356), .B(n410), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n569) );
  XNOR2_X1 U414 ( .A(n569), .B(KEYINPUT41), .ZN(n499) );
  NOR2_X1 U415 ( .A1(n566), .A2(n499), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n359), .B(KEYINPUT46), .ZN(n378) );
  XOR2_X1 U417 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n361) );
  XNOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n367) );
  XOR2_X1 U420 ( .A(n362), .B(G127GAT), .Z(n365) );
  XNOR2_X1 U421 ( .A(n363), .B(G183GAT), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U423 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n377) );
  XOR2_X1 U426 ( .A(G211GAT), .B(G78GAT), .Z(n371) );
  XNOR2_X1 U427 ( .A(G8GAT), .B(G155GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U429 ( .A(KEYINPUT77), .B(G64GAT), .Z(n373) );
  XNOR2_X1 U430 ( .A(G1GAT), .B(G57GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n455) );
  NOR2_X1 U434 ( .A1(n378), .A2(n455), .ZN(n399) );
  XOR2_X1 U435 ( .A(KEYINPUT10), .B(n379), .Z(n382) );
  XNOR2_X1 U436 ( .A(n380), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n394) );
  XOR2_X1 U438 ( .A(KEYINPUT74), .B(KEYINPUT72), .Z(n384) );
  XNOR2_X1 U439 ( .A(KEYINPUT65), .B(KEYINPUT73), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT71), .Z(n386) );
  XNOR2_X1 U442 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U444 ( .A(n388), .B(n387), .Z(n392) );
  XNOR2_X1 U445 ( .A(G36GAT), .B(G190GAT), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n389), .B(KEYINPUT75), .ZN(n417) );
  XNOR2_X1 U447 ( .A(n390), .B(n417), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U449 ( .A(n394), .B(n393), .Z(n396) );
  NAND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n557) );
  NAND2_X1 U453 ( .A1(n399), .A2(n557), .ZN(n400) );
  XNOR2_X1 U454 ( .A(n400), .B(KEYINPUT47), .ZN(n405) );
  XNOR2_X1 U455 ( .A(KEYINPUT36), .B(n557), .ZN(n581) );
  INV_X1 U456 ( .A(n455), .ZN(n575) );
  NOR2_X1 U457 ( .A1(n581), .A2(n575), .ZN(n401) );
  XNOR2_X1 U458 ( .A(KEYINPUT45), .B(n401), .ZN(n402) );
  NAND2_X1 U459 ( .A1(n402), .A2(n566), .ZN(n403) );
  NOR2_X1 U460 ( .A1(n403), .A2(n569), .ZN(n404) );
  NOR2_X1 U461 ( .A1(n405), .A2(n404), .ZN(n407) );
  XOR2_X1 U462 ( .A(G183GAT), .B(KEYINPUT17), .Z(n409) );
  XNOR2_X1 U463 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n437) );
  XNOR2_X1 U465 ( .A(G204GAT), .B(G92GAT), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U467 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U470 ( .A(n416), .B(KEYINPUT97), .Z(n419) );
  XNOR2_X1 U471 ( .A(n417), .B(KEYINPUT96), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n437), .B(n420), .ZN(n423) );
  INV_X1 U474 ( .A(n421), .ZN(n422) );
  XOR2_X1 U475 ( .A(n423), .B(n422), .Z(n515) );
  INV_X1 U476 ( .A(n515), .ZN(n457) );
  NOR2_X1 U477 ( .A1(n524), .A2(n457), .ZN(n424) );
  XOR2_X1 U478 ( .A(KEYINPUT54), .B(n424), .Z(n425) );
  NAND2_X1 U479 ( .A1(n462), .A2(n564), .ZN(n426) );
  XNOR2_X1 U480 ( .A(KEYINPUT55), .B(n426), .ZN(n447) );
  XOR2_X1 U481 ( .A(G176GAT), .B(KEYINPUT78), .Z(n428) );
  XNOR2_X1 U482 ( .A(G169GAT), .B(G15GAT), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n446) );
  XOR2_X1 U484 ( .A(G190GAT), .B(G134GAT), .Z(n430) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G99GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n432) );
  XNOR2_X1 U488 ( .A(G113GAT), .B(G120GAT), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U490 ( .A(n434), .B(n433), .Z(n444) );
  XOR2_X1 U491 ( .A(G71GAT), .B(KEYINPUT82), .Z(n436) );
  XNOR2_X1 U492 ( .A(KEYINPUT81), .B(KEYINPUT20), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n442) );
  XOR2_X1 U494 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U499 ( .A1(n447), .A2(n517), .ZN(n556) );
  NOR2_X1 U500 ( .A1(n566), .A2(n556), .ZN(n450) );
  INV_X1 U501 ( .A(G169GAT), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n448), .B(KEYINPUT118), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(G1348GAT) );
  NOR2_X1 U504 ( .A1(n575), .A2(n556), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n475) );
  NOR2_X1 U506 ( .A1(n566), .A2(n569), .ZN(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT70), .B(n454), .Z(n486) );
  NAND2_X1 U508 ( .A1(n557), .A2(n455), .ZN(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT16), .B(n456), .Z(n473) );
  XOR2_X1 U510 ( .A(KEYINPUT27), .B(n457), .Z(n461) );
  NAND2_X1 U511 ( .A1(n513), .A2(n461), .ZN(n523) );
  NOR2_X1 U512 ( .A1(n526), .A2(n523), .ZN(n458) );
  INV_X1 U513 ( .A(n517), .ZN(n525) );
  NAND2_X1 U514 ( .A1(n458), .A2(n525), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT98), .ZN(n472) );
  NOR2_X1 U516 ( .A1(n462), .A2(n517), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U518 ( .A1(n461), .A2(n563), .ZN(n468) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(KEYINPUT100), .ZN(n466) );
  NAND2_X1 U520 ( .A1(n515), .A2(n517), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT99), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n483) );
  NAND2_X1 U527 ( .A1(n473), .A2(n483), .ZN(n500) );
  NOR2_X1 U528 ( .A1(n486), .A2(n500), .ZN(n481) );
  NAND2_X1 U529 ( .A1(n481), .A2(n513), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U532 ( .A1(n481), .A2(n515), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n479) );
  NAND2_X1 U535 ( .A1(n481), .A2(n517), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U538 ( .A1(n481), .A2(n526), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U540 ( .A1(n575), .A2(n483), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n581), .A2(n484), .ZN(n485) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n485), .ZN(n511) );
  NOR2_X1 U543 ( .A1(n511), .A2(n486), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n487), .B(KEYINPUT38), .ZN(n497) );
  NAND2_X1 U545 ( .A1(n497), .A2(n513), .ZN(n490) );
  XNOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U549 ( .A1(n497), .A2(n515), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n496) );
  XOR2_X1 U553 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n494) );
  NAND2_X1 U554 ( .A1(n517), .A2(n497), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n497), .A2(n526), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n503) );
  INV_X1 U560 ( .A(n499), .ZN(n530) );
  NAND2_X1 U561 ( .A1(n566), .A2(n530), .ZN(n510) );
  NOR2_X1 U562 ( .A1(n500), .A2(n510), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT108), .ZN(n507) );
  NAND2_X1 U564 ( .A1(n507), .A2(n513), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n507), .A2(n515), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n507), .A2(n517), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U572 ( .A1(n526), .A2(n507), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NOR2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U575 ( .A(KEYINPUT109), .B(n512), .Z(n519) );
  NAND2_X1 U576 ( .A1(n519), .A2(n513), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n519), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n519), .A2(n517), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n521) );
  NAND2_X1 U583 ( .A1(n519), .A2(n526), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n522), .Z(G1339GAT) );
  NOR2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n539) );
  NOR2_X1 U587 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n539), .A2(n527), .ZN(n535) );
  NOR2_X1 U589 ( .A1(n566), .A2(n535), .ZN(n529) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT111), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  NOR2_X1 U592 ( .A1(n499), .A2(n535), .ZN(n532) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U595 ( .A1(n575), .A2(n535), .ZN(n533) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(n533), .Z(n534) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U598 ( .A1(n557), .A2(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(KEYINPUT112), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U602 ( .A1(n539), .A2(n563), .ZN(n549) );
  NOR2_X1 U603 ( .A1(n566), .A2(n549), .ZN(n541) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(KEYINPUT113), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n543) );
  XNOR2_X1 U607 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n547) );
  NOR2_X1 U609 ( .A1(n499), .A2(n549), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n575), .A2(n549), .ZN(n548) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n557), .A2(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NOR2_X1 U618 ( .A1(n556), .A2(n499), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  INV_X1 U623 ( .A(KEYINPUT58), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n562) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT121), .B(n565), .Z(n580) );
  NOR2_X1 U632 ( .A1(n566), .A2(n580), .ZN(n567) );
  XOR2_X1 U633 ( .A(n568), .B(n567), .Z(G1352GAT) );
  INV_X1 U634 ( .A(n569), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n580), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n580), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

