//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT99), .B(G92gat), .Z(new_n203));
  INV_X1    g002(.A(G85gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n203), .A2(new_n204), .B1(KEYINPUT8), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n205), .ZN(new_n207));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G92gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(new_n204), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(G85gat), .A3(G92gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n209), .A2(KEYINPUT100), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n207), .A2(new_n208), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT100), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n206), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n205), .A2(KEYINPUT8), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT99), .B(G92gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G85gat), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n211), .A2(new_n213), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n216), .B(new_n215), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G29gat), .A2(G36gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NOR3_X1   g026(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(KEYINPUT15), .A3(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n230), .A2(KEYINPUT15), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(KEYINPUT15), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(G36gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n228), .A2(KEYINPUT91), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n227), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n231), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT17), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(new_n231), .C1(new_n234), .C2(new_n239), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n224), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n224), .ZN(new_n247));
  AND2_X1   g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT41), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(G190gat), .B1(new_n244), .B2(new_n250), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G218gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n202), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n248), .A2(KEYINPUT41), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n252), .A2(G218gat), .A3(new_n253), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G134gat), .B(G162gat), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n256), .B2(new_n259), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n254), .A2(new_n255), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT98), .A3(new_n259), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n257), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n262), .B1(new_n268), .B2(new_n260), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G71gat), .A2(G78gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(G71gat), .A2(G78gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(KEYINPUT95), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(KEYINPUT95), .B2(new_n271), .ZN(new_n274));
  INV_X1    g073(.A(G64gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G57gat), .ZN(new_n276));
  INV_X1    g075(.A(G57gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G64gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n279), .A2(KEYINPUT96), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT9), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n279), .A2(KEYINPUT96), .B1(new_n281), .B2(new_n271), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n274), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(KEYINPUT97), .A3(G57gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n278), .ZN(new_n287));
  OR2_X1    g086(.A1(G71gat), .A2(G78gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n271), .B1(new_n288), .B2(new_n281), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT21), .ZN(new_n292));
  AND2_X1   g091(.A1(G231gat), .A2(G233gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G127gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT92), .ZN(new_n297));
  XOR2_X1   g096(.A(G15gat), .B(G22gat), .Z(new_n298));
  INV_X1    g097(.A(G1gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G15gat), .B(G22gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT16), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(G1gat), .ZN(new_n303));
  INV_X1    g102(.A(G8gat), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n300), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n297), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(new_n303), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G8gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT92), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(KEYINPUT21), .B2(new_n291), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n296), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G183gat), .B(G211gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n296), .A2(new_n313), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n296), .A2(new_n313), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G230gat), .A2(G233gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n291), .A2(new_n224), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n218), .B(new_n223), .C1(new_n283), .C2(new_n290), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(KEYINPUT101), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT101), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n291), .A2(new_n224), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT10), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT10), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n326), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n326), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n336), .A3(new_n331), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G120gat), .B(G148gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT102), .ZN(new_n340));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n335), .A2(new_n337), .A3(new_n342), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n270), .A2(new_n325), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(G183gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n246), .ZN(new_n354));
  NAND3_X1  g153(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT66), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n356), .A2(KEYINPUT66), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n354), .B(new_n355), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT65), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(G169gat), .B2(G176gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(KEYINPUT23), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n367));
  NAND2_X1  g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT23), .ZN(new_n369));
  INV_X1    g168(.A(G169gat), .ZN(new_n370));
  INV_X1    g169(.A(G176gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n367), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n358), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n354), .A3(new_n355), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n372), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT64), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n362), .A2(new_n378), .A3(KEYINPUT23), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n362), .B2(KEYINPUT23), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n376), .B(new_n377), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n361), .A2(new_n374), .B1(new_n381), .B2(new_n367), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT26), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n363), .A2(new_n383), .A3(new_n365), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n372), .A2(KEYINPUT26), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n368), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n353), .A2(KEYINPUT27), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G183gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n389), .A3(new_n246), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n390), .A2(new_n391), .B1(G183gat), .B2(G190gat), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n386), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n352), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397));
  XNOR2_X1  g196(.A(G197gat), .B(G204gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(G211gat), .A2(G218gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(KEYINPUT74), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(KEYINPUT74), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT75), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G211gat), .B(G218gat), .Z(new_n406));
  OR2_X1    g205(.A1(new_n403), .A2(KEYINPUT74), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT75), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n401), .A4(new_n398), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n405), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n397), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(new_n406), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n374), .A2(new_n361), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n381), .A2(new_n367), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n386), .A2(new_n392), .A3(new_n393), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n352), .B(KEYINPUT77), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n396), .A2(new_n418), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n424), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n395), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(G226gat), .A3(G233gat), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n418), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n351), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n424), .B1(new_n423), .B2(new_n428), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n395), .A2(new_n352), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n417), .B(new_n412), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n396), .A2(new_n418), .A3(new_n425), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n350), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n436), .A2(new_n440), .A3(new_n437), .A4(new_n350), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(G1gat), .B(G29gat), .Z(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n447), .A2(KEYINPUT6), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n452));
  INV_X1    g251(.A(G113gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT69), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G113gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(G120gat), .ZN(new_n457));
  INV_X1    g256(.A(G120gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G113gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(KEYINPUT70), .A3(new_n459), .ZN(new_n463));
  INV_X1    g262(.A(G134gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n295), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G127gat), .A2(G134gat), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT1), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT68), .B(G127gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n469), .B2(new_n464), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n453), .A2(G120gat), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT1), .B1(new_n459), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT2), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n476), .A2(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G141gat), .B(G148gat), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(G155gat), .B2(G162gat), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(G141gat), .A2(G148gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G162gat), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT2), .B1(new_n316), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n316), .B2(new_n484), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n483), .B(new_n485), .C1(new_n474), .C2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n473), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n488), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT3), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n480), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n470), .A2(new_n472), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n465), .A2(new_n466), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT1), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n460), .B2(new_n461), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n500), .B2(new_n463), .ZN(new_n501));
  OAI211_X1 g300(.A(KEYINPUT4), .B(new_n490), .C1(new_n495), .C2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n468), .A2(new_n473), .A3(new_n489), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G225gat), .A2(G233gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n452), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n507), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n489), .B1(new_n468), .B2(new_n473), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT80), .ZN(new_n512));
  INV_X1    g311(.A(new_n459), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT69), .B(G113gat), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(G120gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n467), .B1(new_n515), .B2(KEYINPUT70), .ZN(new_n516));
  INV_X1    g315(.A(new_n463), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n473), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n491), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n490), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n509), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n507), .A3(new_n452), .ZN(new_n525));
  AOI211_X1 g324(.A(new_n450), .B(new_n451), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AND4_X1   g325(.A1(new_n449), .A2(new_n524), .A3(new_n525), .A4(new_n448), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n442), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n518), .A2(new_n421), .A3(new_n422), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n501), .B1(new_n382), .B2(new_n394), .ZN(new_n530));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G71gat), .B(G99gat), .Z(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G43gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT33), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n529), .A2(new_n530), .A3(new_n532), .A4(new_n536), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT71), .B1(new_n540), .B2(new_n537), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n529), .A2(new_n530), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT34), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n531), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n532), .B1(new_n529), .B2(new_n530), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G78gat), .B(G106gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT31), .B(G50gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G22gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(new_n555), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT29), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n491), .B1(new_n560), .B2(KEYINPUT3), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n494), .A2(new_n428), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n412), .A2(new_n417), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n561), .A2(new_n563), .A3(G228gat), .A4(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G228gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT83), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n410), .A2(new_n411), .A3(new_n429), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n491), .B1(new_n569), .B2(KEYINPUT3), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n570), .B2(new_n563), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n559), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n550), .B(new_n539), .C1(new_n542), .C2(new_n541), .ZN(new_n573));
  INV_X1    g372(.A(new_n571), .ZN(new_n574));
  INV_X1    g373(.A(new_n559), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n564), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n552), .A2(new_n572), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT35), .B1(new_n528), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT90), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n512), .A2(new_n522), .ZN(new_n581));
  INV_X1    g380(.A(new_n452), .ZN(new_n582));
  AND4_X1   g381(.A1(new_n504), .A2(new_n468), .A3(new_n473), .A4(new_n489), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n504), .B1(new_n501), .B2(new_n489), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n518), .A2(new_n492), .A3(new_n494), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n582), .B1(new_n586), .B2(new_n509), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n525), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n450), .ZN(new_n589));
  INV_X1    g388(.A(new_n451), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n524), .A2(new_n449), .A3(new_n525), .A4(new_n448), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n572), .A2(new_n594), .A3(new_n576), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n593), .A2(new_n595), .A3(new_n442), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n552), .A2(KEYINPUT73), .A3(new_n573), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n543), .A2(new_n551), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(KEYINPUT89), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n599), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT89), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n596), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(KEYINPUT90), .B(KEYINPUT35), .C1(new_n528), .C2(new_n577), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n572), .A2(KEYINPUT85), .A3(new_n576), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT85), .B1(new_n572), .B2(new_n576), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n597), .A2(new_n610), .A3(new_n599), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n552), .A2(KEYINPUT36), .A3(new_n573), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n609), .A2(new_n528), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n520), .A2(new_n509), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n586), .A2(new_n509), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n502), .A2(new_n505), .A3(new_n615), .A4(new_n509), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT86), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n447), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n619), .B2(new_n447), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n618), .B(KEYINPUT40), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT88), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n621), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(KEYINPUT88), .A3(KEYINPUT40), .A4(new_n618), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n447), .B1(new_n524), .B2(new_n525), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n442), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n618), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(KEYINPUT87), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT87), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n627), .A2(new_n621), .B1(new_n617), .B2(new_n616), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(KEYINPUT40), .ZN(new_n638));
  AND4_X1   g437(.A1(new_n630), .A2(new_n632), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n572), .A2(new_n576), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n351), .A2(KEYINPUT37), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n433), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n418), .B1(new_n434), .B2(new_n435), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n396), .A2(new_n425), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n643), .B(KEYINPUT37), .C1(new_n418), .C2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n436), .A2(new_n437), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n433), .A2(new_n641), .B1(new_n648), .B2(KEYINPUT37), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n647), .B(new_n438), .C1(new_n649), .C2(new_n646), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n640), .B1(new_n650), .B2(new_n593), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n613), .B1(new_n639), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n606), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n239), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n655), .A2(new_n225), .A3(new_n233), .A4(new_n232), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n242), .B1(new_n656), .B2(new_n231), .ZN(new_n657));
  INV_X1    g456(.A(new_n243), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n309), .B(new_n310), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT93), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n312), .A2(new_n660), .A3(new_n240), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n312), .B2(new_n240), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n654), .B(new_n659), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n312), .A2(new_n240), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n312), .A2(new_n660), .A3(new_n240), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n669), .A2(KEYINPUT18), .A3(new_n654), .A4(new_n659), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n661), .A2(new_n662), .B1(new_n240), .B2(new_n312), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n654), .B(KEYINPUT13), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G113gat), .B(G141gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G197gat), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT11), .B(G169gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT12), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n670), .A3(new_n673), .A4(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n653), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT94), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n653), .A2(KEYINPUT94), .A3(new_n683), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n347), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n593), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  INV_X1    g491(.A(new_n442), .ZN(new_n693));
  INV_X1    g492(.A(new_n347), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n692), .A2(KEYINPUT103), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT94), .B1(new_n653), .B2(new_n683), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n681), .A2(new_n682), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n685), .B(new_n697), .C1(new_n606), .C2(new_n652), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n693), .B(new_n694), .C1(new_n696), .C2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n695), .A2(new_n701), .A3(G8gat), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n688), .A2(KEYINPUT42), .A3(new_n693), .A4(new_n703), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT42), .B1(new_n702), .B2(new_n703), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n707), .A2(new_n708), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(G1325gat));
  INV_X1    g514(.A(G15gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n603), .A2(new_n600), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n688), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n611), .A2(new_n612), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n688), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n723), .B2(new_n716), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n688), .A2(new_n609), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT43), .B(G22gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  INV_X1    g526(.A(new_n325), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n263), .B1(new_n261), .B2(new_n264), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n268), .A2(new_n262), .A3(new_n260), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n731), .A3(new_n346), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n692), .A2(new_n733), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n734), .A2(G29gat), .A3(new_n593), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n270), .B1(new_n606), .B2(new_n652), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(KEYINPUT107), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n270), .B(new_n741), .C1(new_n606), .C2(new_n652), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n325), .B(KEYINPUT106), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n344), .A2(new_n345), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(new_n697), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n689), .A3(new_n746), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n735), .A2(new_n736), .B1(G29gat), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n736), .B2(new_n735), .ZN(G1328gat));
  OR3_X1    g548(.A1(new_n734), .A2(G36gat), .A3(new_n442), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n743), .A2(new_n693), .A3(new_n746), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n750), .A2(KEYINPUT46), .B1(G36gat), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(KEYINPUT46), .B2(new_n750), .ZN(G1329gat));
  INV_X1    g552(.A(G43gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n734), .B2(new_n717), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n743), .A2(G43gat), .A3(new_n721), .A4(new_n746), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  INV_X1    g558(.A(G50gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n692), .A2(new_n760), .A3(new_n609), .A4(new_n733), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT48), .ZN(new_n762));
  INV_X1    g561(.A(new_n640), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n763), .B(new_n746), .C1(new_n739), .C2(new_n742), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n609), .B(new_n746), .C1(new_n739), .C2(new_n742), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G50gat), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n761), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n759), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n771), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n766), .A2(new_n767), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n773), .B(KEYINPUT109), .C1(new_n774), .C2(new_n762), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(G1331gat));
  NOR4_X1   g575(.A1(new_n728), .A2(new_n731), .A3(new_n683), .A4(new_n346), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n653), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n689), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g579(.A1(new_n778), .A2(new_n693), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  NAND2_X1  g584(.A1(new_n778), .A2(new_n721), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n717), .A2(G71gat), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n786), .A2(G71gat), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n778), .A2(new_n609), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n325), .A2(new_n683), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n737), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n794));
  NOR2_X1   g593(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n794), .B1(new_n737), .B2(new_n792), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(new_n745), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n204), .A3(new_n689), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n325), .A2(new_n683), .A3(new_n346), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n743), .A2(new_n689), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n204), .B2(new_n804), .ZN(G1336gat));
  NAND3_X1  g604(.A1(new_n743), .A2(new_n693), .A3(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n693), .A2(new_n745), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n806), .A2(new_n220), .B1(new_n799), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n809), .B(KEYINPUT52), .Z(G1337gat));
  INV_X1    g609(.A(G99gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n800), .A2(new_n811), .A3(new_n718), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n743), .A2(new_n721), .A3(new_n802), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G99gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n814), .B2(new_n816), .ZN(G1338gat));
  NOR2_X1   g616(.A1(new_n640), .A2(G106gat), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n745), .B(new_n818), .C1(new_n797), .C2(new_n798), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n609), .B(new_n802), .C1(new_n739), .C2(new_n742), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT53), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n822), .B2(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n743), .A2(new_n763), .A3(new_n802), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT53), .B1(new_n826), .B2(G106gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n819), .A2(KEYINPUT113), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n819), .A2(KEYINPUT113), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n824), .A2(new_n825), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  NOR2_X1   g630(.A1(new_n347), .A2(new_n683), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n343), .B1(new_n335), .B2(KEYINPUT54), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n329), .A2(new_n331), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n334), .B1(new_n835), .B2(new_n333), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n336), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(KEYINPUT54), .A3(new_n335), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n837), .A2(new_n840), .A3(KEYINPUT54), .A4(new_n335), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n834), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n345), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n833), .B1(new_n847), .B2(new_n841), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(KEYINPUT55), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n654), .B1(new_n669), .B2(new_n659), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n312), .A2(new_n240), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n851), .B(new_n672), .C1(new_n667), .C2(new_n668), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n678), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n682), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n731), .A2(new_n845), .A3(new_n849), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n682), .A2(new_n853), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n346), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n697), .B1(new_n843), .B2(new_n844), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n849), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n855), .B1(new_n859), .B2(new_n731), .ZN(new_n860));
  INV_X1    g659(.A(new_n744), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n832), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n593), .ZN(new_n863));
  INV_X1    g662(.A(new_n577), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n693), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n514), .A3(new_n683), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n860), .A2(new_n861), .ZN(new_n869));
  INV_X1    g668(.A(new_n832), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n609), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n862), .A2(KEYINPUT115), .A3(new_n609), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n693), .A2(new_n593), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n718), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n697), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n867), .B1(new_n878), .B2(new_n453), .ZN(G1340gat));
  AOI21_X1  g678(.A(G120gat), .B1(new_n866), .B2(new_n745), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n875), .A2(new_n877), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n346), .A2(new_n458), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(G1341gat));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n469), .A3(new_n325), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n875), .A2(new_n861), .A3(new_n877), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n469), .ZN(G1342gat));
  NAND2_X1  g685(.A1(new_n731), .A2(new_n442), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT116), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n865), .A2(G134gat), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT56), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n875), .A2(new_n270), .A3(new_n877), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n464), .B2(new_n891), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n721), .A2(new_n640), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT55), .B(new_n834), .C1(new_n839), .C2(new_n842), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n345), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n683), .B1(new_n848), .B2(KEYINPUT55), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n270), .B1(new_n897), .B2(new_n857), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n744), .B1(new_n898), .B2(new_n855), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n689), .B(new_n893), .C1(new_n899), .C2(new_n832), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n697), .A2(G141gat), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(new_n693), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n854), .A2(KEYINPUT117), .A3(new_n745), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n346), .B2(new_n856), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n858), .B2(new_n849), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n855), .B1(new_n907), .B2(new_n731), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n832), .B1(new_n908), .B2(new_n728), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n872), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n763), .C1(new_n899), .C2(new_n832), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n720), .A2(new_n876), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n910), .A2(new_n912), .A3(new_n683), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n902), .B1(new_n914), .B2(G141gat), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT118), .B1(new_n914), .B2(G141gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT58), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  AOI221_X4 g717(.A(new_n902), .B1(KEYINPUT118), .B2(new_n918), .C1(G141gat), .C2(new_n914), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n919), .ZN(G1344gat));
  OAI21_X1  g719(.A(KEYINPUT57), .B1(new_n862), .B2(new_n640), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n270), .B1(new_n897), .B2(new_n906), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n325), .B1(new_n922), .B2(new_n855), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n911), .B(new_n609), .C1(new_n923), .C2(new_n832), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n913), .A2(new_n745), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G148gat), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n912), .A3(new_n745), .A4(new_n913), .ZN(new_n928));
  INV_X1    g727(.A(G148gat), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(KEYINPUT59), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n927), .A2(KEYINPUT59), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n863), .A2(new_n442), .A3(new_n893), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n745), .A2(new_n929), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT119), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n936));
  INV_X1    g735(.A(new_n934), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n928), .A2(new_n930), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n926), .B2(G148gat), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n936), .B(new_n937), .C1(new_n938), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n935), .A2(new_n941), .ZN(G1345gat));
  NAND3_X1  g741(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n316), .A3(new_n861), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n932), .A2(new_n728), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n945), .A2(KEYINPUT120), .ZN(new_n946));
  AOI21_X1  g745(.A(G155gat), .B1(new_n945), .B2(KEYINPUT120), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1346gat));
  NAND4_X1  g747(.A1(new_n910), .A2(new_n912), .A3(new_n731), .A4(new_n913), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G162gat), .ZN(new_n950));
  OR3_X1    g749(.A1(new_n900), .A2(G162gat), .A3(new_n888), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(G1347gat));
  NOR2_X1   g753(.A1(new_n862), .A2(new_n689), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n864), .A2(new_n693), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT122), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(KEYINPUT123), .A3(new_n957), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n960), .A2(new_n370), .A3(new_n683), .A4(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n689), .A2(new_n442), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n966), .A2(new_n717), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT115), .B1(new_n862), .B2(new_n609), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n868), .B(new_n872), .C1(new_n899), .C2(new_n832), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(new_n683), .ZN(new_n972));
  OAI22_X1  g771(.A1(new_n963), .A2(new_n964), .B1(new_n370), .B2(new_n972), .ZN(G1348gat));
  NAND3_X1  g772(.A1(new_n960), .A2(new_n745), .A3(new_n961), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n974), .A2(new_n371), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n971), .A2(G176gat), .A3(new_n745), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(G1349gat));
  AOI21_X1  g779(.A(new_n353), .B1(new_n971), .B2(new_n744), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n387), .A2(new_n389), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n958), .A2(new_n983), .A3(new_n728), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n981), .A2(KEYINPUT60), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(KEYINPUT60), .B1(new_n981), .B2(new_n984), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1350gat));
  AOI211_X1 g786(.A(new_n270), .B(new_n968), .C1(new_n969), .C2(new_n970), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT126), .B1(new_n988), .B2(new_n246), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n731), .B(new_n967), .C1(new_n873), .C2(new_n874), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n990), .A2(new_n991), .A3(G190gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n989), .A2(KEYINPUT61), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n994));
  OAI211_X1 g793(.A(KEYINPUT126), .B(new_n994), .C1(new_n988), .C2(new_n246), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n960), .A2(new_n246), .A3(new_n731), .A4(new_n961), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(G1351gat));
  AND2_X1   g796(.A1(new_n921), .A2(new_n924), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n966), .A2(new_n721), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(G197gat), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n1000), .A2(new_n1001), .A3(new_n697), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n955), .A2(new_n893), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1003), .A2(new_n442), .ZN(new_n1004));
  AOI21_X1  g803(.A(G197gat), .B1(new_n1004), .B2(new_n683), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1002), .A2(new_n1005), .ZN(G1352gat));
  INV_X1    g805(.A(G204gat), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1007), .B1(new_n1008), .B2(KEYINPUT127), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n1003), .A2(new_n807), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(KEYINPUT127), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g811(.A(G204gat), .B1(new_n1000), .B2(new_n346), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(new_n1013), .ZN(G1353gat));
  INV_X1    g813(.A(G211gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1004), .A2(new_n1015), .A3(new_n325), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n325), .A3(new_n999), .ZN(new_n1017));
  AND3_X1   g816(.A1(new_n1017), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1018));
  AOI21_X1  g817(.A(KEYINPUT63), .B1(new_n1017), .B2(G211gat), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(G1354gat));
  OAI21_X1  g819(.A(G218gat), .B1(new_n1000), .B2(new_n270), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1004), .A2(new_n255), .A3(new_n731), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1021), .A2(new_n1022), .ZN(G1355gat));
endmodule


