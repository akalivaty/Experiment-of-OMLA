//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n192));
  AOI22_X1  g006(.A1(KEYINPUT66), .A2(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n196));
  OAI211_X1 g010(.A(G134), .B(new_n189), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n189), .B2(G134), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n193), .A2(new_n194), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT67), .B1(new_n189), .B2(G134), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n204), .A3(new_n191), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n200), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n205), .B2(G131), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT70), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(new_n213), .A3(new_n200), .A4(new_n207), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G128), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n220), .B(G146), .C1(new_n215), .C2(new_n216), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n219), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n210), .A2(new_n214), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n232), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n192), .B1(new_n203), .B2(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n203), .A2(KEYINPUT66), .A3(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n199), .A3(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n191), .B1(new_n240), .B2(new_n192), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n200), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n225), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT64), .B1(new_n218), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n225), .A2(new_n248), .A3(new_n249), .A4(new_n244), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n236), .B1(new_n243), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n229), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n254), .A2(G210), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT26), .B(G101), .Z(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT72), .B1(new_n253), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n262), .B(new_n259), .C1(new_n229), .C2(new_n252), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n236), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n237), .A2(new_n199), .A3(new_n238), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n194), .B1(new_n266), .B2(new_n197), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n239), .A2(new_n241), .A3(G131), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n251), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n229), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT30), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n212), .A2(new_n228), .A3(new_n200), .A4(new_n207), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n265), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n188), .B1(new_n264), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n269), .A2(new_n265), .ZN(new_n277));
  INV_X1    g091(.A(new_n228), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n212), .A2(new_n200), .A3(new_n207), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(KEYINPUT70), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n214), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n262), .B1(new_n281), .B2(new_n259), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n253), .A2(KEYINPUT72), .A3(new_n260), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n272), .B1(new_n229), .B2(new_n269), .ZN(new_n285));
  INV_X1    g099(.A(new_n274), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n236), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(KEYINPUT31), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n253), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n269), .A2(new_n273), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n229), .A2(new_n252), .B1(new_n236), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n292), .B2(new_n289), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n276), .A2(new_n288), .B1(new_n293), .B2(new_n259), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  INV_X1    g112(.A(G472), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n290), .B(new_n260), .C1(new_n292), .C2(new_n289), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n280), .A2(new_n214), .B1(new_n243), .B2(new_n251), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n274), .B1(new_n302), .B2(new_n272), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n281), .B1(new_n303), .B2(new_n236), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n300), .B(new_n301), .C1(new_n304), .C2(new_n260), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT74), .B(G902), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n281), .A2(KEYINPUT28), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n253), .B1(new_n302), .B2(new_n265), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(KEYINPUT28), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n259), .A2(new_n300), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n299), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n276), .A2(new_n288), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n293), .A2(new_n259), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n296), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n316), .B2(KEYINPUT32), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n284), .A2(KEYINPUT31), .A3(new_n287), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT31), .B1(new_n284), .B2(new_n287), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n295), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n187), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n298), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n298), .A2(new_n317), .A3(new_n323), .A4(KEYINPUT75), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT98), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT9), .B(G234), .Z(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT81), .ZN(new_n331));
  INV_X1    g145(.A(G902), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G221), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT82), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n220), .A2(KEYINPUT1), .A3(G146), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n219), .A2(new_n227), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  INV_X1    g152(.A(G104), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(G107), .ZN(new_n340));
  INV_X1    g154(.A(G107), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT3), .A3(G104), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G101), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT83), .B1(new_n341), .B2(G104), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n339), .A3(G107), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n339), .A2(G107), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n341), .A2(G104), .ZN(new_n350));
  OAI21_X1  g164(.A(G101), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n337), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n348), .A2(new_n351), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n228), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n243), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT12), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G101), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n348), .A2(KEYINPUT4), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n345), .A2(new_n347), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n344), .B1(new_n363), .B2(new_n343), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n251), .B(new_n361), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n353), .A2(KEYINPUT10), .A3(new_n228), .ZN(new_n366));
  INV_X1    g180(.A(new_n243), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n358), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G140), .ZN(new_n369));
  INV_X1    g183(.A(G953), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G227), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n369), .B(new_n371), .Z(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT12), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n354), .A2(new_n374), .A3(new_n243), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n356), .A2(new_n368), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n358), .A2(new_n365), .A3(new_n366), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n243), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n373), .B1(new_n378), .B2(new_n368), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n379), .B2(KEYINPUT84), .ZN(new_n380));
  INV_X1    g194(.A(new_n375), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n374), .B1(new_n354), .B2(new_n243), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n368), .A4(new_n373), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G469), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n306), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n307), .B1(new_n380), .B2(new_n385), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT85), .A3(new_n387), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n356), .A2(new_n368), .A3(new_n372), .A4(new_n375), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n378), .A2(new_n368), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n394), .B1(new_n395), .B2(new_n372), .ZN(new_n396));
  OAI21_X1  g210(.A(G469), .B1(new_n396), .B2(G902), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n335), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G214), .B1(G237), .B2(G902), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n236), .B(new_n361), .C1(new_n362), .C2(new_n364), .ZN(new_n400));
  INV_X1    g214(.A(G119), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G116), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n403));
  INV_X1    g217(.A(G113), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G116), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G119), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n407), .A3(KEYINPUT5), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(new_n233), .A3(new_n348), .A4(new_n351), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n400), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT6), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n400), .A2(new_n410), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G125), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n219), .A2(new_n421), .A3(new_n227), .A4(new_n221), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n251), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n370), .A2(G224), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT87), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n408), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n232), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n405), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(new_n233), .A3(new_n348), .A4(new_n351), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT89), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n353), .A2(new_n434), .A3(new_n233), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n409), .A2(new_n233), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n348), .A2(new_n351), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n411), .B(KEYINPUT8), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n423), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n422), .B(new_n445), .C1(new_n251), .C2(new_n421), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n442), .A2(KEYINPUT90), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n432), .A2(KEYINPUT89), .B1(new_n437), .B2(new_n436), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n440), .B1(new_n449), .B2(new_n435), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n446), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n452), .A3(new_n412), .ZN(new_n453));
  OAI21_X1  g267(.A(G210), .B1(G237), .B2(G902), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n427), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n427), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n399), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G140), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G125), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n421), .A2(G140), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n458), .A2(KEYINPUT77), .A3(G125), .ZN(new_n464));
  XNOR2_X1  g278(.A(G125), .B(G140), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT77), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n463), .B1(new_n467), .B2(new_n462), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n254), .A2(G143), .A3(G214), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(G143), .B1(new_n254), .B2(G214), .ZN(new_n471));
  OAI21_X1  g285(.A(G131), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G237), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n370), .A3(G214), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n220), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n194), .A3(new_n469), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n468), .A2(new_n222), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT16), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT78), .B1(new_n467), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n421), .A2(G140), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n478), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n459), .A2(new_n460), .A3(new_n466), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(KEYINPUT77), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT78), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT16), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n479), .A2(G146), .A3(new_n481), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(KEYINPUT18), .A2(G131), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n470), .B2(new_n471), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT91), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n475), .A2(new_n469), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n490), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n493), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n482), .A2(new_n483), .A3(G146), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n465), .A2(new_n222), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n497), .A2(new_n489), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n488), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n339), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n477), .A2(new_n487), .B1(new_n496), .B2(new_n500), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT92), .B1(new_n508), .B2(new_n505), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n486), .A2(new_n481), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(new_n485), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n222), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n472), .A2(new_n514), .A3(new_n476), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n493), .A2(KEYINPUT17), .A3(G131), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n517), .A3(new_n487), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n505), .A3(new_n501), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n507), .A2(new_n509), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT20), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n518), .A2(new_n505), .A3(new_n501), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n505), .B1(new_n518), .B2(new_n501), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n332), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT93), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT93), .B(new_n332), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(G475), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n220), .A2(G128), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n226), .A2(G143), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(G134), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n538), .A3(G134), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n534), .A2(new_n535), .A3(new_n538), .A4(G134), .ZN(new_n541));
  INV_X1    g355(.A(G122), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT94), .B1(new_n542), .B2(G116), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n406), .A3(G122), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n406), .A2(G122), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n341), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n548), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(G107), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n540), .B(new_n541), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n546), .A2(KEYINPUT14), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT14), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n543), .B2(new_n545), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n547), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n553), .B1(new_n556), .B2(KEYINPUT95), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n555), .B2(new_n547), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n341), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n537), .B1(G107), .B2(new_n550), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n552), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n331), .A2(G217), .A3(new_n370), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n563), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n552), .B(new_n565), .C1(new_n560), .C2(new_n561), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n307), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n567), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G952), .ZN(new_n574));
  AOI211_X1 g388(.A(G953), .B(new_n574), .C1(G234), .C2(G237), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI211_X1 g390(.A(new_n370), .B(new_n306), .C1(G234), .C2(G237), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT21), .B(G898), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT97), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n526), .A2(new_n533), .A3(new_n573), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n457), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n329), .B1(new_n398), .B2(new_n583), .ZN(new_n584));
  AND4_X1   g398(.A1(KEYINPUT85), .A2(new_n386), .A3(new_n387), .A4(new_n306), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT85), .B1(new_n391), .B2(new_n387), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n397), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n335), .ZN(new_n588));
  AND4_X1   g402(.A1(new_n329), .A2(new_n583), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G217), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n306), .B2(G234), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n513), .A2(new_n487), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n226), .A2(G119), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n401), .A2(G128), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT24), .B(G110), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT76), .B1(new_n226), .B2(G119), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT23), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n603), .B2(G110), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G110), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n601), .A2(new_n606), .A3(new_n595), .A4(new_n602), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n596), .A2(new_n597), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n607), .A2(new_n608), .B1(new_n222), .B2(new_n465), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n487), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n370), .A2(G221), .A3(G234), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT79), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT22), .B(G137), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n614), .ZN(new_n616));
  INV_X1    g430(.A(new_n604), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n513), .B2(new_n487), .ZN(new_n618));
  INV_X1    g432(.A(new_n610), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT25), .B1(new_n621), .B2(new_n306), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT25), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n623), .B(new_n307), .C1(new_n615), .C2(new_n620), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n592), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT80), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT80), .B(new_n592), .C1(new_n622), .C2(new_n624), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n592), .A2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n328), .A2(new_n590), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  OAI21_X1  g448(.A(G472), .B1(new_n294), .B2(new_n307), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n635), .A2(KEYINPUT99), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n316), .B1(new_n635), .B2(KEYINPUT99), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n398), .A2(new_n632), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT100), .ZN(new_n641));
  INV_X1    g455(.A(new_n457), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n642), .A2(new_n581), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n564), .A2(new_n566), .ZN(new_n644));
  OAI211_X1 g458(.A(KEYINPUT103), .B(new_n568), .C1(new_n644), .C2(new_n307), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n567), .B2(G478), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n644), .B2(KEYINPUT33), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT33), .B1(new_n564), .B2(new_n566), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT101), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n566), .A2(KEYINPUT102), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n566), .A2(KEYINPUT102), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(KEYINPUT33), .A3(new_n564), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n650), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n307), .A2(new_n568), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n648), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n526), .A2(new_n533), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n643), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n641), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NOR2_X1   g482(.A1(new_n661), .A2(new_n573), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n641), .A2(new_n643), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND2_X1  g486(.A1(new_n605), .A2(new_n610), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n614), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n629), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n627), .A2(new_n628), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n638), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n590), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  NOR2_X1   g496(.A1(new_n678), .A2(new_n457), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n575), .B(KEYINPUT104), .Z(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n578), .B2(G900), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n661), .A2(new_n573), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n683), .A2(new_n687), .A3(new_n398), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n328), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  INV_X1    g504(.A(new_n456), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n427), .A2(new_n453), .A3(new_n454), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT38), .Z(new_n694));
  INV_X1    g508(.A(new_n399), .ZN(new_n695));
  INV_X1    g509(.A(new_n573), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n661), .A2(new_n696), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n694), .A2(new_n695), .A3(new_n677), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n685), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n398), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n322), .B1(new_n321), .B2(new_n187), .ZN(new_n704));
  AOI211_X1 g518(.A(KEYINPUT73), .B(KEYINPUT32), .C1(new_n320), .C2(new_n295), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n284), .A2(new_n287), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n309), .A2(new_n259), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n299), .B1(new_n709), .B2(new_n332), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n316), .B2(KEYINPUT32), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT105), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n703), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n220), .ZN(G45));
  NOR3_X1   g529(.A1(new_n660), .A2(new_n662), .A3(new_n686), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n683), .A2(new_n398), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n328), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  NOR2_X1   g533(.A1(new_n391), .A2(new_n387), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n393), .A2(new_n334), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n664), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n328), .A2(new_n632), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND2_X1  g540(.A1(new_n643), .A2(new_n669), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n722), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT75), .B1(new_n706), .B2(new_n317), .ZN(new_n729));
  INV_X1    g543(.A(new_n327), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n632), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  NOR4_X1   g546(.A1(new_n722), .A2(new_n678), .A3(new_n582), .A4(new_n457), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n328), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n697), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n661), .A2(KEYINPUT106), .A3(new_n696), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n334), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n740), .B(new_n720), .C1(new_n390), .C2(new_n392), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n643), .A3(new_n741), .ZN(new_n742));
  OAI22_X1  g556(.A1(new_n318), .A2(new_n319), .B1(new_n260), .B2(new_n310), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n295), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n632), .A2(new_n635), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT107), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n642), .A2(new_n581), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n722), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n635), .A2(new_n744), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n631), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n739), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NAND3_X1  g568(.A1(new_n716), .A2(new_n741), .A3(new_n642), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n749), .B2(new_n678), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n677), .A2(new_n635), .A3(KEYINPUT108), .A4(new_n744), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n421), .ZN(G27));
  NOR2_X1   g574(.A1(new_n693), .A2(new_n695), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n397), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n396), .A2(KEYINPUT109), .A3(G469), .A4(new_n332), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n393), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n716), .A2(new_n334), .A3(new_n761), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n631), .B1(new_n317), .B2(new_n297), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(KEYINPUT42), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n631), .B1(new_n326), .B2(new_n327), .ZN(new_n772));
  INV_X1    g586(.A(new_n766), .ZN(new_n773));
  INV_X1    g587(.A(new_n761), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n740), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n716), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n771), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n194), .ZN(G33));
  NAND4_X1  g593(.A1(new_n328), .A2(new_n632), .A3(new_n687), .A4(new_n775), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n660), .A2(new_n661), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT43), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n638), .A3(new_n677), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n782), .B1(new_n786), .B2(KEYINPUT44), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(KEYINPUT44), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n387), .B1(new_n396), .B2(KEYINPUT45), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(KEYINPUT45), .B2(new_n396), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(KEYINPUT46), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n393), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n334), .A3(new_n699), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n774), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n787), .A2(new_n789), .A3(new_n790), .A4(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT112), .B(G137), .Z(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(G39));
  XNOR2_X1  g618(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n799), .A2(new_n334), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n805), .B1(new_n799), .B2(new_n334), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n716), .A2(new_n761), .A3(new_n631), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n328), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND4_X1  g624(.A1(new_n783), .A2(new_n632), .A3(new_n588), .A4(new_n399), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n393), .A2(new_n721), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(KEYINPUT49), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT114), .ZN(new_n814));
  INV_X1    g628(.A(new_n713), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n694), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n684), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n784), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(new_n750), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n695), .A2(new_n820), .A3(new_n694), .A4(new_n741), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n757), .A2(new_n758), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n722), .A2(new_n774), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n821), .A2(new_n822), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n815), .A2(new_n632), .A3(new_n575), .A4(new_n825), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n662), .A3(new_n660), .ZN(new_n830));
  OAI22_X1  g644(.A1(new_n806), .A2(new_n807), .B1(new_n588), .B2(new_n812), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n761), .A3(new_n820), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n823), .A2(new_n827), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n826), .A2(new_n769), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(KEYINPUT120), .A3(KEYINPUT48), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n741), .A2(new_n642), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n574), .B(G953), .C1(new_n820), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n839), .B(new_n844), .C1(new_n663), .C2(new_n829), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n835), .A2(new_n836), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  INV_X1    g661(.A(new_n759), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n773), .A2(new_n740), .A3(new_n677), .A4(new_n686), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n457), .B1(new_n737), .B2(new_n738), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n712), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n689), .A2(new_n718), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n759), .B1(new_n328), .B2(new_n688), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .A3(new_n718), .A4(new_n851), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(KEYINPUT117), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n724), .A2(new_n731), .A3(new_n734), .A4(new_n753), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n661), .A2(new_n696), .A3(new_n686), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n398), .A2(new_n863), .A3(new_n677), .A4(new_n761), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n328), .A2(new_n864), .B1(new_n824), .B2(new_n768), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n780), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n776), .A2(new_n777), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n770), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n640), .A2(new_n665), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n633), .A2(KEYINPUT115), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n727), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n640), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n680), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n633), .A2(new_n870), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n867), .A2(new_n869), .A3(new_n871), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT116), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n877), .A2(new_n871), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n778), .A2(new_n862), .A3(new_n866), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n861), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n854), .B2(new_n856), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n878), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n854), .A2(new_n887), .A3(new_n856), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n847), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n880), .A3(new_n881), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n885), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n880), .A4(new_n881), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n847), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT119), .B1(new_n892), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n894), .A2(new_n885), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n885), .B2(new_n884), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n900), .B(new_n897), .C1(new_n902), .C2(new_n847), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n846), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n817), .B1(new_n904), .B2(new_n905), .ZN(G75));
  AOI21_X1  g720(.A(KEYINPUT53), .B1(new_n889), .B2(new_n890), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n854), .A2(KEYINPUT117), .A3(new_n856), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT117), .B1(new_n854), .B2(new_n856), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT53), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n306), .ZN(new_n914));
  INV_X1    g728(.A(new_n454), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n420), .B(new_n426), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT55), .Z(new_n918));
  AND2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n370), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n916), .B2(new_n918), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n922), .ZN(G51));
  NOR3_X1   g737(.A1(new_n913), .A2(new_n306), .A3(new_n792), .ZN(new_n924));
  INV_X1    g738(.A(new_n386), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT54), .B1(new_n907), .B2(new_n912), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n897), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n793), .B(KEYINPUT57), .Z(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(KEYINPUT121), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n931));
  INV_X1    g745(.A(new_n928), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n926), .B2(new_n897), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n933), .B2(new_n925), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n920), .B1(new_n930), .B2(new_n934), .ZN(G54));
  NAND2_X1  g749(.A1(new_n895), .A2(new_n896), .ZN(new_n936));
  AND2_X1   g750(.A1(KEYINPUT58), .A2(G475), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n307), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n520), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n921), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT122), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n914), .A2(new_n520), .A3(new_n937), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n944), .A2(new_n945), .A3(new_n921), .A4(new_n940), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(G60));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT59), .Z(new_n949));
  NOR2_X1   g763(.A1(new_n656), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n927), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n921), .ZN(new_n952));
  INV_X1    g766(.A(new_n949), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n899), .A2(new_n903), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n954), .B2(new_n656), .ZN(G63));
  XNOR2_X1  g769(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n591), .A2(new_n332), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n936), .A2(new_n675), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n936), .A2(new_n958), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n621), .B(KEYINPUT124), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n921), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G66));
  AOI21_X1  g778(.A(new_n370), .B1(new_n580), .B2(G224), .ZN(new_n965));
  INV_X1    g779(.A(new_n862), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n880), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n967), .B2(new_n370), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n418), .B(new_n419), .C1(G898), .C2(new_n370), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT125), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(G69));
  NAND2_X1  g785(.A1(new_n769), .A2(new_n850), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT126), .B1(new_n800), .B2(new_n972), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n800), .A2(KEYINPUT126), .A3(new_n972), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n809), .A2(new_n780), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n855), .A2(new_n718), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n802), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n975), .A2(new_n977), .A3(new_n778), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n370), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n303), .B(new_n468), .ZN(new_n980));
  NAND2_X1  g794(.A1(G900), .A2(G953), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n761), .B1(new_n663), .B2(new_n669), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n700), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n772), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n809), .A2(new_n802), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n714), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n976), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(KEYINPUT62), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  AOI21_X1  g804(.A(G953), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n982), .B1(new_n991), .B2(new_n980), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n370), .B1(G227), .B2(G900), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n967), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n978), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n304), .A2(new_n259), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n921), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n304), .A2(new_n259), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n989), .A2(new_n998), .A3(new_n990), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n996), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n707), .B1(new_n260), .B2(new_n304), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n996), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n902), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT127), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1006), .B(new_n1011), .C1(new_n902), .C2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(G57));
endmodule


