//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(KEYINPUT89), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n217), .A2(new_n218), .B1(new_n214), .B2(new_n215), .ZN(new_n219));
  OR3_X1    g018(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT17), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT17), .B1(new_n219), .B2(new_n220), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n207), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n219), .A2(new_n206), .A3(new_n220), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n224), .A2(KEYINPUT18), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n218), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n214), .A2(new_n215), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n220), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n225), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n226), .B(KEYINPUT13), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n206), .B1(new_n237), .B2(new_n221), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n225), .A2(new_n226), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n227), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G141gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G197gat), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT11), .B(G169gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n227), .A2(new_n240), .A3(new_n246), .A4(new_n234), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(KEYINPUT90), .A3(new_n247), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n258), .A3(G113gat), .ZN(new_n259));
  INV_X1    g058(.A(G113gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G120gat), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT66), .B1(new_n259), .B2(new_n261), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264));
  AND2_X1   g063(.A1(G127gat), .A2(G134gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G127gat), .A2(G134gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n262), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(new_n266), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT64), .B(KEYINPUT28), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT27), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n274), .A3(new_n280), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  AND2_X1   g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(KEYINPUT26), .B2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n282), .A2(new_n284), .A3(new_n286), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n287), .A2(new_n291), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  INV_X1    g092(.A(G169gat), .ZN(new_n294));
  INV_X1    g093(.A(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G183gat), .B(G190gat), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n292), .B(new_n298), .C1(new_n291), .C2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(KEYINPUT24), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n276), .A2(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n280), .A2(G183gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n308), .B2(KEYINPUT24), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT25), .B1(new_n309), .B2(new_n298), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n290), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n273), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G227gat), .A2(G233gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT34), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n314), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G15gat), .B(G43gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(G71gat), .B(G99gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n259), .A2(new_n261), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n261), .ZN(new_n325));
  INV_X1    g124(.A(new_n267), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n271), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n311), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(G227gat), .A3(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT33), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n321), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(KEYINPUT32), .C1(new_n331), .C2(new_n321), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n318), .B1(new_n334), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n254), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n335), .ZN(new_n340));
  INV_X1    g139(.A(new_n318), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT87), .A3(new_n336), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n346));
  INV_X1    g145(.A(G197gat), .ZN(new_n347));
  INV_X1    g146(.A(G204gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G197gat), .A2(G204gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n345), .B1(new_n351), .B2(KEYINPUT69), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(KEYINPUT69), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n345), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AND2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G141gat), .B(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT2), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(G155gat), .B2(G162gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G141gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G148gat), .ZN(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G155gat), .B(G162gat), .ZN(new_n369));
  INV_X1    g168(.A(G155gat), .ZN(new_n370));
  INV_X1    g169(.A(G162gat), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT2), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n363), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n355), .B1(new_n356), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G228gat), .ZN(new_n377));
  INV_X1    g176(.A(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n373), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n354), .A2(KEYINPUT29), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n355), .A2(new_n385), .A3(new_n356), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT81), .B1(new_n354), .B2(KEYINPUT29), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n374), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n376), .B1(new_n388), .B2(new_n381), .ZN(new_n389));
  INV_X1    g188(.A(new_n379), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n384), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT31), .B(G50gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n392), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n384), .B(new_n394), .C1(new_n389), .C2(new_n390), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G22gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(new_n398), .A3(new_n395), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT35), .ZN(new_n403));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n328), .A2(new_n375), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n271), .A2(new_n363), .A3(new_n373), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n327), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n415), .B2(KEYINPUT4), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417));
  AOI211_X1 g216(.A(KEYINPUT76), .B(new_n417), .C1(new_n327), .C2(new_n414), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n271), .A2(new_n363), .A3(new_n373), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n268), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n327), .B2(new_n414), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n417), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n412), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT77), .B1(new_n268), .B2(new_n420), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n381), .B1(new_n268), .B2(new_n272), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n327), .A2(new_n414), .A3(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n411), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT78), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n425), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT4), .B1(new_n421), .B2(new_n423), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n415), .A2(new_n417), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n440));
  INV_X1    g239(.A(new_n412), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n408), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n419), .A2(new_n424), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n441), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT78), .B1(new_n431), .B2(KEYINPUT5), .ZN(new_n448));
  AOI211_X1 g247(.A(new_n433), .B(new_n440), .C1(new_n429), .C2(new_n430), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(new_n407), .A3(new_n442), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n407), .B1(new_n450), .B2(new_n442), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n344), .A2(new_n402), .A3(new_n403), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n311), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT70), .B(new_n290), .C1(new_n302), .C2(new_n310), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT71), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n459), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n300), .A2(new_n301), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n309), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT70), .B1(new_n467), .B2(new_n290), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n356), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT71), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n461), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n311), .A2(new_n462), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n463), .A2(new_n471), .A3(new_n355), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n462), .A3(new_n459), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n311), .A2(new_n356), .A3(new_n461), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n354), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G8gat), .B(G36gat), .Z(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT72), .ZN(new_n479));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT73), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(KEYINPUT30), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n473), .A2(new_n476), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n476), .A3(new_n481), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n488), .B1(new_n487), .B2(new_n491), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n456), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT79), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n445), .B(new_n451), .C1(new_n453), .C2(new_n498), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT79), .B(new_n407), .C1(new_n450), .C2(new_n442), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n454), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n473), .A2(new_n476), .A3(new_n485), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n482), .B1(new_n473), .B2(new_n476), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT74), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT74), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n505), .A3(new_n486), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n504), .A2(new_n506), .B1(new_n489), .B2(new_n490), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT80), .B1(new_n501), .B2(new_n507), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n318), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n336), .B(new_n511), .C1(new_n342), .C2(new_n510), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n402), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n508), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n497), .B1(new_n514), .B2(new_n403), .ZN(new_n515));
  INV_X1    g314(.A(new_n402), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n508), .B2(new_n509), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT36), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(KEYINPUT36), .B2(new_n512), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT37), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n473), .A2(new_n520), .A3(new_n476), .ZN(new_n521));
  INV_X1    g320(.A(new_n481), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n473), .B2(new_n476), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT38), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n477), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT38), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n482), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n463), .A2(new_n471), .A3(new_n354), .A4(new_n472), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n474), .A2(new_n355), .A3(new_n475), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n530), .A2(KEYINPUT37), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n526), .A2(new_n481), .B1(new_n532), .B2(new_n521), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n525), .A2(new_n452), .A3(new_n454), .A4(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n534), .A2(new_n402), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT40), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n429), .A2(new_n430), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n537), .A2(KEYINPUT39), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n437), .A2(new_n410), .A3(new_n438), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n430), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n430), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT84), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n543), .A2(new_n544), .A3(new_n407), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n543), .B2(new_n407), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n541), .B(KEYINPUT86), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n444), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n407), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT84), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n544), .A3(new_n407), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT86), .B1(new_n552), .B2(new_n541), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n540), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n545), .B2(new_n546), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT85), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n552), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n559), .A3(new_n536), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n554), .B(new_n560), .C1(new_n494), .C2(new_n492), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n519), .B1(new_n535), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n517), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n253), .B1(new_n515), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n454), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n450), .A2(new_n442), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n498), .B1(new_n566), .B2(new_n408), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n451), .A2(new_n445), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n500), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n565), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT96), .ZN(new_n573));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G99gat), .B(G106gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n577), .B1(new_n587), .B2(new_n230), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n587), .B1(new_n222), .B2(new_n223), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n576), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n591), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n592), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n594), .A3(new_n575), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(G57gat), .A2(G64gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(G57gat), .A2(G64gat), .ZN(new_n603));
  AND2_X1   g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(KEYINPUT9), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n606), .B2(new_n604), .ZN(new_n607));
  XNOR2_X1  g406(.A(G71gat), .B(G78gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n207), .B1(new_n610), .B2(new_n609), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT93), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT92), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n615), .B(new_n622), .Z(new_n623));
  NOR2_X1   g422(.A1(new_n601), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n587), .A2(new_n609), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n585), .A2(new_n586), .ZN(new_n627));
  INV_X1    g426(.A(new_n586), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n628), .B1(new_n582), .B2(new_n584), .ZN(new_n629));
  OR3_X1    g428(.A1(new_n627), .A2(new_n609), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n587), .A2(KEYINPUT97), .A3(new_n609), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT10), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n625), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n633), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n625), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n639), .B(new_n642), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n624), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n564), .A2(new_n571), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g446(.A1(new_n564), .A2(new_n496), .A3(new_n645), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n648), .A2(G8gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT16), .B(G8gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT42), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(KEYINPUT42), .B2(new_n651), .ZN(G1325gat));
  NAND2_X1  g452(.A1(new_n564), .A2(new_n645), .ZN(new_n654));
  INV_X1    g453(.A(new_n519), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n344), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n654), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n654), .A2(new_n402), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(new_n601), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n515), .B2(new_n563), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n639), .B(new_n642), .ZN(new_n665));
  INV_X1    g464(.A(new_n623), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n665), .A2(new_n253), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(G29gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n571), .A2(new_n669), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n668), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  INV_X1    g473(.A(new_n667), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n456), .A2(new_n496), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT80), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n504), .A2(new_n506), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n491), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n571), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n507), .ZN(new_n681));
  INV_X1    g480(.A(new_n513), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n676), .B1(new_n683), .B2(KEYINPUT35), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n535), .A2(new_n561), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n655), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n402), .B1(new_n680), .B2(new_n681), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT100), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n517), .A2(new_n562), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n684), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n663), .A2(KEYINPUT44), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT101), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n517), .A2(new_n562), .A3(new_n689), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n689), .B1(new_n517), .B2(new_n562), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n515), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n692), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT99), .B1(new_n664), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n601), .B1(new_n703), .B2(new_n684), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n675), .B1(new_n700), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(new_n571), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n674), .B1(new_n669), .B2(new_n709), .ZN(G1328gat));
  INV_X1    g509(.A(G36gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n496), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT46), .B1(new_n668), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n668), .A2(new_n712), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n717), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n715), .A2(new_n716), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n708), .A2(new_n496), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n711), .B2(new_n724), .ZN(G1329gat));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n708), .B2(new_n519), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n664), .A2(new_n727), .A3(new_n344), .A4(new_n667), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n726), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n655), .B(new_n675), .C1(new_n700), .C2(new_n707), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT47), .B(new_n729), .C1(new_n732), .C2(new_n727), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1330gat));
  XOR2_X1   g533(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n735));
  INV_X1    g534(.A(G50gat), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n708), .B2(new_n516), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n664), .A2(new_n736), .A3(new_n516), .A4(new_n667), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI211_X1 g539(.A(new_n402), .B(new_n675), .C1(new_n700), .C2(new_n707), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT48), .B(new_n738), .C1(new_n741), .C2(new_n736), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1331gat));
  NAND3_X1  g542(.A1(new_n624), .A2(new_n253), .A3(new_n665), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n691), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n571), .B(KEYINPUT105), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  INV_X1    g547(.A(new_n496), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n691), .A2(new_n749), .A3(new_n744), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  NAND2_X1  g553(.A1(new_n745), .A2(new_n519), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n657), .A2(G71gat), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n755), .A2(G71gat), .B1(new_n745), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n745), .A2(new_n516), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n251), .A2(new_n252), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n666), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n663), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n691), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n697), .A2(KEYINPUT51), .A3(new_n765), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n769), .A2(new_n579), .A3(new_n571), .A4(new_n665), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n764), .A2(new_n643), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n700), .B2(new_n707), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n571), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n774), .B2(new_n579), .ZN(G1336gat));
  NAND3_X1  g574(.A1(new_n767), .A2(KEYINPUT106), .A3(new_n768), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n777), .B(new_n761), .C1(new_n691), .C2(new_n766), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n749), .A2(G92gat), .A3(new_n643), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n691), .A2(KEYINPUT101), .A3(new_n693), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n698), .B1(new_n697), .B2(new_n692), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n664), .A2(KEYINPUT99), .A3(new_n701), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n705), .B1(new_n704), .B2(KEYINPUT44), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n781), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n496), .A3(new_n771), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n780), .B1(G92gat), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n580), .B1(new_n773), .B2(new_n496), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n769), .A2(new_n779), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT107), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n769), .A2(new_n792), .A3(new_n779), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n794), .ZN(G1337gat));
  XNOR2_X1  g594(.A(KEYINPUT109), .B(G99gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n657), .A2(new_n643), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n769), .A2(new_n797), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n655), .B(new_n772), .C1(new_n700), .C2(new_n707), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n799), .B2(KEYINPUT108), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n773), .A2(KEYINPUT108), .A3(new_n519), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(G1338gat));
  NOR3_X1   g601(.A1(new_n643), .A2(new_n402), .A3(G106gat), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT111), .Z(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n769), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n402), .B(new_n772), .C1(new_n700), .C2(new_n707), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT110), .B(G106gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n776), .A2(new_n778), .A3(new_n804), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n773), .A2(new_n516), .ZN(new_n810));
  INV_X1    g609(.A(new_n807), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n624), .A2(new_n643), .A3(new_n253), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n624), .A2(new_n643), .A3(KEYINPUT112), .A4(new_n253), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n636), .B1(new_n638), .B2(new_n635), .ZN(new_n820));
  INV_X1    g619(.A(new_n625), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n637), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n824), .B(new_n625), .C1(new_n634), .C2(new_n636), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n642), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n226), .B1(new_n224), .B2(new_n225), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n232), .A2(new_n233), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n245), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n250), .B1(new_n829), .B2(KEYINPUT113), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n831));
  INV_X1    g630(.A(new_n225), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n238), .A2(new_n832), .ZN(new_n833));
  OAI22_X1  g632(.A1(new_n833), .A2(new_n226), .B1(new_n232), .B2(new_n233), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n831), .B1(new_n834), .B2(new_n245), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n601), .A2(new_n826), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n639), .A2(new_n642), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n825), .A2(new_n642), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n637), .A2(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n822), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n842), .B2(KEYINPUT55), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n665), .A2(new_n836), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n826), .A2(new_n252), .A3(new_n251), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n663), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n819), .B1(new_n848), .B2(new_n666), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n516), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n496), .A2(new_n657), .A3(new_n501), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n260), .A3(new_n253), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n746), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(new_n496), .A3(new_n513), .ZN(new_n856));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n762), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n854), .A2(new_n857), .ZN(G1340gat));
  NAND4_X1  g657(.A1(new_n856), .A2(new_n256), .A3(new_n258), .A4(new_n665), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n851), .A2(new_n665), .A3(new_n852), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n860), .A2(KEYINPUT114), .A3(G120gat), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT114), .B1(new_n860), .B2(G120gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n853), .B2(new_n623), .ZN(new_n864));
  INV_X1    g663(.A(G127gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n856), .A2(new_n865), .A3(new_n666), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n856), .A2(new_n868), .A3(new_n601), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT115), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n853), .B2(new_n663), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n871), .B(new_n872), .C1(KEYINPUT56), .C2(new_n869), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT121), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT122), .Z(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n749), .A2(new_n655), .A3(new_n571), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n849), .A2(new_n516), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT116), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n882), .B(KEYINPUT57), .C1(new_n849), .C2(new_n516), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n402), .A2(new_n880), .ZN(new_n885));
  INV_X1    g684(.A(new_n844), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n823), .A2(new_n642), .A3(new_n825), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT55), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n762), .A2(new_n889), .A3(new_n839), .A4(new_n826), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n601), .B1(new_n890), .B2(new_n845), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n847), .A2(new_n663), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT118), .B(new_n623), .C1(new_n893), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n819), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n891), .A2(new_n892), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n886), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT118), .B1(new_n900), .B2(new_n623), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n885), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n878), .B1(new_n884), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n364), .B1(new_n903), .B2(new_n762), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n855), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n849), .A2(KEYINPUT119), .A3(new_n746), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n519), .A2(new_n402), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT120), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n496), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n253), .A2(G141gat), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n912), .A2(new_n914), .B1(KEYINPUT121), .B2(new_n874), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n877), .B1(new_n904), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n915), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n253), .B(new_n878), .C1(new_n884), .C2(new_n902), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n917), .B(new_n876), .C1(new_n918), .C2(new_n364), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1344gat));
  OAI21_X1  g719(.A(KEYINPUT59), .B1(new_n912), .B2(new_n643), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n366), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n815), .B1(new_n848), .B2(new_n666), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n402), .B1(new_n923), .B2(KEYINPUT123), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT57), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n849), .A2(new_n885), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n878), .A2(new_n643), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT59), .B(G148gat), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n884), .A2(new_n902), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n930), .A2(KEYINPUT59), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n922), .B(new_n931), .C1(new_n932), .C2(new_n933), .ZN(G1345gat));
  AOI21_X1  g733(.A(new_n370), .B1(new_n903), .B2(new_n666), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n912), .A2(G155gat), .A3(new_n623), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT124), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n936), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n623), .B(new_n878), .C1(new_n884), .C2(new_n902), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n370), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n937), .A2(new_n941), .ZN(G1346gat));
  INV_X1    g741(.A(new_n912), .ZN(new_n943));
  AOI21_X1  g742(.A(G162gat), .B1(new_n943), .B2(new_n601), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n663), .A2(new_n371), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n903), .B2(new_n945), .ZN(G1347gat));
  NOR3_X1   g745(.A1(new_n850), .A2(new_n571), .A3(new_n749), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n682), .ZN(new_n948));
  AOI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n762), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n746), .A2(new_n749), .A3(new_n657), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n851), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n253), .A2(new_n294), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1348gat));
  INV_X1    g752(.A(new_n951), .ZN(new_n954));
  OAI21_X1  g753(.A(G176gat), .B1(new_n954), .B2(new_n643), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n948), .A2(new_n295), .A3(new_n665), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n958), .A2(KEYINPUT60), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n958), .A2(KEYINPUT60), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n948), .A2(new_n283), .A3(new_n666), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n851), .A2(new_n666), .A3(new_n950), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G183gat), .ZN(new_n963));
  AOI211_X1 g762(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  AND4_X1   g763(.A1(new_n958), .A2(new_n961), .A3(KEYINPUT60), .A4(new_n963), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n280), .A3(new_n601), .ZN(new_n967));
  OAI21_X1  g766(.A(G190gat), .B1(new_n954), .B2(new_n663), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NAND2_X1  g770(.A1(new_n947), .A2(new_n909), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n762), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n746), .A2(new_n749), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n655), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n928), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n253), .A2(new_n347), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NOR3_X1   g778(.A1(new_n972), .A2(G204gat), .A3(new_n643), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n928), .A2(new_n643), .A3(new_n976), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n348), .B2(new_n982), .ZN(G1353gat));
  OR3_X1    g782(.A1(new_n972), .A2(G211gat), .A3(new_n623), .ZN(new_n984));
  INV_X1    g783(.A(new_n976), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n666), .B(new_n985), .C1(new_n926), .C2(new_n927), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  NAND2_X1  g788(.A1(new_n601), .A2(G218gat), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT126), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n985), .B(new_n991), .C1(new_n926), .C2(new_n927), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n972), .A2(new_n663), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n992), .B1(G218gat), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


