//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(G116), .B(G119), .Z(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(new_n188), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n198), .A2(KEYINPUT65), .A3(G146), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT65), .B1(new_n198), .B2(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n201), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G134), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G137), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n214), .A2(G131), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n215), .A2(new_n217), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n207), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n197), .A3(new_n199), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n198), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n196), .B2(G143), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n198), .A2(KEYINPUT65), .A3(G146), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n225), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n227), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(G137), .B1(new_n209), .B2(new_n211), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n212), .B2(G134), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n208), .A3(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n221), .A2(new_n220), .A3(new_n222), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n234), .A2(new_n240), .A3(new_n241), .A4(KEYINPUT68), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n224), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n234), .A2(new_n240), .A3(new_n241), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n195), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  AND4_X1   g061(.A1(new_n195), .A2(new_n246), .A3(new_n242), .A4(new_n224), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n187), .B(KEYINPUT28), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n250));
  INV_X1    g064(.A(new_n246), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n224), .A2(new_n242), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n194), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n246), .A2(new_n195), .A3(new_n242), .A4(new_n224), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n224), .A2(new_n195), .A3(new_n244), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n249), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT26), .B(G101), .Z(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n260), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n259), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n246), .A2(KEYINPUT30), .A3(new_n242), .A4(new_n224), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n271));
  INV_X1    g085(.A(new_n244), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n200), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n200), .A2(new_n205), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n232), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G131), .B1(new_n214), .B2(new_n218), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n241), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n271), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n270), .A2(new_n194), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n254), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n266), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n266), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n195), .B1(new_n224), .B2(new_n244), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n250), .B2(new_n256), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n243), .A2(KEYINPUT28), .A3(new_n195), .A4(new_n246), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n267), .B1(new_n290), .B2(new_n266), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n269), .A2(KEYINPUT73), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n293), .B(G902), .C1(new_n259), .C2(new_n268), .ZN(new_n294));
  OAI21_X1  g108(.A(G472), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n270), .A2(new_n194), .A3(new_n279), .ZN(new_n299));
  INV_X1    g113(.A(new_n266), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n254), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n300), .A2(new_n254), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT31), .A3(new_n280), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n300), .B1(new_n288), .B2(new_n289), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n297), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI211_X1 g122(.A(KEYINPUT70), .B(new_n306), .C1(new_n302), .C2(new_n304), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n296), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n296), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(new_n311), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n308), .B2(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n299), .A2(new_n298), .A3(new_n301), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT31), .B1(new_n303), .B2(new_n280), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n307), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n305), .A2(new_n297), .A3(new_n307), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n314), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n295), .A2(new_n312), .A3(new_n316), .A4(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G210), .B1(G237), .B2(G902), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT86), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n192), .A2(new_n188), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G116), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT82), .A4(G116), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G113), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n329), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n340));
  XNOR2_X1  g154(.A(G104), .B(G107), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G104), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT3), .B1(new_n344), .B2(G107), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  INV_X1    g160(.A(G107), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G104), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(G107), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n345), .A2(new_n348), .A3(new_n342), .A4(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n344), .A2(G107), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n347), .A2(G104), .ZN(new_n352));
  OAI211_X1 g166(.A(KEYINPUT80), .B(G101), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n343), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n339), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n356), .A2(G113), .A3(new_n334), .A4(new_n335), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n191), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n343), .A2(new_n350), .A3(new_n353), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G122), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT8), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT1), .ZN(new_n366));
  OAI21_X1  g180(.A(G128), .B1(new_n228), .B2(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n204), .A2(new_n367), .B1(new_n273), .B2(new_n226), .ZN(new_n368));
  INV_X1    g182(.A(G125), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n276), .A2(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n262), .A2(G224), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n370), .A2(KEYINPUT7), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n371), .ZN(new_n374));
  OR2_X1    g188(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n364), .A2(new_n365), .A3(new_n373), .A4(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n383), .A3(G101), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n194), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n355), .A2(new_n385), .A3(new_n362), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n361), .A2(new_n363), .B1(new_n374), .B2(new_n377), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n365), .B1(new_n388), .B2(new_n373), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n328), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n374), .B(new_n372), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n355), .A2(new_n385), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n355), .A2(new_n385), .A3(KEYINPUT83), .ZN(new_n395));
  INV_X1    g209(.A(new_n362), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(KEYINPUT6), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n362), .B1(new_n392), .B2(new_n393), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n391), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n327), .B1(new_n390), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n391), .ZN(new_n404));
  INV_X1    g218(.A(new_n401), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n400), .A2(new_n395), .B1(KEYINPUT6), .B2(new_n386), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n327), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n364), .A2(new_n373), .A3(new_n378), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT85), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n386), .A3(new_n379), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n407), .A2(new_n328), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n403), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT87), .B(new_n327), .C1(new_n390), .C2(new_n402), .ZN(new_n415));
  INV_X1    g229(.A(G952), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n416), .A2(KEYINPUT96), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(KEYINPUT96), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n262), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(G234), .B2(G237), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT97), .Z(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(G898), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n422), .B(KEYINPUT98), .Z(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n328), .B(new_n262), .C1(G234), .C2(G237), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n414), .A2(new_n415), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G113), .B(G122), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(new_n344), .ZN(new_n436));
  INV_X1    g250(.A(G140), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G125), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n369), .A2(G140), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT77), .ZN(new_n440));
  OR3_X1    g254(.A1(new_n369), .A2(KEYINPUT77), .A3(G140), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(G146), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n438), .A2(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n196), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT89), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n261), .A2(new_n262), .A3(G214), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n198), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n261), .A2(new_n262), .A3(G143), .A4(G214), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(KEYINPUT18), .A2(G131), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT16), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT16), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n438), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G146), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n453), .A2(G131), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n451), .A2(new_n220), .A3(new_n452), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n443), .A2(KEYINPUT19), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n440), .A2(new_n441), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(KEYINPUT19), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n462), .B(new_n465), .C1(new_n468), .C2(G146), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n436), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n455), .B1(new_n448), .B2(new_n446), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n472), .A3(new_n464), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n458), .A2(new_n196), .A3(new_n460), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n196), .B1(new_n458), .B2(new_n460), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n472), .B(new_n220), .C1(new_n451), .C2(new_n452), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n478), .B2(KEYINPUT90), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n458), .A2(new_n196), .A3(new_n460), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n462), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n482), .B2(new_n477), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n471), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n470), .B1(new_n484), .B2(new_n436), .ZN(new_n485));
  NOR2_X1   g299(.A1(G475), .A2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT91), .B(new_n434), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n453), .A2(KEYINPUT17), .A3(G131), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n462), .A2(KEYINPUT90), .A3(new_n481), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n473), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n436), .B(new_n457), .C1(new_n490), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n436), .ZN(new_n495));
  INV_X1    g309(.A(new_n469), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n471), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n487), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n489), .B1(new_n498), .B2(new_n433), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n488), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G122), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G116), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n347), .B1(new_n504), .B2(KEYINPUT14), .ZN(new_n505));
  XNOR2_X1  g319(.A(G116), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n198), .A2(G128), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n225), .A2(KEYINPUT92), .A3(G143), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT92), .B1(new_n225), .B2(G143), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n209), .A2(new_n211), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT94), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n511), .B(new_n512), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n506), .B(new_n347), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n508), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n198), .A2(KEYINPUT13), .A3(G128), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n523), .B(new_n524), .C1(new_n509), .C2(new_n510), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n525), .A2(KEYINPUT93), .A3(G134), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT93), .B1(new_n525), .B2(G134), .ZN(new_n527));
  OAI221_X1 g341(.A(new_n521), .B1(new_n512), .B2(new_n511), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT9), .B(G234), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(G217), .A3(new_n262), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n532), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n520), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n536), .B(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n484), .A2(new_n436), .ZN(new_n543));
  INV_X1    g357(.A(new_n494), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n328), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G475), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n502), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G221), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n531), .B2(new_n328), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n227), .B1(new_n233), .B2(new_n273), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(new_n350), .A3(new_n353), .A4(new_n343), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n354), .B2(new_n234), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n219), .A2(new_n223), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT12), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G140), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n262), .A2(G227), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n354), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT10), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n552), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n382), .A2(new_n207), .A3(new_n384), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n564), .A3(new_n565), .A4(new_n554), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n553), .A2(new_n555), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n557), .A2(new_n561), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT81), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n555), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n566), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n569), .A2(new_n570), .B1(new_n573), .B2(new_n560), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n368), .A2(new_n359), .ZN(new_n575));
  AOI221_X4 g389(.A(KEYINPUT12), .B1(new_n241), .B2(new_n277), .C1(new_n575), .C2(new_n552), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n567), .B1(new_n553), .B2(new_n555), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(KEYINPUT81), .A3(new_n561), .A4(new_n566), .ZN(new_n579));
  AOI211_X1 g393(.A(G469), .B(G902), .C1(new_n574), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n572), .A2(new_n561), .A3(new_n566), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n578), .A2(new_n566), .ZN(new_n582));
  OAI211_X1 g396(.A(G469), .B(new_n581), .C1(new_n582), .C2(new_n561), .ZN(new_n583));
  NAND2_X1  g397(.A1(G469), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n550), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n432), .A2(new_n547), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT24), .B(G110), .Z(new_n588));
  INV_X1    g402(.A(KEYINPUT75), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n225), .A2(G119), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n331), .A2(G128), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n588), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT24), .B(G110), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT75), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT76), .B1(new_n331), .B2(G128), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT23), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT23), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n590), .A2(KEYINPUT76), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n599), .A3(new_n591), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n592), .A2(new_n595), .B1(new_n600), .B2(G110), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n475), .B2(new_n476), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT78), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n601), .B(new_n604), .C1(new_n475), .C2(new_n476), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n593), .A2(new_n594), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n600), .B2(G110), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n462), .A2(new_n608), .A3(new_n444), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT22), .B(G137), .ZN(new_n610));
  INV_X1    g424(.A(G234), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n548), .A2(new_n611), .A3(G953), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n610), .B(new_n612), .Z(new_n613));
  AND3_X1   g427(.A1(new_n606), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n606), .B2(new_n609), .ZN(new_n615));
  OAI21_X1  g429(.A(G217), .B1(new_n611), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n328), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT79), .ZN(new_n619));
  INV_X1    g433(.A(new_n605), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n604), .B1(new_n482), .B2(new_n601), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n609), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n613), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n606), .A2(new_n609), .A3(new_n613), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n328), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n616), .B1(new_n626), .B2(KEYINPUT25), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n614), .A2(new_n615), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT25), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n328), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n619), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n325), .A2(new_n587), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  NOR2_X1   g449(.A1(new_n632), .A2(new_n586), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n328), .B1(new_n308), .B2(new_n309), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n637), .A2(G472), .B1(new_n322), .B2(new_n296), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n537), .A2(new_n328), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n536), .B2(new_n537), .ZN(new_n641));
  INV_X1    g455(.A(new_n535), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n534), .B1(new_n520), .B2(new_n528), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT33), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n533), .A2(new_n645), .A3(new_n535), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(G478), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n502), .B2(new_n546), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n430), .B1(new_n403), .B2(new_n412), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n649), .A2(new_n427), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n639), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT99), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n488), .A2(new_n499), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n498), .A2(new_n433), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(new_n488), .B2(new_n499), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT101), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n488), .A2(new_n499), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT100), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n657), .A4(new_n658), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n542), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n546), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n666), .A2(new_n427), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n666), .A2(new_n672), .A3(new_n427), .A4(new_n669), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n671), .A2(new_n639), .A3(new_n650), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  INV_X1    g490(.A(new_n432), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n547), .A2(new_n586), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n623), .A2(KEYINPUT36), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n622), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n622), .A2(new_n679), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n680), .A2(new_n681), .A3(new_n617), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n627), .B2(new_n630), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n677), .A2(new_n638), .A3(new_n678), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT37), .B(G110), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AND2_X1   g502(.A1(new_n583), .A2(new_n584), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n569), .A2(new_n570), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n573), .A2(new_n560), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n579), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(G469), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n328), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n549), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n695), .A2(new_n650), .A3(new_n684), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n325), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(G900), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n425), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n421), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n668), .B(new_n700), .C1(new_n661), .C2(new_n665), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  NAND2_X1  g517(.A1(new_n414), .A2(new_n415), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT38), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n700), .B(KEYINPUT39), .Z(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n586), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n253), .A2(new_n254), .A3(new_n266), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n328), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n266), .B1(new_n280), .B2(new_n254), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n312), .A2(new_n316), .A3(new_n324), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n502), .A2(new_n546), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n429), .A3(new_n667), .A4(new_n683), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n710), .B2(KEYINPUT40), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n706), .A2(new_n711), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  INV_X1    g535(.A(new_n700), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n649), .A2(KEYINPUT104), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT104), .B1(new_n649), .B2(new_n722), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n697), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n693), .B1(new_n692), .B2(new_n328), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n580), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n730), .B2(new_n550), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n580), .A2(new_n729), .A3(KEYINPUT105), .A4(new_n549), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n325), .A2(new_n733), .A3(new_n633), .A4(new_n651), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  AND3_X1   g550(.A1(new_n325), .A2(new_n733), .A3(new_n633), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n671), .A2(new_n737), .A3(new_n650), .A4(new_n673), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NAND2_X1  g553(.A1(new_n692), .A2(new_n328), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G469), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n694), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT105), .B1(new_n742), .B2(new_n549), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n730), .A2(new_n728), .A3(new_n550), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n743), .A2(new_n650), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n547), .A2(new_n428), .A3(new_n683), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n325), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G119), .ZN(G21));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n249), .B(new_n266), .C1(new_n255), .C2(new_n258), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n313), .B1(new_n750), .B2(new_n305), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n753));
  INV_X1    g567(.A(G472), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n632), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n428), .B(new_n542), .C1(new_n502), .C2(new_n546), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n743), .A3(new_n650), .A4(new_n744), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n749), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n745), .A2(KEYINPUT106), .A3(new_n756), .A4(new_n758), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n684), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n723), .A2(new_n724), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n766), .B2(new_n745), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n751), .B(new_n683), .C1(new_n637), .C2(G472), .ZN(new_n768));
  INV_X1    g582(.A(new_n648), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n717), .A2(new_n769), .A3(new_n722), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n649), .A2(KEYINPUT104), .A3(new_n722), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n768), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n743), .A2(new_n650), .A3(new_n744), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n774), .A2(KEYINPUT107), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  INV_X1    g593(.A(new_n725), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n704), .A2(new_n429), .A3(new_n695), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n325), .A2(new_n781), .A3(new_n633), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n430), .B1(new_n414), .B2(new_n415), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n695), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n779), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n312), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n310), .A2(KEYINPUT108), .A3(new_n311), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n295), .A3(new_n315), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n725), .A2(new_n786), .A3(new_n790), .A4(new_n633), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n783), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  NAND3_X1  g607(.A1(new_n666), .A2(new_n669), .A3(new_n722), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n782), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n208), .ZN(G36));
  INV_X1    g610(.A(new_n717), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n769), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT43), .Z(new_n799));
  NOR2_X1   g613(.A1(new_n638), .A2(new_n683), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT44), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT109), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(KEYINPUT44), .A3(new_n800), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n581), .B1(new_n582), .B2(new_n561), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n693), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(new_n584), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(KEYINPUT46), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n694), .B1(new_n808), .B2(KEYINPUT46), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n550), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n708), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n803), .A2(new_n812), .A3(new_n784), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n801), .A2(KEYINPUT109), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n802), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n811), .B(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n784), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n325), .A2(new_n633), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n725), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  NAND3_X1  g636(.A1(new_n633), .A2(new_n429), .A3(new_n550), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n742), .A2(KEYINPUT49), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n742), .A2(KEYINPUT49), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n823), .A2(new_n798), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n716), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n705), .ZN(new_n828));
  INV_X1    g642(.A(new_n421), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n799), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n756), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n745), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT115), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n819), .A2(new_n731), .A3(new_n732), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n790), .A2(new_n633), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT48), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n835), .A2(new_n836), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n835), .A2(new_n836), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n837), .A3(new_n838), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n633), .A2(new_n834), .A3(new_n827), .A4(new_n829), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n419), .B1(new_n844), .B2(new_n649), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n833), .A2(new_n841), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n697), .B1(new_n701), .B2(new_n725), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n717), .A2(new_n650), .A3(new_n667), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n684), .A2(new_n586), .A3(new_n700), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n716), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n848), .B(new_n851), .C1(new_n767), .C2(new_n776), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT52), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n546), .A2(new_n684), .A3(new_n542), .A4(new_n722), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n325), .A2(new_n666), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n774), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n781), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n782), .A2(new_n794), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(KEYINPUT111), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n785), .B1(new_n855), .B2(new_n774), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n861), .B2(new_n795), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n747), .A2(new_n734), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n738), .A2(new_n864), .A3(new_n762), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n667), .A2(new_n502), .A3(new_n546), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n797), .B2(new_n648), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n677), .A3(new_n636), .A4(new_n638), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n634), .A2(new_n685), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT110), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT110), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n634), .A2(new_n871), .A3(new_n685), .A4(new_n868), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n870), .A2(new_n872), .B1(new_n783), .B2(new_n791), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n865), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n847), .B1(new_n853), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n777), .A2(KEYINPUT52), .A3(new_n848), .A4(new_n851), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n852), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n870), .A2(new_n872), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n792), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n738), .A2(new_n864), .A3(new_n762), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n879), .A2(new_n883), .A3(KEYINPUT53), .A4(new_n863), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT54), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n733), .A2(new_n430), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT112), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n831), .A2(new_n705), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT50), .Z(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(KEYINPUT51), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n835), .A2(new_n768), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n844), .A2(new_n797), .A3(new_n648), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n831), .A2(new_n784), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n742), .A2(new_n550), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n818), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n895), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n892), .B(new_n900), .C1(new_n891), .C2(new_n890), .ZN(new_n901));
  INV_X1    g715(.A(new_n895), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n899), .B(KEYINPUT114), .Z(new_n903));
  OAI211_X1 g717(.A(new_n890), .B(new_n902), .C1(new_n903), .C2(new_n896), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT51), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n846), .B(new_n886), .C1(new_n901), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(G952), .A2(G953), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n828), .B1(new_n906), .B2(new_n907), .ZN(G75));
  NOR2_X1   g722(.A1(new_n262), .A2(G952), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n885), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n328), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n327), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n405), .A2(new_n406), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n391), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n407), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT55), .Z(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n913), .A2(KEYINPUT118), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT118), .B1(new_n913), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n910), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n913), .A2(KEYINPUT117), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT56), .B1(new_n913), .B2(KEYINPUT117), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(G51));
  NOR3_X1   g740(.A1(new_n911), .A2(new_n328), .A3(new_n807), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT119), .Z(new_n928));
  INV_X1    g742(.A(new_n886), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n584), .B(KEYINPUT57), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n692), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n909), .B1(new_n928), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(new_n485), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n485), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n909), .ZN(G60));
  AND2_X1   g750(.A1(new_n644), .A2(new_n646), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n640), .B(KEYINPUT59), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n910), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n929), .A2(new_n937), .A3(new_n938), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n875), .B2(new_n884), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n628), .B(KEYINPUT121), .Z(new_n946));
  OAI211_X1 g760(.A(KEYINPUT122), .B(new_n910), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n680), .A2(new_n681), .ZN(new_n948));
  INV_X1    g762(.A(new_n944), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n853), .A2(new_n874), .A3(new_n847), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n863), .A2(new_n865), .A3(new_n873), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT53), .B1(new_n951), .B2(new_n879), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n948), .B(new_n949), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n945), .A2(KEYINPUT120), .A3(new_n948), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n947), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT122), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n945), .A2(new_n946), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n909), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT61), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n962), .B(new_n909), .C1(new_n945), .C2(new_n948), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n945), .A2(KEYINPUT123), .A3(new_n946), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT123), .B1(new_n945), .B2(new_n946), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT124), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n960), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n947), .A2(new_n955), .A3(new_n956), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n962), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n972), .A3(new_n966), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(new_n973), .ZN(G66));
  AOI21_X1  g788(.A(new_n262), .B1(new_n423), .B2(G224), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n882), .B1(new_n872), .B2(new_n870), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n977), .B2(new_n262), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n914), .B1(G898), .B2(new_n262), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n978), .B(new_n979), .Z(G69));
  NAND3_X1  g794(.A1(new_n777), .A2(new_n720), .A3(new_n848), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n710), .A2(new_n819), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(new_n325), .A3(new_n633), .A4(new_n867), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n821), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n982), .A2(new_n985), .A3(new_n815), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n262), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n270), .A2(new_n279), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(new_n468), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n815), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n812), .A2(new_n836), .A3(new_n849), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n821), .A2(new_n858), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n792), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n777), .A2(new_n848), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n998), .A2(new_n262), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n991), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G72));
  NAND3_X1  g819(.A1(new_n998), .A2(new_n976), .A3(new_n999), .ZN(new_n1006));
  XNOR2_X1  g820(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n754), .A2(new_n328), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  AOI211_X1 g823(.A(new_n300), .B(new_n281), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n987), .B2(new_n977), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1011), .A2(new_n714), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n299), .A2(new_n301), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1009), .B1(new_n286), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT127), .Z(new_n1015));
  NOR2_X1   g829(.A1(new_n911), .A2(new_n1015), .ZN(new_n1016));
  NOR4_X1   g830(.A1(new_n1010), .A2(new_n909), .A3(new_n1012), .A4(new_n1016), .ZN(G57));
endmodule


