

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791;

  XNOR2_X1 U371 ( .A(n408), .B(n407), .ZN(n425) );
  XOR2_X1 U372 ( .A(KEYINPUT4), .B(KEYINPUT65), .Z(n772) );
  NOR2_X1 U373 ( .A1(n703), .A2(n704), .ZN(n564) );
  NAND2_X1 U374 ( .A1(n375), .A2(n372), .ZN(n790) );
  XNOR2_X2 U375 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n441) );
  NOR2_X2 U376 ( .A1(n385), .A2(n384), .ZN(n551) );
  NAND2_X2 U377 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X2 U378 ( .A(n510), .B(n355), .ZN(n773) );
  XNOR2_X2 U379 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n408) );
  XNOR2_X2 U380 ( .A(n540), .B(n539), .ZN(n708) );
  INV_X2 U381 ( .A(G953), .ZN(n412) );
  NAND2_X1 U382 ( .A1(n361), .A2(n393), .ZN(n394) );
  AND2_X1 U383 ( .A1(n788), .A2(n360), .ZN(n392) );
  AND2_X1 U384 ( .A1(n417), .A2(n416), .ZN(n415) );
  XNOR2_X1 U385 ( .A(n598), .B(KEYINPUT6), .ZN(n607) );
  XNOR2_X1 U386 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U387 ( .A(n463), .B(n462), .ZN(n592) );
  XNOR2_X1 U388 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U389 ( .A(n518), .B(n517), .ZN(n598) );
  XNOR2_X1 U390 ( .A(n659), .B(n660), .ZN(n661) );
  XNOR2_X1 U391 ( .A(n524), .B(n523), .ZN(n659) );
  NAND2_X1 U392 ( .A1(n607), .A2(n608), .ZN(n391) );
  NOR2_X1 U393 ( .A1(n352), .A2(n607), .ZN(n423) );
  NAND2_X1 U394 ( .A1(n390), .A2(n609), .ZN(n389) );
  XNOR2_X1 U395 ( .A(n391), .B(n438), .ZN(n390) );
  INV_X1 U396 ( .A(KEYINPUT104), .ZN(n438) );
  XNOR2_X1 U397 ( .A(n548), .B(n547), .ZN(n729) );
  INV_X1 U398 ( .A(KEYINPUT33), .ZN(n547) );
  INV_X1 U399 ( .A(KEYINPUT106), .ZN(n610) );
  OR2_X1 U400 ( .A1(n651), .A2(G902), .ZN(n518) );
  NAND2_X2 U401 ( .A1(n401), .A2(n400), .ZN(n546) );
  AND2_X1 U402 ( .A1(n403), .A2(n404), .ZN(n400) );
  NAND2_X1 U403 ( .A1(n370), .A2(n369), .ZN(n368) );
  INV_X1 U404 ( .A(n790), .ZN(n370) );
  NAND2_X1 U405 ( .A1(n790), .A2(n605), .ZN(n367) );
  NOR2_X1 U406 ( .A1(n556), .A2(KEYINPUT44), .ZN(n552) );
  INV_X1 U407 ( .A(G237), .ZN(n458) );
  NOR2_X1 U408 ( .A1(G953), .A2(G237), .ZN(n511) );
  NAND2_X1 U409 ( .A1(n399), .A2(n398), .ZN(n397) );
  OR2_X1 U410 ( .A1(n615), .A2(n623), .ZN(n393) );
  XNOR2_X1 U411 ( .A(G116), .B(G113), .ZN(n453) );
  NOR2_X1 U412 ( .A1(n433), .A2(n432), .ZN(n431) );
  AND2_X1 U413 ( .A1(n611), .A2(n614), .ZN(n432) );
  AND2_X1 U414 ( .A1(n387), .A2(n388), .ZN(n386) );
  NAND2_X1 U415 ( .A1(n475), .A2(KEYINPUT0), .ZN(n416) );
  OR2_X1 U416 ( .A1(n659), .A2(G902), .ZN(n380) );
  NOR2_X1 U417 ( .A1(n620), .A2(n604), .ZN(n409) );
  AND2_X1 U418 ( .A1(n630), .A2(n378), .ZN(n377) );
  NOR2_X1 U419 ( .A1(n609), .A2(KEYINPUT40), .ZN(n376) );
  OR2_X1 U420 ( .A1(n612), .A2(n435), .ZN(n434) );
  XNOR2_X1 U421 ( .A(n538), .B(n440), .ZN(n539) );
  NAND2_X1 U422 ( .A1(n546), .A2(n519), .ZN(n422) );
  INV_X1 U423 ( .A(KEYINPUT82), .ZN(n421) );
  NAND2_X1 U424 ( .A1(n366), .A2(n365), .ZN(n615) );
  NAND2_X1 U425 ( .A1(n791), .A2(n379), .ZN(n365) );
  NAND2_X1 U426 ( .A1(n368), .A2(n367), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n446), .B(G128), .ZN(n490) );
  XNOR2_X1 U428 ( .A(G131), .B(G143), .ZN(n478) );
  XOR2_X1 U429 ( .A(KEYINPUT11), .B(G104), .Z(n479) );
  XOR2_X1 U430 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n482) );
  XOR2_X1 U431 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n443) );
  INV_X1 U432 ( .A(G101), .ZN(n407) );
  NOR2_X1 U433 ( .A1(n394), .A2(n632), .ZN(n364) );
  NAND2_X1 U434 ( .A1(G234), .A2(G237), .ZN(n466) );
  INV_X1 U435 ( .A(KEYINPUT36), .ZN(n613) );
  XNOR2_X1 U436 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U437 ( .A(n524), .B(n516), .ZN(n651) );
  XNOR2_X1 U438 ( .A(KEYINPUT75), .B(G110), .ZN(n449) );
  XNOR2_X1 U439 ( .A(n477), .B(G140), .ZN(n774) );
  XNOR2_X1 U440 ( .A(n490), .B(G134), .ZN(n510) );
  XNOR2_X1 U441 ( .A(G116), .B(G107), .ZN(n491) );
  INV_X1 U442 ( .A(KEYINPUT35), .ZN(n550) );
  AND2_X1 U443 ( .A1(n729), .A2(KEYINPUT34), .ZN(n384) );
  NAND2_X1 U444 ( .A1(n414), .A2(n359), .ZN(n413) );
  NAND2_X1 U445 ( .A1(n601), .A2(n410), .ZN(n620) );
  AND2_X1 U446 ( .A1(n603), .A2(n600), .ZN(n410) );
  XNOR2_X1 U447 ( .A(n525), .B(KEYINPUT1), .ZN(n439) );
  XNOR2_X1 U448 ( .A(n406), .B(G475), .ZN(n489) );
  OR2_X1 U449 ( .A1(n640), .A2(G902), .ZN(n406) );
  AND2_X1 U450 ( .A1(n411), .A2(G953), .ZN(n763) );
  AND2_X1 U451 ( .A1(n645), .A2(G953), .ZN(n759) );
  NAND2_X1 U452 ( .A1(n374), .A2(n373), .ZN(n372) );
  NOR2_X1 U453 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U454 ( .A1(n692), .A2(n378), .ZN(n373) );
  NAND2_X1 U455 ( .A1(n351), .A2(n434), .ZN(n427) );
  XNOR2_X1 U456 ( .A(n419), .B(KEYINPUT83), .ZN(n576) );
  XNOR2_X1 U457 ( .A(n422), .B(n421), .ZN(n420) );
  AND2_X1 U458 ( .A1(n430), .A2(n362), .ZN(n351) );
  OR2_X1 U459 ( .A1(n703), .A2(n708), .ZN(n352) );
  AND2_X1 U460 ( .A1(n383), .A2(n549), .ZN(n353) );
  AND2_X1 U461 ( .A1(n622), .A2(n648), .ZN(n354) );
  OR2_X1 U462 ( .A1(n395), .A2(n394), .ZN(n776) );
  XOR2_X1 U463 ( .A(G137), .B(G131), .Z(n355) );
  XOR2_X1 U464 ( .A(n531), .B(n530), .Z(n356) );
  XNOR2_X1 U465 ( .A(n389), .B(KEYINPUT105), .ZN(n624) );
  AND2_X1 U466 ( .A1(n364), .A2(n363), .ZN(n357) );
  AND2_X1 U467 ( .A1(n430), .A2(n431), .ZN(n358) );
  NAND2_X2 U468 ( .A1(n415), .A2(n413), .ZN(n566) );
  NOR2_X1 U469 ( .A1(n475), .A2(KEYINPUT0), .ZN(n359) );
  INV_X1 U470 ( .A(n626), .ZN(n433) );
  AND2_X1 U471 ( .A1(n354), .A2(n623), .ZN(n360) );
  AND2_X1 U472 ( .A1(n649), .A2(n698), .ZN(n361) );
  INV_X1 U473 ( .A(n609), .ZN(n692) );
  AND2_X1 U474 ( .A1(n570), .A2(n569), .ZN(n609) );
  AND2_X1 U475 ( .A1(n431), .A2(n428), .ZN(n362) );
  XNOR2_X1 U476 ( .A(n457), .B(n459), .ZN(n632) );
  INV_X1 U477 ( .A(n395), .ZN(n363) );
  NAND2_X1 U478 ( .A1(n371), .A2(n605), .ZN(n369) );
  INV_X1 U479 ( .A(n791), .ZN(n371) );
  INV_X1 U480 ( .A(n630), .ZN(n374) );
  INV_X1 U481 ( .A(KEYINPUT40), .ZN(n378) );
  INV_X1 U482 ( .A(n605), .ZN(n379) );
  XNOR2_X2 U483 ( .A(n559), .B(n439), .ZN(n703) );
  XNOR2_X2 U484 ( .A(n380), .B(G469), .ZN(n559) );
  INV_X1 U485 ( .A(n566), .ZN(n383) );
  INV_X1 U486 ( .A(n729), .ZN(n382) );
  NAND2_X1 U487 ( .A1(n381), .A2(n386), .ZN(n385) );
  NAND2_X1 U488 ( .A1(n382), .A2(n353), .ZN(n381) );
  NAND2_X1 U489 ( .A1(n566), .A2(KEYINPUT34), .ZN(n387) );
  INV_X1 U490 ( .A(n619), .ZN(n388) );
  NAND2_X1 U491 ( .A1(n788), .A2(n354), .ZN(n399) );
  NAND2_X1 U492 ( .A1(n392), .A2(n615), .ZN(n396) );
  NAND2_X1 U493 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U494 ( .A(n623), .ZN(n398) );
  XNOR2_X1 U495 ( .A(n557), .B(KEYINPUT84), .ZN(n554) );
  NOR2_X2 U496 ( .A1(n650), .A2(n682), .ZN(n557) );
  NAND2_X1 U497 ( .A1(n566), .A2(n508), .ZN(n403) );
  NAND2_X1 U498 ( .A1(n546), .A2(n423), .ZN(n542) );
  NAND2_X1 U499 ( .A1(n402), .A2(n418), .ZN(n401) );
  NOR2_X1 U500 ( .A1(n566), .A2(n508), .ZN(n402) );
  NAND2_X1 U501 ( .A1(n507), .A2(n508), .ZN(n404) );
  NOR2_X1 U502 ( .A1(n741), .A2(n616), .ZN(n596) );
  XNOR2_X1 U503 ( .A(n595), .B(KEYINPUT41), .ZN(n741) );
  BUF_X1 U504 ( .A(n688), .Z(n405) );
  XNOR2_X1 U505 ( .A(n409), .B(KEYINPUT39), .ZN(n630) );
  NAND2_X1 U506 ( .A1(n412), .A2(G224), .ZN(n442) );
  NAND2_X1 U507 ( .A1(n412), .A2(G234), .ZN(n497) );
  NAND2_X1 U508 ( .A1(n412), .A2(G227), .ZN(n520) );
  INV_X1 U509 ( .A(G898), .ZN(n411) );
  NOR2_X1 U510 ( .A1(n781), .A2(n412), .ZN(n782) );
  NAND2_X1 U511 ( .A1(n700), .A2(n412), .ZN(n769) );
  INV_X1 U512 ( .A(n688), .ZN(n414) );
  NAND2_X1 U513 ( .A1(n688), .A2(KEYINPUT0), .ZN(n417) );
  XNOR2_X2 U514 ( .A(n611), .B(n465), .ZN(n688) );
  INV_X1 U515 ( .A(n507), .ZN(n418) );
  NAND2_X1 U516 ( .A1(n420), .A2(n433), .ZN(n419) );
  AND2_X2 U517 ( .A1(n699), .A2(n583), .ZN(n631) );
  NAND2_X2 U518 ( .A1(n592), .A2(n720), .ZN(n611) );
  XNOR2_X2 U519 ( .A(n424), .B(n773), .ZN(n524) );
  XNOR2_X2 U520 ( .A(n509), .B(G146), .ZN(n424) );
  XNOR2_X2 U521 ( .A(n425), .B(n772), .ZN(n509) );
  NAND2_X1 U522 ( .A1(n426), .A2(KEYINPUT108), .ZN(n429) );
  NAND2_X1 U523 ( .A1(n358), .A2(n434), .ZN(n426) );
  NAND2_X2 U524 ( .A1(n429), .A2(n427), .ZN(n788) );
  INV_X1 U525 ( .A(KEYINPUT108), .ZN(n428) );
  NAND2_X1 U526 ( .A1(n612), .A2(n614), .ZN(n430) );
  NAND2_X1 U527 ( .A1(n436), .A2(n437), .ZN(n435) );
  INV_X1 U528 ( .A(n611), .ZN(n436) );
  INV_X1 U529 ( .A(n614), .ZN(n437) );
  XNOR2_X1 U530 ( .A(n551), .B(n550), .ZN(n556) );
  XOR2_X1 U531 ( .A(n537), .B(n536), .Z(n440) );
  BUF_X1 U532 ( .A(n729), .Z(n740) );
  XNOR2_X1 U533 ( .A(n613), .B(KEYINPUT107), .ZN(n614) );
  BUF_X1 U534 ( .A(n750), .Z(n755) );
  XNOR2_X1 U535 ( .A(n751), .B(KEYINPUT122), .ZN(n752) );
  XNOR2_X1 U536 ( .A(n753), .B(n752), .ZN(n754) );
  XNOR2_X1 U537 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n444), .B(n443), .ZN(n448) );
  INV_X1 U539 ( .A(G146), .ZN(n445) );
  XNOR2_X1 U540 ( .A(n445), .B(G125), .ZN(n476) );
  INV_X1 U541 ( .A(G143), .ZN(n446) );
  XNOR2_X1 U542 ( .A(n490), .B(n476), .ZN(n447) );
  XNOR2_X1 U543 ( .A(n448), .B(n447), .ZN(n451) );
  XOR2_X1 U544 ( .A(G104), .B(G107), .Z(n450) );
  XNOR2_X1 U545 ( .A(n450), .B(n449), .ZN(n760) );
  XNOR2_X1 U546 ( .A(n760), .B(KEYINPUT73), .ZN(n522) );
  XNOR2_X1 U547 ( .A(n451), .B(n522), .ZN(n456) );
  XNOR2_X1 U548 ( .A(KEYINPUT3), .B(G119), .ZN(n452) );
  XNOR2_X1 U549 ( .A(n453), .B(n452), .ZN(n514) );
  XNOR2_X1 U550 ( .A(KEYINPUT16), .B(G122), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n514), .B(n454), .ZN(n761) );
  XNOR2_X1 U552 ( .A(n509), .B(n761), .ZN(n455) );
  XNOR2_X1 U553 ( .A(n456), .B(n455), .ZN(n665) );
  XNOR2_X1 U554 ( .A(KEYINPUT87), .B(KEYINPUT15), .ZN(n457) );
  INV_X1 U555 ( .A(G902), .ZN(n459) );
  NAND2_X1 U556 ( .A1(n665), .A2(n632), .ZN(n463) );
  NAND2_X1 U557 ( .A1(n459), .A2(n458), .ZN(n464) );
  NAND2_X1 U558 ( .A1(n464), .A2(G210), .ZN(n461) );
  INV_X1 U559 ( .A(KEYINPUT90), .ZN(n460) );
  NAND2_X1 U560 ( .A1(n464), .A2(G214), .ZN(n720) );
  INV_X1 U561 ( .A(KEYINPUT19), .ZN(n465) );
  XNOR2_X1 U562 ( .A(n466), .B(KEYINPUT14), .ZN(n470) );
  NAND2_X1 U563 ( .A1(n470), .A2(G952), .ZN(n467) );
  XOR2_X1 U564 ( .A(KEYINPUT91), .B(n467), .Z(n736) );
  NOR2_X1 U565 ( .A1(G953), .A2(n736), .ZN(n469) );
  INV_X1 U566 ( .A(KEYINPUT92), .ZN(n468) );
  XNOR2_X1 U567 ( .A(n469), .B(n468), .ZN(n588) );
  NAND2_X1 U568 ( .A1(G902), .A2(n470), .ZN(n585) );
  INV_X1 U569 ( .A(n585), .ZN(n471) );
  NAND2_X1 U570 ( .A1(n471), .A2(n763), .ZN(n473) );
  INV_X1 U571 ( .A(KEYINPUT93), .ZN(n472) );
  XNOR2_X1 U572 ( .A(n473), .B(n472), .ZN(n474) );
  AND2_X1 U573 ( .A1(n588), .A2(n474), .ZN(n475) );
  XNOR2_X1 U574 ( .A(n476), .B(KEYINPUT10), .ZN(n477) );
  XNOR2_X1 U575 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n774), .B(n480), .ZN(n487) );
  NAND2_X1 U577 ( .A1(G214), .A2(n511), .ZN(n481) );
  XNOR2_X1 U578 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U579 ( .A(n483), .B(KEYINPUT100), .Z(n485) );
  XNOR2_X1 U580 ( .A(G113), .B(G122), .ZN(n484) );
  XNOR2_X1 U581 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U582 ( .A(n487), .B(n486), .ZN(n640) );
  INV_X1 U583 ( .A(KEYINPUT13), .ZN(n488) );
  XNOR2_X1 U584 ( .A(n489), .B(n488), .ZN(n570) );
  XOR2_X1 U585 ( .A(KEYINPUT102), .B(G122), .Z(n492) );
  XNOR2_X1 U586 ( .A(n492), .B(n491), .ZN(n496) );
  XOR2_X1 U587 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n494) );
  XNOR2_X1 U588 ( .A(KEYINPUT9), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U589 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U590 ( .A(n496), .B(n495), .Z(n499) );
  XOR2_X1 U591 ( .A(KEYINPUT8), .B(n497), .Z(n532) );
  NAND2_X1 U592 ( .A1(G217), .A2(n532), .ZN(n498) );
  XNOR2_X1 U593 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U594 ( .A(n510), .B(n500), .ZN(n751) );
  NOR2_X1 U595 ( .A1(n751), .A2(G902), .ZN(n502) );
  INV_X1 U596 ( .A(G478), .ZN(n501) );
  XNOR2_X1 U597 ( .A(n502), .B(n501), .ZN(n571) );
  NOR2_X1 U598 ( .A1(n570), .A2(n571), .ZN(n594) );
  NAND2_X1 U599 ( .A1(n632), .A2(G234), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n503), .B(KEYINPUT20), .ZN(n535) );
  NAND2_X1 U601 ( .A1(n535), .A2(G221), .ZN(n506) );
  INV_X1 U602 ( .A(KEYINPUT96), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n504), .B(KEYINPUT21), .ZN(n505) );
  XNOR2_X1 U604 ( .A(n506), .B(n505), .ZN(n707) );
  NAND2_X1 U605 ( .A1(n594), .A2(n707), .ZN(n507) );
  INV_X1 U606 ( .A(KEYINPUT22), .ZN(n508) );
  XOR2_X1 U607 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n513) );
  NAND2_X1 U608 ( .A1(n511), .A2(G210), .ZN(n512) );
  XNOR2_X1 U609 ( .A(n513), .B(n512), .ZN(n515) );
  XNOR2_X1 U610 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U611 ( .A(G472), .ZN(n517) );
  INV_X1 U612 ( .A(n607), .ZN(n519) );
  XNOR2_X1 U613 ( .A(n520), .B(G140), .ZN(n521) );
  XNOR2_X1 U614 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U615 ( .A(KEYINPUT68), .ZN(n525) );
  XOR2_X1 U616 ( .A(G110), .B(G128), .Z(n527) );
  XNOR2_X1 U617 ( .A(G119), .B(G137), .ZN(n526) );
  XNOR2_X1 U618 ( .A(n527), .B(n526), .ZN(n531) );
  XOR2_X1 U619 ( .A(KEYINPUT78), .B(KEYINPUT94), .Z(n529) );
  XNOR2_X1 U620 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n528) );
  XNOR2_X1 U621 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U622 ( .A1(G221), .A2(n532), .ZN(n533) );
  XNOR2_X1 U623 ( .A(n356), .B(n533), .ZN(n534) );
  XNOR2_X1 U624 ( .A(n534), .B(n774), .ZN(n756) );
  NOR2_X1 U625 ( .A1(n756), .A2(G902), .ZN(n540) );
  NAND2_X1 U626 ( .A1(G217), .A2(n535), .ZN(n538) );
  XOR2_X1 U627 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n537) );
  XNOR2_X1 U628 ( .A(KEYINPUT25), .B(KEYINPUT95), .ZN(n536) );
  XNOR2_X1 U629 ( .A(KEYINPUT67), .B(KEYINPUT32), .ZN(n541) );
  XNOR2_X1 U630 ( .A(n542), .B(n541), .ZN(n650) );
  INV_X1 U631 ( .A(n598), .ZN(n561) );
  INV_X1 U632 ( .A(n561), .ZN(n714) );
  INV_X1 U633 ( .A(n708), .ZN(n543) );
  AND2_X1 U634 ( .A1(n714), .A2(n543), .ZN(n544) );
  AND2_X1 U635 ( .A1(n703), .A2(n544), .ZN(n545) );
  AND2_X1 U636 ( .A1(n546), .A2(n545), .ZN(n682) );
  NAND2_X1 U637 ( .A1(n708), .A2(n707), .ZN(n704) );
  NAND2_X1 U638 ( .A1(n564), .A2(n607), .ZN(n548) );
  INV_X1 U639 ( .A(KEYINPUT34), .ZN(n549) );
  NAND2_X1 U640 ( .A1(n570), .A2(n571), .ZN(n619) );
  XNOR2_X1 U641 ( .A(n552), .B(KEYINPUT72), .ZN(n553) );
  NAND2_X1 U642 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U643 ( .A(n555), .B(KEYINPUT74), .ZN(n580) );
  INV_X1 U644 ( .A(n556), .ZN(n786) );
  NAND2_X1 U645 ( .A1(n786), .A2(n557), .ZN(n558) );
  NAND2_X1 U646 ( .A1(n558), .A2(KEYINPUT44), .ZN(n575) );
  INV_X1 U647 ( .A(n704), .ZN(n560) );
  NAND2_X1 U648 ( .A1(n559), .A2(n560), .ZN(n602) );
  NOR2_X1 U649 ( .A1(n602), .A2(n561), .ZN(n562) );
  NAND2_X1 U650 ( .A1(n383), .A2(n562), .ZN(n563) );
  XNOR2_X1 U651 ( .A(KEYINPUT98), .B(n563), .ZN(n676) );
  INV_X1 U652 ( .A(n564), .ZN(n565) );
  OR2_X1 U653 ( .A1(n714), .A2(n565), .ZN(n715) );
  OR2_X1 U654 ( .A1(n566), .A2(n715), .ZN(n568) );
  INV_X1 U655 ( .A(KEYINPUT31), .ZN(n567) );
  XNOR2_X1 U656 ( .A(n568), .B(n567), .ZN(n694) );
  NAND2_X1 U657 ( .A1(n676), .A2(n694), .ZN(n573) );
  INV_X1 U658 ( .A(n571), .ZN(n569) );
  INV_X1 U659 ( .A(n570), .ZN(n572) );
  NAND2_X1 U660 ( .A1(n572), .A2(n571), .ZN(n695) );
  NAND2_X1 U661 ( .A1(n692), .A2(n695), .ZN(n724) );
  NAND2_X1 U662 ( .A1(n573), .A2(n724), .ZN(n574) );
  NAND2_X1 U663 ( .A1(n575), .A2(n574), .ZN(n578) );
  INV_X1 U664 ( .A(n703), .ZN(n626) );
  NAND2_X1 U665 ( .A1(n576), .A2(n708), .ZN(n672) );
  INV_X1 U666 ( .A(n672), .ZN(n577) );
  NOR2_X1 U667 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U668 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X2 U669 ( .A(n581), .B(KEYINPUT45), .ZN(n699) );
  NOR2_X1 U670 ( .A1(n632), .A2(KEYINPUT80), .ZN(n582) );
  OR2_X1 U671 ( .A1(n582), .A2(KEYINPUT2), .ZN(n583) );
  INV_X1 U672 ( .A(n707), .ZN(n584) );
  NOR2_X1 U673 ( .A1(n708), .A2(n584), .ZN(n589) );
  NOR2_X1 U674 ( .A1(G900), .A2(n585), .ZN(n586) );
  NAND2_X1 U675 ( .A1(G953), .A2(n586), .ZN(n587) );
  NAND2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n589), .A2(n600), .ZN(n606) );
  NOR2_X1 U678 ( .A1(n606), .A2(n714), .ZN(n590) );
  XNOR2_X1 U679 ( .A(KEYINPUT28), .B(n590), .ZN(n591) );
  NAND2_X1 U680 ( .A1(n591), .A2(n559), .ZN(n616) );
  BUF_X1 U681 ( .A(n592), .Z(n593) );
  XNOR2_X1 U682 ( .A(n593), .B(KEYINPUT38), .ZN(n604) );
  INV_X1 U683 ( .A(n604), .ZN(n721) );
  NAND2_X1 U684 ( .A1(n721), .A2(n720), .ZN(n725) );
  INV_X1 U685 ( .A(n594), .ZN(n723) );
  NOR2_X1 U686 ( .A1(n725), .A2(n723), .ZN(n595) );
  XNOR2_X1 U687 ( .A(n596), .B(KEYINPUT42), .ZN(n791) );
  INV_X1 U688 ( .A(n720), .ZN(n597) );
  OR2_X1 U689 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U690 ( .A(KEYINPUT30), .B(n599), .Z(n601) );
  INV_X1 U691 ( .A(n602), .ZN(n603) );
  XNOR2_X1 U692 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n605) );
  INV_X1 U693 ( .A(n606), .ZN(n608) );
  XNOR2_X1 U694 ( .A(n624), .B(n610), .ZN(n612) );
  INV_X1 U695 ( .A(n616), .ZN(n687) );
  NAND2_X1 U696 ( .A1(n687), .A2(n724), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n617), .A2(n405), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n618), .B(KEYINPUT47), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n621), .A2(n593), .ZN(n648) );
  XNOR2_X1 U701 ( .A(KEYINPUT48), .B(KEYINPUT81), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n720), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U704 ( .A(n627), .B(KEYINPUT43), .Z(n629) );
  INV_X1 U705 ( .A(n593), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n649) );
  OR2_X1 U707 ( .A1(n630), .A2(n695), .ZN(n698) );
  INV_X1 U708 ( .A(n776), .ZN(n701) );
  NAND2_X1 U709 ( .A1(n631), .A2(n701), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n699), .A2(n357), .ZN(n635) );
  OR2_X1 U711 ( .A1(n632), .A2(n738), .ZN(n633) );
  AND2_X1 U712 ( .A1(n633), .A2(KEYINPUT80), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  INV_X1 U714 ( .A(KEYINPUT66), .ZN(n638) );
  XNOR2_X2 U715 ( .A(n639), .B(n638), .ZN(n750) );
  NAND2_X1 U716 ( .A1(n750), .A2(G475), .ZN(n644) );
  XOR2_X1 U717 ( .A(KEYINPUT69), .B(KEYINPUT59), .Z(n642) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT121), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(n646) );
  INV_X1 U720 ( .A(G952), .ZN(n645) );
  NOR2_X2 U721 ( .A1(n646), .A2(n759), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n647), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U723 ( .A(n648), .B(G143), .ZN(G45) );
  XNOR2_X1 U724 ( .A(n649), .B(G140), .ZN(G42) );
  XOR2_X1 U725 ( .A(n650), .B(G119), .Z(G21) );
  NAND2_X1 U726 ( .A1(n750), .A2(G472), .ZN(n654) );
  XNOR2_X1 U727 ( .A(KEYINPUT86), .B(KEYINPUT62), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n651), .B(n652), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X2 U730 ( .A1(n655), .A2(n759), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT109), .B(KEYINPUT63), .ZN(n656) );
  XOR2_X1 U732 ( .A(n656), .B(KEYINPUT85), .Z(n657) );
  XNOR2_X1 U733 ( .A(n658), .B(n657), .ZN(G57) );
  NAND2_X1 U734 ( .A1(n750), .A2(G469), .ZN(n662) );
  XOR2_X1 U735 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n660) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X2 U737 ( .A1(n663), .A2(n759), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n664), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U739 ( .A1(n750), .A2(G210), .ZN(n669) );
  BUF_X1 U740 ( .A(n665), .Z(n667) );
  XNOR2_X1 U741 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X2 U743 ( .A1(n670), .A2(n759), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U745 ( .A(G101), .B(KEYINPUT110), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(G3) );
  NOR2_X1 U747 ( .A1(n676), .A2(n692), .ZN(n675) );
  XNOR2_X1 U748 ( .A(G104), .B(KEYINPUT111), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n675), .B(n674), .ZN(G6) );
  NOR2_X1 U750 ( .A1(n676), .A2(n695), .ZN(n681) );
  XOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n678) );
  XNOR2_X1 U752 ( .A(G107), .B(KEYINPUT26), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U754 ( .A(KEYINPUT112), .B(n679), .ZN(n680) );
  XNOR2_X1 U755 ( .A(n681), .B(n680), .ZN(G9) );
  XOR2_X1 U756 ( .A(G110), .B(n682), .Z(G12) );
  INV_X1 U757 ( .A(n695), .ZN(n683) );
  NAND2_X1 U758 ( .A1(n687), .A2(n683), .ZN(n684) );
  NOR2_X1 U759 ( .A1(n684), .A2(n405), .ZN(n686) );
  XNOR2_X1 U760 ( .A(G128), .B(KEYINPUT29), .ZN(n685) );
  XNOR2_X1 U761 ( .A(n686), .B(n685), .ZN(G30) );
  NAND2_X1 U762 ( .A1(n687), .A2(n609), .ZN(n689) );
  NOR2_X1 U763 ( .A1(n689), .A2(n405), .ZN(n690) );
  XOR2_X1 U764 ( .A(KEYINPUT114), .B(n690), .Z(n691) );
  XNOR2_X1 U765 ( .A(G146), .B(n691), .ZN(G48) );
  NOR2_X1 U766 ( .A1(n692), .A2(n694), .ZN(n693) );
  XOR2_X1 U767 ( .A(G113), .B(n693), .Z(G15) );
  NOR2_X1 U768 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U769 ( .A(G116), .B(KEYINPUT115), .ZN(n696) );
  XNOR2_X1 U770 ( .A(n697), .B(n696), .ZN(G18) );
  XNOR2_X1 U771 ( .A(G134), .B(n698), .ZN(G36) );
  BUF_X1 U772 ( .A(n699), .Z(n700) );
  NAND2_X1 U773 ( .A1(n701), .A2(n700), .ZN(n737) );
  NOR2_X1 U774 ( .A1(n738), .A2(KEYINPUT79), .ZN(n702) );
  NAND2_X1 U775 ( .A1(n737), .A2(n702), .ZN(n748) );
  NAND2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U777 ( .A(n705), .B(KEYINPUT50), .ZN(n706) );
  XNOR2_X1 U778 ( .A(KEYINPUT117), .B(n706), .ZN(n712) );
  NOR2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U780 ( .A(KEYINPUT49), .B(n709), .Z(n710) );
  XNOR2_X1 U781 ( .A(KEYINPUT116), .B(n710), .ZN(n711) );
  NOR2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n717), .B(KEYINPUT118), .ZN(n718) );
  XNOR2_X1 U786 ( .A(n718), .B(KEYINPUT51), .ZN(n719) );
  NOR2_X1 U787 ( .A1(n741), .A2(n719), .ZN(n733) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n728) );
  INV_X1 U790 ( .A(n724), .ZN(n726) );
  NOR2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U792 ( .A1(n728), .A2(n727), .ZN(n730) );
  NOR2_X1 U793 ( .A1(n730), .A2(n740), .ZN(n731) );
  XOR2_X1 U794 ( .A(KEYINPUT119), .B(n731), .Z(n732) );
  NOR2_X1 U795 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U796 ( .A(n734), .B(KEYINPUT52), .ZN(n735) );
  NOR2_X1 U797 ( .A1(n736), .A2(n735), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n737), .B(KEYINPUT79), .ZN(n739) );
  INV_X1 U799 ( .A(KEYINPUT2), .ZN(n738) );
  NAND2_X1 U800 ( .A1(n739), .A2(n738), .ZN(n744) );
  NOR2_X1 U801 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U802 ( .A1(G953), .A2(n742), .ZN(n743) );
  NAND2_X1 U803 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U804 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U805 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U806 ( .A(KEYINPUT53), .B(n749), .Z(G75) );
  NAND2_X1 U807 ( .A1(n755), .A2(G478), .ZN(n753) );
  NOR2_X1 U808 ( .A1(n759), .A2(n754), .ZN(G63) );
  NAND2_X1 U809 ( .A1(n755), .A2(G217), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n757), .B(n756), .ZN(n758) );
  NOR2_X1 U811 ( .A1(n759), .A2(n758), .ZN(G66) );
  XOR2_X1 U812 ( .A(G101), .B(n760), .Z(n762) );
  XNOR2_X1 U813 ( .A(n762), .B(n761), .ZN(n765) );
  INV_X1 U814 ( .A(n763), .ZN(n764) );
  AND2_X1 U815 ( .A1(n765), .A2(n764), .ZN(n771) );
  NAND2_X1 U816 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n766), .B(KEYINPUT61), .ZN(n767) );
  NAND2_X1 U818 ( .A1(n767), .A2(G898), .ZN(n768) );
  NAND2_X1 U819 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U820 ( .A(n771), .B(n770), .ZN(G69) );
  XNOR2_X1 U821 ( .A(n772), .B(n773), .ZN(n775) );
  XNOR2_X1 U822 ( .A(n775), .B(n774), .ZN(n778) );
  XOR2_X1 U823 ( .A(n778), .B(n776), .Z(n777) );
  NOR2_X1 U824 ( .A1(G953), .A2(n777), .ZN(n784) );
  XNOR2_X1 U825 ( .A(G227), .B(n778), .ZN(n779) );
  NAND2_X1 U826 ( .A1(n779), .A2(G900), .ZN(n780) );
  XNOR2_X1 U827 ( .A(KEYINPUT123), .B(n780), .ZN(n781) );
  XNOR2_X1 U828 ( .A(n782), .B(KEYINPUT124), .ZN(n783) );
  NOR2_X1 U829 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U830 ( .A(KEYINPUT125), .B(n785), .ZN(G72) );
  XNOR2_X1 U831 ( .A(G122), .B(KEYINPUT126), .ZN(n787) );
  XNOR2_X1 U832 ( .A(n787), .B(n786), .ZN(G24) );
  XOR2_X1 U833 ( .A(n788), .B(G125), .Z(n789) );
  XNOR2_X1 U834 ( .A(KEYINPUT37), .B(n789), .ZN(G27) );
  XOR2_X1 U835 ( .A(G131), .B(n790), .Z(G33) );
  XOR2_X1 U836 ( .A(G137), .B(n791), .Z(G39) );
endmodule

