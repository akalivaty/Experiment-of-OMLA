

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767;

  NOR2_X1 U371 ( .A1(n375), .A2(n372), .ZN(n367) );
  XNOR2_X1 U372 ( .A(n585), .B(KEYINPUT35), .ZN(n651) );
  XNOR2_X1 U373 ( .A(n551), .B(KEYINPUT40), .ZN(n764) );
  BUF_X1 U374 ( .A(n677), .Z(n350) );
  XNOR2_X1 U375 ( .A(n541), .B(KEYINPUT1), .ZN(n677) );
  XNOR2_X1 U376 ( .A(n450), .B(n449), .ZN(n541) );
  OR2_X1 U377 ( .A1(n720), .A2(G902), .ZN(n450) );
  XNOR2_X1 U378 ( .A(n749), .B(n442), .ZN(n467) );
  XNOR2_X1 U379 ( .A(KEYINPUT68), .B(G101), .ZN(n502) );
  INV_X1 U380 ( .A(G146), .ZN(n424) );
  XNOR2_X2 U381 ( .A(n507), .B(n353), .ZN(n749) );
  NOR2_X2 U382 ( .A1(n647), .A2(n733), .ZN(n649) );
  XNOR2_X1 U383 ( .A(n387), .B(KEYINPUT46), .ZN(n557) );
  NOR2_X1 U384 ( .A1(n583), .A2(n582), .ZN(n698) );
  XNOR2_X2 U385 ( .A(n521), .B(n520), .ZN(n578) );
  XNOR2_X2 U386 ( .A(n393), .B(n420), .ZN(n519) );
  XNOR2_X2 U387 ( .A(n409), .B(n362), .ZN(n599) );
  XNOR2_X2 U388 ( .A(n490), .B(n441), .ZN(n507) );
  XNOR2_X2 U389 ( .A(n395), .B(n394), .ZN(n527) );
  XNOR2_X2 U390 ( .A(G110), .B(G107), .ZN(n443) );
  INV_X2 U391 ( .A(G953), .ZN(n741) );
  INV_X1 U392 ( .A(KEYINPUT80), .ZN(n394) );
  NAND2_X1 U393 ( .A1(n379), .A2(n412), .ZN(n378) );
  AND2_X1 U394 ( .A1(n565), .A2(n351), .ZN(n399) );
  XNOR2_X1 U395 ( .A(n594), .B(n593), .ZN(n673) );
  XNOR2_X1 U396 ( .A(n407), .B(n406), .ZN(n712) );
  NAND2_X1 U397 ( .A1(n599), .A2(n356), .ZN(n601) );
  AND2_X1 U398 ( .A1(n537), .A2(n536), .ZN(n561) );
  BUF_X1 U399 ( .A(n615), .Z(n604) );
  NAND2_X2 U400 ( .A1(n652), .A2(n667), .ZN(n411) );
  NAND2_X1 U401 ( .A1(n398), .A2(n400), .ZN(n746) );
  XNOR2_X2 U402 ( .A(n501), .B(n500), .ZN(n740) );
  INV_X1 U403 ( .A(KEYINPUT10), .ZN(n425) );
  INV_X1 U404 ( .A(n417), .ZN(n416) );
  XNOR2_X1 U405 ( .A(n382), .B(n354), .ZN(n615) );
  OR2_X1 U406 ( .A1(n729), .A2(G902), .ZN(n382) );
  NAND2_X1 U407 ( .A1(n764), .A2(n767), .ZN(n387) );
  AND2_X1 U408 ( .A1(n651), .A2(KEYINPUT44), .ZN(n608) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n469) );
  XNOR2_X1 U410 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n475) );
  XOR2_X1 U411 ( .A(KEYINPUT97), .B(KEYINPUT99), .Z(n474) );
  INV_X1 U412 ( .A(n650), .ZN(n402) );
  XNOR2_X1 U413 ( .A(n574), .B(n573), .ZN(n702) );
  NAND2_X1 U414 ( .A1(n578), .A2(n577), .ZN(n409) );
  XNOR2_X1 U415 ( .A(n471), .B(n426), .ZN(n747) );
  XNOR2_X1 U416 ( .A(G119), .B(G128), .ZN(n422) );
  XOR2_X1 U417 ( .A(KEYINPUT77), .B(G110), .Z(n423) );
  XNOR2_X1 U418 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n428) );
  NAND2_X1 U419 ( .A1(n380), .A2(KEYINPUT2), .ZN(n379) );
  NAND2_X1 U420 ( .A1(n417), .A2(n414), .ZN(n413) );
  BUF_X1 U421 ( .A(n563), .Z(n386) );
  INV_X1 U422 ( .A(KEYINPUT41), .ZN(n406) );
  XNOR2_X1 U423 ( .A(n549), .B(n548), .ZN(n567) );
  INV_X1 U424 ( .A(KEYINPUT39), .ZN(n548) );
  AND2_X1 U425 ( .A1(n547), .A2(n546), .ZN(n549) );
  NAND2_X1 U426 ( .A1(n702), .A2(n590), .ZN(n581) );
  NAND2_X1 U427 ( .A1(n384), .A2(n383), .ZN(n688) );
  AND2_X1 U428 ( .A1(n683), .A2(n592), .ZN(n383) );
  XNOR2_X1 U429 ( .A(n484), .B(n391), .ZN(n583) );
  XNOR2_X1 U430 ( .A(n485), .B(n392), .ZN(n391) );
  XNOR2_X1 U431 ( .A(n644), .B(KEYINPUT62), .ZN(n645) );
  XNOR2_X1 U432 ( .A(n640), .B(n639), .ZN(n733) );
  INV_X1 U433 ( .A(KEYINPUT85), .ZN(n410) );
  XNOR2_X1 U434 ( .A(KEYINPUT5), .B(G137), .ZN(n459) );
  XNOR2_X1 U435 ( .A(KEYINPUT70), .B(G131), .ZN(n479) );
  XNOR2_X1 U436 ( .A(G113), .B(G143), .ZN(n473) );
  XOR2_X1 U437 ( .A(G137), .B(G140), .Z(n444) );
  XNOR2_X1 U438 ( .A(G116), .B(G113), .ZN(n464) );
  XNOR2_X1 U439 ( .A(KEYINPUT3), .B(G119), .ZN(n463) );
  NOR2_X1 U440 ( .A1(n352), .A2(n365), .ZN(n417) );
  AND2_X1 U441 ( .A1(n587), .A2(n680), .ZN(n518) );
  NOR2_X1 U442 ( .A1(n615), .A2(n517), .ZN(n531) );
  XNOR2_X1 U443 ( .A(n552), .B(n408), .ZN(n693) );
  INV_X1 U444 ( .A(KEYINPUT108), .ZN(n408) );
  XNOR2_X1 U445 ( .A(n563), .B(KEYINPUT38), .ZN(n696) );
  OR2_X1 U446 ( .A1(n565), .A2(n401), .ZN(n400) );
  NOR2_X1 U447 ( .A1(n399), .A2(n360), .ZN(n398) );
  XOR2_X1 U448 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n487) );
  XNOR2_X1 U449 ( .A(G116), .B(G134), .ZN(n486) );
  XNOR2_X1 U450 ( .A(n443), .B(G104), .ZN(n499) );
  XNOR2_X1 U451 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n441) );
  XNOR2_X1 U452 ( .A(n499), .B(n498), .ZN(n501) );
  XNOR2_X1 U453 ( .A(KEYINPUT16), .B(G122), .ZN(n498) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n545) );
  INV_X1 U455 ( .A(KEYINPUT30), .ZN(n388) );
  INV_X1 U456 ( .A(KEYINPUT6), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n385), .B(n432), .ZN(n729) );
  XNOR2_X1 U458 ( .A(n431), .B(n359), .ZN(n432) );
  XNOR2_X1 U459 ( .A(n747), .B(n433), .ZN(n385) );
  NAND2_X1 U460 ( .A1(n371), .A2(n370), .ZN(n655) );
  NOR2_X1 U461 ( .A1(n378), .A2(n392), .ZN(n371) );
  INV_X1 U462 ( .A(G210), .ZN(n373) );
  AND2_X1 U463 ( .A1(n564), .A2(n386), .ZN(n650) );
  NOR2_X1 U464 ( .A1(n712), .A2(n554), .ZN(n556) );
  NAND2_X1 U465 ( .A1(n567), .A2(n671), .ZN(n551) );
  XNOR2_X1 U466 ( .A(n543), .B(KEYINPUT111), .ZN(n759) );
  NAND2_X1 U467 ( .A1(n584), .A2(n419), .ZN(n585) );
  XNOR2_X1 U468 ( .A(n581), .B(n580), .ZN(n584) );
  OR2_X1 U469 ( .A1(n688), .A2(n598), .ZN(n594) );
  NOR2_X1 U470 ( .A1(n566), .A2(n527), .ZN(n668) );
  XNOR2_X1 U471 ( .A(n591), .B(n381), .ZN(n662) );
  INV_X1 U472 ( .A(KEYINPUT94), .ZN(n381) );
  NOR2_X1 U473 ( .A1(n766), .A2(KEYINPUT82), .ZN(n351) );
  NOR2_X1 U474 ( .A1(n631), .A2(n630), .ZN(n352) );
  INV_X1 U475 ( .A(KEYINPUT66), .ZN(n418) );
  XOR2_X1 U476 ( .A(n479), .B(G134), .Z(n353) );
  XNOR2_X1 U477 ( .A(n437), .B(n436), .ZN(n354) );
  OR2_X1 U478 ( .A1(G237), .A2(G902), .ZN(n355) );
  AND2_X1 U479 ( .A1(n698), .A2(n680), .ZN(n356) );
  NAND2_X1 U480 ( .A1(n628), .A2(n627), .ZN(n357) );
  AND2_X1 U481 ( .A1(n650), .A2(n403), .ZN(n358) );
  XOR2_X1 U482 ( .A(n430), .B(n429), .Z(n359) );
  INV_X1 U483 ( .A(n677), .ZN(n384) );
  AND2_X1 U484 ( .A1(n358), .A2(n569), .ZN(n360) );
  INV_X1 U485 ( .A(n378), .ZN(n368) );
  AND2_X1 U486 ( .A1(n402), .A2(KEYINPUT82), .ZN(n361) );
  XOR2_X1 U487 ( .A(n579), .B(KEYINPUT0), .Z(n362) );
  AND2_X1 U488 ( .A1(n631), .A2(n418), .ZN(n363) );
  NOR2_X1 U489 ( .A1(n633), .A2(KEYINPUT81), .ZN(n364) );
  AND2_X1 U490 ( .A1(n364), .A2(n631), .ZN(n365) );
  XNOR2_X1 U491 ( .A(G902), .B(KEYINPUT15), .ZN(n629) );
  AND2_X1 U492 ( .A1(n417), .A2(KEYINPUT66), .ZN(n366) );
  INV_X1 U493 ( .A(KEYINPUT82), .ZN(n403) );
  INV_X1 U494 ( .A(G475), .ZN(n392) );
  NAND2_X1 U495 ( .A1(n367), .A2(n368), .ZN(n646) );
  NAND2_X1 U496 ( .A1(n369), .A2(n368), .ZN(n396) );
  NOR2_X1 U497 ( .A1(n375), .A2(n373), .ZN(n369) );
  NOR2_X1 U498 ( .A1(n375), .A2(n378), .ZN(n728) );
  INV_X1 U499 ( .A(n375), .ZN(n370) );
  INV_X1 U500 ( .A(G472), .ZN(n372) );
  INV_X1 U501 ( .A(n632), .ZN(n380) );
  NAND2_X2 U502 ( .A1(n734), .A2(n746), .ZN(n632) );
  XNOR2_X2 U503 ( .A(n404), .B(KEYINPUT45), .ZN(n734) );
  NAND2_X1 U504 ( .A1(n380), .A2(n363), .ZN(n377) );
  XNOR2_X2 U505 ( .A(n374), .B(G143), .ZN(n490) );
  XNOR2_X2 U506 ( .A(G128), .B(KEYINPUT65), .ZN(n374) );
  NAND2_X2 U507 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U508 ( .A1(n632), .A2(n366), .ZN(n376) );
  NOR2_X1 U509 ( .A1(n673), .A2(n662), .ZN(n596) );
  XNOR2_X1 U510 ( .A(n397), .B(n425), .ZN(n471) );
  XNOR2_X2 U511 ( .A(n468), .B(G472), .ZN(n587) );
  NAND2_X1 U512 ( .A1(n415), .A2(n413), .ZN(n412) );
  XNOR2_X1 U513 ( .A(n397), .B(n502), .ZN(n506) );
  NAND2_X1 U514 ( .A1(n587), .A2(n695), .ZN(n389) );
  INV_X1 U515 ( .A(n609), .ZN(n602) );
  NAND2_X1 U516 ( .A1(n532), .A2(n609), .ZN(n534) );
  XNOR2_X2 U517 ( .A(n587), .B(n390), .ZN(n609) );
  NOR2_X2 U518 ( .A1(n641), .A2(n733), .ZN(n642) );
  XNOR2_X1 U519 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U520 ( .A1(n518), .A2(n531), .ZN(n393) );
  XNOR2_X1 U521 ( .A(n396), .B(n637), .ZN(n641) );
  NOR2_X2 U522 ( .A1(n554), .A2(n522), .ZN(n395) );
  XNOR2_X2 U523 ( .A(n424), .B(G125), .ZN(n397) );
  XNOR2_X1 U524 ( .A(n624), .B(n623), .ZN(n405) );
  NAND2_X1 U525 ( .A1(n361), .A2(n569), .ZN(n401) );
  NAND2_X1 U526 ( .A1(n405), .A2(n357), .ZN(n404) );
  NAND2_X1 U527 ( .A1(n693), .A2(n698), .ZN(n407) );
  INV_X1 U528 ( .A(n599), .ZN(n598) );
  INV_X1 U529 ( .A(n618), .ZN(n628) );
  XNOR2_X2 U530 ( .A(n411), .B(n410), .ZN(n618) );
  NAND2_X1 U531 ( .A1(n617), .A2(n616), .ZN(n667) );
  XNOR2_X2 U532 ( .A(n614), .B(KEYINPUT32), .ZN(n652) );
  NAND2_X1 U533 ( .A1(n629), .A2(KEYINPUT66), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n416), .A2(KEYINPUT66), .ZN(n415) );
  AND2_X1 U535 ( .A1(n583), .A2(n582), .ZN(n419) );
  XNOR2_X1 U536 ( .A(KEYINPUT28), .B(KEYINPUT107), .ZN(n420) );
  XOR2_X1 U537 ( .A(KEYINPUT105), .B(n561), .Z(n421) );
  INV_X1 U538 ( .A(KEYINPUT48), .ZN(n559) );
  INV_X1 U539 ( .A(n695), .ZN(n535) );
  NOR2_X1 U540 ( .A1(n550), .A2(n535), .ZN(n536) );
  INV_X1 U541 ( .A(KEYINPUT84), .ZN(n623) );
  INV_X1 U542 ( .A(KEYINPUT19), .ZN(n520) );
  INV_X1 U543 ( .A(KEYINPUT34), .ZN(n580) );
  BUF_X1 U544 ( .A(n587), .Z(n683) );
  XNOR2_X1 U545 ( .A(n729), .B(KEYINPUT122), .ZN(n730) );
  INV_X1 U546 ( .A(KEYINPUT63), .ZN(n648) );
  XNOR2_X1 U547 ( .A(n731), .B(n730), .ZN(n732) );
  XOR2_X1 U548 ( .A(n423), .B(n422), .Z(n433) );
  INV_X1 U549 ( .A(n444), .ZN(n426) );
  NAND2_X1 U550 ( .A1(G234), .A2(n741), .ZN(n427) );
  XNOR2_X1 U551 ( .A(n428), .B(n427), .ZN(n493) );
  NAND2_X1 U552 ( .A1(G221), .A2(n493), .ZN(n431) );
  XOR2_X1 U553 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n430) );
  XNOR2_X1 U554 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n429) );
  XOR2_X1 U555 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n437) );
  XOR2_X1 U556 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n435) );
  NAND2_X1 U557 ( .A1(G234), .A2(n629), .ZN(n434) );
  XNOR2_X1 U558 ( .A(n435), .B(n434), .ZN(n438) );
  NAND2_X1 U559 ( .A1(n438), .A2(G217), .ZN(n436) );
  NAND2_X1 U560 ( .A1(n438), .A2(G221), .ZN(n440) );
  XOR2_X1 U561 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n439) );
  XNOR2_X1 U562 ( .A(n440), .B(n439), .ZN(n680) );
  AND2_X1 U563 ( .A1(n615), .A2(n680), .ZN(n592) );
  INV_X1 U564 ( .A(n592), .ZN(n676) );
  XNOR2_X1 U565 ( .A(n502), .B(G146), .ZN(n442) );
  XNOR2_X1 U566 ( .A(KEYINPUT78), .B(n444), .ZN(n446) );
  NAND2_X1 U567 ( .A1(n741), .A2(G227), .ZN(n445) );
  XNOR2_X1 U568 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U569 ( .A(n499), .B(n447), .ZN(n448) );
  XNOR2_X1 U570 ( .A(n467), .B(n448), .ZN(n720) );
  XNOR2_X1 U571 ( .A(KEYINPUT71), .B(G469), .ZN(n449) );
  INV_X1 U572 ( .A(n541), .ZN(n586) );
  NAND2_X1 U573 ( .A1(G234), .A2(G237), .ZN(n451) );
  XNOR2_X1 U574 ( .A(n451), .B(KEYINPUT14), .ZN(n707) );
  INV_X1 U575 ( .A(G952), .ZN(n638) );
  NAND2_X1 U576 ( .A1(n741), .A2(n638), .ZN(n454) );
  INV_X1 U577 ( .A(G902), .ZN(n452) );
  NAND2_X1 U578 ( .A1(G953), .A2(n452), .ZN(n453) );
  AND2_X1 U579 ( .A1(n454), .A2(n453), .ZN(n455) );
  AND2_X1 U580 ( .A1(n707), .A2(n455), .ZN(n576) );
  NAND2_X1 U581 ( .A1(G953), .A2(G900), .ZN(n456) );
  NAND2_X1 U582 ( .A1(n576), .A2(n456), .ZN(n517) );
  INV_X1 U583 ( .A(n517), .ZN(n457) );
  NAND2_X1 U584 ( .A1(n586), .A2(n457), .ZN(n458) );
  NOR2_X1 U585 ( .A1(n676), .A2(n458), .ZN(n546) );
  NAND2_X1 U586 ( .A1(n469), .A2(G210), .ZN(n460) );
  XNOR2_X1 U587 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U588 ( .A(KEYINPUT75), .B(KEYINPUT93), .ZN(n461) );
  XNOR2_X1 U589 ( .A(n462), .B(n461), .ZN(n465) );
  XNOR2_X1 U590 ( .A(n464), .B(n463), .ZN(n500) );
  XNOR2_X1 U591 ( .A(n465), .B(n500), .ZN(n466) );
  XNOR2_X1 U592 ( .A(n467), .B(n466), .ZN(n643) );
  OR2_X2 U593 ( .A1(n643), .A2(G902), .ZN(n468) );
  XNOR2_X1 U594 ( .A(KEYINPUT74), .B(n355), .ZN(n510) );
  NAND2_X1 U595 ( .A1(n510), .A2(G214), .ZN(n695) );
  NAND2_X1 U596 ( .A1(n546), .A2(n545), .ZN(n515) );
  NAND2_X1 U597 ( .A1(G214), .A2(n469), .ZN(n470) );
  XOR2_X1 U598 ( .A(G104), .B(n472), .Z(n483) );
  XNOR2_X1 U599 ( .A(n474), .B(n473), .ZN(n478) );
  XOR2_X1 U600 ( .A(G140), .B(KEYINPUT98), .Z(n476) );
  XNOR2_X1 U601 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U602 ( .A(n478), .B(n477), .ZN(n481) );
  XNOR2_X1 U603 ( .A(n479), .B(G122), .ZN(n480) );
  XNOR2_X1 U604 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U605 ( .A(n483), .B(n482), .ZN(n653) );
  NOR2_X1 U606 ( .A1(G902), .A2(n653), .ZN(n484) );
  INV_X1 U607 ( .A(KEYINPUT13), .ZN(n485) );
  XNOR2_X1 U608 ( .A(n487), .B(n486), .ZN(n492) );
  XOR2_X1 U609 ( .A(KEYINPUT7), .B(G107), .Z(n488) );
  XNOR2_X1 U610 ( .A(n488), .B(G122), .ZN(n489) );
  XNOR2_X1 U611 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U612 ( .A(n492), .B(n491), .Z(n495) );
  NAND2_X1 U613 ( .A1(G217), .A2(n493), .ZN(n494) );
  XNOR2_X1 U614 ( .A(n495), .B(n494), .ZN(n724) );
  NOR2_X1 U615 ( .A1(G902), .A2(n724), .ZN(n497) );
  XOR2_X1 U616 ( .A(KEYINPUT101), .B(G478), .Z(n496) );
  XNOR2_X1 U617 ( .A(n497), .B(n496), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n504) );
  NAND2_X1 U619 ( .A1(n741), .A2(G224), .ZN(n503) );
  XNOR2_X1 U620 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U621 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U622 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U623 ( .A(n509), .B(n740), .ZN(n636) );
  INV_X1 U624 ( .A(n629), .ZN(n631) );
  OR2_X2 U625 ( .A1(n636), .A2(n631), .ZN(n512) );
  NAND2_X1 U626 ( .A1(n510), .A2(G210), .ZN(n511) );
  XNOR2_X2 U627 ( .A(n512), .B(n511), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n553), .A2(n386), .ZN(n513) );
  NAND2_X1 U629 ( .A1(n583), .A2(n513), .ZN(n514) );
  NOR2_X1 U630 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U631 ( .A(KEYINPUT106), .B(n516), .Z(n762) );
  NAND2_X1 U632 ( .A1(n519), .A2(n586), .ZN(n554) );
  NOR2_X2 U633 ( .A1(n563), .A2(n535), .ZN(n521) );
  INV_X1 U634 ( .A(n578), .ZN(n522) );
  INV_X1 U635 ( .A(n527), .ZN(n524) );
  OR2_X1 U636 ( .A1(n583), .A2(n553), .ZN(n523) );
  XNOR2_X1 U637 ( .A(n523), .B(KEYINPUT102), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n583), .A2(n553), .ZN(n550) );
  NAND2_X1 U639 ( .A1(n566), .A2(n550), .ZN(n694) );
  NAND2_X1 U640 ( .A1(n524), .A2(n694), .ZN(n525) );
  NAND2_X1 U641 ( .A1(KEYINPUT47), .A2(n525), .ZN(n526) );
  NAND2_X1 U642 ( .A1(n762), .A2(n526), .ZN(n530) );
  NOR2_X1 U643 ( .A1(n527), .A2(n550), .ZN(n670) );
  NOR2_X1 U644 ( .A1(n668), .A2(n670), .ZN(n528) );
  NOR2_X1 U645 ( .A1(n528), .A2(KEYINPUT47), .ZN(n529) );
  NOR2_X1 U646 ( .A1(n530), .A2(n529), .ZN(n544) );
  AND2_X1 U647 ( .A1(n680), .A2(n531), .ZN(n532) );
  INV_X1 U648 ( .A(KEYINPUT104), .ZN(n533) );
  XNOR2_X1 U649 ( .A(n534), .B(n533), .ZN(n537) );
  INV_X1 U650 ( .A(n386), .ZN(n538) );
  NAND2_X1 U651 ( .A1(n561), .A2(n538), .ZN(n540) );
  XOR2_X1 U652 ( .A(KEYINPUT36), .B(KEYINPUT110), .Z(n539) );
  XNOR2_X1 U653 ( .A(n540), .B(n539), .ZN(n542) );
  AND2_X1 U654 ( .A1(n542), .A2(n384), .ZN(n543) );
  NAND2_X1 U655 ( .A1(n544), .A2(n759), .ZN(n558) );
  AND2_X1 U656 ( .A1(n545), .A2(n696), .ZN(n547) );
  INV_X1 U657 ( .A(n550), .ZN(n671) );
  NAND2_X1 U658 ( .A1(n696), .A2(n695), .ZN(n552) );
  INV_X1 U659 ( .A(n553), .ZN(n582) );
  XNOR2_X1 U660 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n555) );
  XNOR2_X1 U661 ( .A(n556), .B(n555), .ZN(n767) );
  NOR2_X2 U662 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U663 ( .A(n560), .B(n559), .ZN(n565) );
  NAND2_X1 U664 ( .A1(n421), .A2(n350), .ZN(n562) );
  XNOR2_X1 U665 ( .A(n562), .B(KEYINPUT43), .ZN(n564) );
  INV_X1 U666 ( .A(n566), .ZN(n674) );
  AND2_X1 U667 ( .A1(n567), .A2(n674), .ZN(n568) );
  XNOR2_X1 U668 ( .A(n568), .B(KEYINPUT112), .ZN(n766) );
  INV_X1 U669 ( .A(n766), .ZN(n569) );
  NOR2_X1 U670 ( .A1(n677), .A2(n676), .ZN(n570) );
  NAND2_X1 U671 ( .A1(n570), .A2(n609), .ZN(n574) );
  XNOR2_X1 U672 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n572) );
  INV_X1 U673 ( .A(KEYINPUT72), .ZN(n571) );
  XNOR2_X1 U674 ( .A(n572), .B(n571), .ZN(n573) );
  NAND2_X1 U675 ( .A1(G953), .A2(G898), .ZN(n575) );
  AND2_X1 U676 ( .A1(n576), .A2(n575), .ZN(n577) );
  INV_X1 U677 ( .A(KEYINPUT87), .ZN(n579) );
  INV_X1 U678 ( .A(n598), .ZN(n590) );
  NAND2_X1 U679 ( .A1(n592), .A2(n586), .ZN(n588) );
  NOR2_X1 U680 ( .A1(n588), .A2(n683), .ZN(n589) );
  NAND2_X1 U681 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U682 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n593) );
  INV_X1 U683 ( .A(KEYINPUT96), .ZN(n595) );
  XNOR2_X1 U684 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n597), .A2(n694), .ZN(n606) );
  XNOR2_X1 U686 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n600) );
  XNOR2_X1 U687 ( .A(n601), .B(n600), .ZN(n613) );
  AND2_X1 U688 ( .A1(n613), .A2(n350), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n617), .A2(n602), .ZN(n603) );
  XNOR2_X1 U690 ( .A(n603), .B(KEYINPUT83), .ZN(n605) );
  NAND2_X1 U691 ( .A1(n605), .A2(n604), .ZN(n660) );
  NAND2_X1 U692 ( .A1(n606), .A2(n660), .ZN(n607) );
  NOR2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n609), .B(KEYINPUT79), .ZN(n611) );
  NOR2_X1 U695 ( .A1(n677), .A2(n604), .ZN(n610) );
  AND2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n604), .A2(n683), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n618), .A2(KEYINPUT44), .ZN(n620) );
  INV_X1 U700 ( .A(KEYINPUT67), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n620), .B(n619), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n624) );
  INV_X1 U703 ( .A(n651), .ZN(n626) );
  INV_X1 U704 ( .A(KEYINPUT44), .ZN(n625) );
  AND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n627) );
  INV_X1 U706 ( .A(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U707 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n630) );
  XNOR2_X1 U708 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n634) );
  XOR2_X1 U709 ( .A(n634), .B(KEYINPUT86), .Z(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(G953), .ZN(n640) );
  INV_X1 U712 ( .A(KEYINPUT88), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n642), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U714 ( .A(n643), .Z(n644) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(G57) );
  XOR2_X1 U717 ( .A(n650), .B(G140), .Z(G42) );
  XOR2_X1 U718 ( .A(n651), .B(G122), .Z(G24) );
  XNOR2_X1 U719 ( .A(n652), .B(G119), .ZN(G21) );
  XNOR2_X1 U720 ( .A(n653), .B(KEYINPUT59), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(n657) );
  INV_X1 U722 ( .A(n733), .ZN(n656) );
  NAND2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n659) );
  INV_X1 U724 ( .A(KEYINPUT60), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n659), .B(n658), .ZN(G60) );
  XNOR2_X1 U726 ( .A(G101), .B(n660), .ZN(G3) );
  NAND2_X1 U727 ( .A1(n662), .A2(n671), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n661), .B(G104), .ZN(G6) );
  XOR2_X1 U729 ( .A(G107), .B(KEYINPUT27), .Z(n664) );
  NAND2_X1 U730 ( .A1(n662), .A2(n674), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(G9) );
  XNOR2_X1 U734 ( .A(n667), .B(G110), .ZN(G12) );
  XNOR2_X1 U735 ( .A(n668), .B(G128), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n669), .B(KEYINPUT29), .ZN(G30) );
  XOR2_X1 U737 ( .A(n670), .B(G146), .Z(G48) );
  NAND2_X1 U738 ( .A1(n673), .A2(n671), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(G113), .ZN(G15) );
  NAND2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n675), .B(G116), .ZN(G18) );
  XOR2_X1 U742 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n691) );
  NAND2_X1 U743 ( .A1(n350), .A2(n676), .ZN(n679) );
  XOR2_X1 U744 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n678) );
  XNOR2_X1 U745 ( .A(n679), .B(n678), .ZN(n687) );
  XNOR2_X1 U746 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n604), .A2(n680), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n682), .B(n681), .ZN(n685) );
  INV_X1 U749 ( .A(n683), .ZN(n684) );
  AND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U753 ( .A(n691), .B(n690), .Z(n692) );
  NOR2_X1 U754 ( .A1(n712), .A2(n692), .ZN(n705) );
  NAND2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n701) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U757 ( .A(KEYINPUT119), .B(n697), .ZN(n699) );
  NAND2_X1 U758 ( .A1(n699), .A2(n698), .ZN(n700) );
  AND2_X1 U759 ( .A1(n701), .A2(n700), .ZN(n703) );
  INV_X1 U760 ( .A(n702), .ZN(n711) );
  NOR2_X1 U761 ( .A1(n703), .A2(n711), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U763 ( .A(KEYINPUT52), .B(n706), .ZN(n709) );
  NAND2_X1 U764 ( .A1(G952), .A2(n707), .ZN(n708) );
  NOR2_X1 U765 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U766 ( .A1(G953), .A2(n710), .ZN(n716) );
  XNOR2_X1 U767 ( .A(n632), .B(KEYINPUT2), .ZN(n714) );
  NOR2_X1 U768 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U770 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U771 ( .A(KEYINPUT53), .B(n717), .Z(G75) );
  NAND2_X1 U772 ( .A1(n728), .A2(G469), .ZN(n722) );
  XOR2_X1 U773 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n718) );
  XNOR2_X1 U774 ( .A(n718), .B(KEYINPUT120), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n733), .A2(n723), .ZN(G54) );
  NAND2_X1 U778 ( .A1(n728), .A2(G478), .ZN(n726) );
  XOR2_X1 U779 ( .A(n724), .B(KEYINPUT121), .Z(n725) );
  XNOR2_X1 U780 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U781 ( .A1(n727), .A2(n733), .ZN(G63) );
  NAND2_X1 U782 ( .A1(n728), .A2(G217), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n733), .A2(n732), .ZN(G66) );
  NAND2_X1 U784 ( .A1(n734), .A2(n741), .ZN(n739) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n735) );
  XNOR2_X1 U786 ( .A(KEYINPUT61), .B(n735), .ZN(n736) );
  NAND2_X1 U787 ( .A1(n736), .A2(G898), .ZN(n737) );
  XOR2_X1 U788 ( .A(KEYINPUT123), .B(n737), .Z(n738) );
  NAND2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n745) );
  XNOR2_X1 U790 ( .A(n740), .B(G101), .ZN(n743) );
  NOR2_X1 U791 ( .A1(n741), .A2(G898), .ZN(n742) );
  NOR2_X1 U792 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n747), .B(KEYINPUT124), .ZN(n748) );
  XNOR2_X1 U795 ( .A(n749), .B(n748), .ZN(n752) );
  XOR2_X1 U796 ( .A(n746), .B(n752), .Z(n750) );
  NOR2_X1 U797 ( .A1(G953), .A2(n750), .ZN(n751) );
  XNOR2_X1 U798 ( .A(KEYINPUT125), .B(n751), .ZN(n758) );
  INV_X1 U799 ( .A(n752), .ZN(n753) );
  XNOR2_X1 U800 ( .A(G227), .B(n753), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n754), .A2(G900), .ZN(n755) );
  XNOR2_X1 U802 ( .A(KEYINPUT126), .B(n755), .ZN(n756) );
  NAND2_X1 U803 ( .A1(n756), .A2(G953), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n758), .A2(n757), .ZN(G72) );
  XNOR2_X1 U805 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n760) );
  XNOR2_X1 U806 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U807 ( .A(G125), .B(n761), .ZN(G27) );
  XNOR2_X1 U808 ( .A(G143), .B(n762), .ZN(n763) );
  XNOR2_X1 U809 ( .A(n763), .B(KEYINPUT114), .ZN(G45) );
  XOR2_X1 U810 ( .A(G131), .B(n764), .Z(n765) );
  XNOR2_X1 U811 ( .A(KEYINPUT127), .B(n765), .ZN(G33) );
  XOR2_X1 U812 ( .A(G134), .B(n766), .Z(G36) );
  XNOR2_X1 U813 ( .A(G137), .B(n767), .ZN(G39) );
endmodule

