//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT66), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT65), .Z(new_n210));
  OR3_X1    g009(.A1(new_n205), .A2(KEYINPUT69), .A3(new_n207), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT69), .B1(new_n205), .B2(new_n207), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n208), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT68), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(KEYINPUT28), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT28), .B1(new_n214), .B2(new_n216), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n204), .B(new_n213), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OR3_X1    g019(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n221), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n227));
  INV_X1    g026(.A(new_n205), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n210), .A2(new_n226), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n204), .B1(KEYINPUT67), .B2(KEYINPUT24), .ZN(new_n235));
  AND2_X1   g034(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n236));
  OAI221_X1 g035(.A(new_n225), .B1(G183gat), .B2(G190gat), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n232), .B1(new_n228), .B2(new_n229), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n234), .A2(new_n237), .A3(new_n210), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n203), .B1(new_n220), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n220), .A2(new_n240), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n241), .B1(new_n244), .B2(new_n203), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT73), .B(G197gat), .ZN(new_n246));
  INV_X1    g045(.A(G204gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT22), .ZN(new_n249));
  INV_X1    g048(.A(G211gat), .ZN(new_n250));
  INV_X1    g049(.A(G218gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G211gat), .B(G218gat), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n253), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT77), .B1(new_n245), .B2(new_n258), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n242), .A2(new_n243), .B1(G226gat), .B2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n261));
  NOR4_X1   g060(.A1(new_n260), .A2(new_n261), .A3(new_n257), .A4(new_n241), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT75), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n213), .A2(new_n204), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n219), .B1(new_n215), .B2(new_n217), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n240), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n203), .B1(new_n269), .B2(KEYINPUT29), .ZN(new_n270));
  INV_X1    g069(.A(new_n241), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n260), .A2(KEYINPUT75), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n257), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT76), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT75), .B1(new_n260), .B2(new_n241), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n270), .A2(new_n264), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(KEYINPUT76), .A3(new_n257), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n263), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  OAI21_X1  g083(.A(KEYINPUT78), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n259), .A2(new_n262), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT76), .B1(new_n279), .B2(new_n257), .ZN(new_n287));
  AOI211_X1 g086(.A(new_n275), .B(new_n258), .C1(new_n277), .C2(new_n278), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT78), .ZN(new_n290));
  INV_X1    g089(.A(new_n284), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n281), .A2(new_n294), .A3(new_n284), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n286), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT30), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G134gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n299), .B2(G127gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(KEYINPUT1), .ZN(new_n302));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  XNOR2_X1  g103(.A(G155gat), .B(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n306), .A2(KEYINPUT79), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(KEYINPUT79), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT2), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT80), .ZN(new_n311));
  XOR2_X1   g110(.A(G141gat), .B(G148gat), .Z(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(KEYINPUT80), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n307), .B(new_n308), .C1(new_n311), .C2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(G141gat), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n305), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT82), .B(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT2), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n319), .B(new_n322), .C1(new_n316), .C2(new_n312), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT4), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n315), .A2(new_n323), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n304), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(KEYINPUT3), .B2(new_n326), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT5), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n326), .B(new_n304), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT5), .B1(new_n332), .B2(new_n330), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n325), .A2(new_n328), .ZN(new_n334));
  INV_X1    g133(.A(new_n330), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT0), .ZN(new_n339));
  XNOR2_X1  g138(.A(G57gat), .B(G85gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  AOI21_X1  g140(.A(KEYINPUT6), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n331), .A2(new_n343), .A3(new_n336), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n342), .B(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n293), .A2(new_n298), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G15gat), .B(G43gat), .Z(new_n347));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n269), .A2(new_n304), .ZN(new_n350));
  INV_X1    g149(.A(new_n304), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n242), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(G227gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n349), .B1(new_n356), .B2(KEYINPUT33), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT34), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n350), .B(new_n352), .C1(KEYINPUT72), .C2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n359), .B(new_n355), .C1(new_n353), .C2(KEYINPUT72), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT32), .B1(new_n353), .B2(new_n355), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n358), .A2(KEYINPUT71), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n350), .A2(new_n352), .A3(new_n355), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n358), .A2(KEYINPUT71), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n361), .B1(new_n360), .B2(new_n365), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n357), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  INV_X1    g169(.A(new_n357), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n366), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G78gat), .B(G106gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G50gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g178(.A(new_n253), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n243), .B1(new_n380), .B2(new_n254), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n253), .A2(new_n255), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n326), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n243), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n257), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G228gat), .ZN(new_n388));
  INV_X1    g187(.A(G233gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n379), .B1(new_n257), .B2(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n326), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n392), .A2(G228gat), .A3(G233gat), .A4(new_n386), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n378), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(G22gat), .B1(new_n394), .B2(KEYINPUT84), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n394), .A2(KEYINPUT84), .A3(G22gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n390), .A2(new_n393), .ZN(new_n398));
  OAI22_X1  g197(.A1(new_n396), .A2(new_n397), .B1(new_n377), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n397), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n377), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n395), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n373), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT35), .B1(new_n346), .B2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n373), .A2(new_n399), .A3(new_n402), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n285), .A2(new_n292), .B1(new_n295), .B2(new_n297), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT35), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(new_n345), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n399), .A2(new_n402), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n293), .A2(new_n298), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n334), .A2(new_n335), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT39), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n343), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n332), .B2(new_n330), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n416), .A2(KEYINPUT85), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(KEYINPUT85), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT86), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT40), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n344), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n421), .B2(new_n420), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n411), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT87), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT37), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n281), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n426), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT87), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n279), .A2(new_n258), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n426), .B1(new_n245), .B2(new_n257), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT38), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n291), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n296), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n345), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n284), .B1(new_n427), .B2(new_n429), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n289), .A2(KEYINPUT37), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n410), .B(new_n424), .C1(new_n437), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n373), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n369), .A2(new_n372), .A3(KEYINPUT36), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n346), .B2(new_n409), .ZN(new_n447));
  AOI221_X4 g246(.A(new_n202), .B1(new_n404), .B2(new_n408), .C1(new_n442), .C2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n437), .A2(new_n441), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n424), .A2(new_n410), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n408), .A2(new_n404), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT88), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT94), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G22gat), .ZN(new_n456));
  INV_X1    g255(.A(G1gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT16), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n456), .A2(G1gat), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n459), .A2(new_n460), .A3(G8gat), .ZN(new_n461));
  INV_X1    g260(.A(G8gat), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n456), .A2(G1gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n456), .A2(new_n458), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n455), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G43gat), .B(G50gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n468));
  OR3_X1    g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT15), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT15), .B1(new_n467), .B2(new_n468), .ZN(new_n470));
  NOR2_X1   g269(.A1(G29gat), .A2(G36gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n471), .B(KEYINPUT14), .Z(new_n472));
  NAND2_X1  g271(.A1(G29gat), .A2(G36gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT92), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n469), .A2(new_n470), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n471), .B(KEYINPUT14), .ZN(new_n476));
  INV_X1    g275(.A(new_n473), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT15), .B(new_n467), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(G8gat), .B1(new_n459), .B2(new_n460), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n462), .A3(new_n464), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT94), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n466), .A2(new_n475), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n475), .A2(new_n478), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT94), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT94), .B1(new_n479), .B2(new_n480), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT13), .Z(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT95), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT95), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT18), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n461), .B2(new_n465), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT93), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT17), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n475), .A2(new_n498), .A3(new_n478), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n475), .B2(new_n478), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n496), .B(new_n497), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n488), .A3(new_n486), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n491), .A2(new_n493), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT96), .ZN(new_n504));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G169gat), .B(G197gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n501), .A2(KEYINPUT18), .A3(new_n488), .A4(new_n486), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n503), .A2(new_n504), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(new_n494), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n487), .A2(new_n492), .A3(new_n489), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n492), .B1(new_n487), .B2(new_n489), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n515), .B(new_n513), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT96), .B1(new_n518), .B2(new_n511), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n514), .A2(new_n519), .B1(new_n511), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n454), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  INV_X1    g321(.A(G71gat), .ZN(new_n523));
  INV_X1    g322(.A(G78gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT9), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n522), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(G71gat), .A2(G78gat), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT97), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n532), .A3(new_n522), .ZN(new_n533));
  AND2_X1   g332(.A1(G57gat), .A2(G64gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(G57gat), .A2(G64gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT98), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n522), .A2(new_n538), .A3(new_n527), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n522), .B2(new_n527), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n528), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G127gat), .B(G155gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT20), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n546), .B(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n466), .B(new_n481), .C1(new_n543), .C2(new_n542), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT100), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n549), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G183gat), .B(G211gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n552), .B(new_n555), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G134gat), .B(G162gat), .Z(new_n558));
  AND2_X1   g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT41), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n558), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n563), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(new_n572), .A3(new_n566), .A4(new_n570), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(KEYINPUT101), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n566), .A2(new_n570), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT101), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n578), .A2(new_n579), .A3(new_n572), .A4(new_n575), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n499), .B2(new_n500), .ZN(new_n583));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584));
  AOI22_X1  g383(.A1(new_n483), .A2(new_n581), .B1(KEYINPUT41), .B2(new_n559), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT102), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT103), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n561), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n583), .A2(new_n585), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n587), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n591), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT104), .B1(new_n557), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT104), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n597), .A3(new_n556), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n577), .A2(new_n542), .A3(new_n580), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT105), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT105), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n577), .A2(new_n542), .A3(new_n602), .A4(new_n580), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n574), .A2(new_n576), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n542), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n600), .A2(new_n601), .A3(new_n603), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT106), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n605), .B1(new_n599), .B2(KEYINPUT105), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT106), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n601), .A4(new_n603), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n582), .A2(new_n601), .A3(new_n542), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT107), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n609), .A2(new_n603), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n619), .A2(new_n621), .A3(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n521), .A2(new_n595), .A3(new_n598), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n345), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n457), .ZN(G1324gat));
  NAND2_X1  g432(.A1(new_n595), .A2(new_n598), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n634), .A2(new_n406), .A3(new_n629), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT108), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n521), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n462), .B1(new_n521), .B2(new_n635), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT42), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(KEYINPUT42), .B2(new_n638), .ZN(G1325gat));
  INV_X1    g440(.A(new_n446), .ZN(new_n642));
  OAI21_X1  g441(.A(G15gat), .B1(new_n631), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(G15gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n373), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n631), .B2(new_n645), .ZN(G1326gat));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n410), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT43), .B(G22gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  NOR3_X1   g448(.A1(new_n596), .A2(new_n556), .A3(new_n629), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n521), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT45), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n345), .A2(G29gat), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n596), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n448), .B2(new_n453), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n442), .A2(new_n447), .B1(new_n404), .B2(new_n408), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n655), .B1(new_n658), .B2(new_n596), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n556), .A2(new_n520), .A3(new_n629), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G29gat), .B1(new_n662), .B2(new_n345), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n654), .A2(new_n663), .A3(new_n664), .ZN(G1328gat));
  OR2_X1    g464(.A1(new_n406), .A2(G36gat), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n651), .A2(KEYINPUT46), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G36gat), .B1(new_n662), .B2(new_n406), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT46), .B1(new_n651), .B2(new_n666), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(G1329gat));
  NAND4_X1  g469(.A1(new_n657), .A2(new_n446), .A3(new_n659), .A4(new_n661), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G43gat), .ZN(new_n672));
  INV_X1    g471(.A(G43gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n373), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n672), .B1(new_n651), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1330gat));
  NOR2_X1   g476(.A1(new_n410), .A2(G50gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n521), .A2(new_n650), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n657), .A2(new_n409), .A3(new_n659), .A4(new_n661), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT109), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G50gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(KEYINPUT109), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT48), .B(new_n679), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT48), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n680), .A2(G50gat), .ZN(new_n686));
  INV_X1    g485(.A(new_n679), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(G1331gat));
  NAND2_X1  g488(.A1(new_n451), .A2(new_n452), .ZN(new_n690));
  INV_X1    g489(.A(new_n520), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n634), .A2(new_n691), .A3(new_n630), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n345), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g496(.A1(new_n693), .A2(new_n406), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  AND2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n698), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT110), .ZN(G1333gat));
  NAND2_X1  g502(.A1(new_n694), .A2(new_n373), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705));
  AOI21_X1  g504(.A(G71gat), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n705), .B2(new_n704), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n694), .A2(G71gat), .A3(new_n446), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT50), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(new_n711), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1334gat));
  NOR2_X1   g512(.A1(new_n693), .A2(new_n410), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(new_n524), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n691), .A2(new_n556), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n629), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n660), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n719), .A2(new_n567), .A3(new_n345), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n690), .A2(new_n594), .A3(new_n716), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n594), .A4(new_n716), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n630), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n695), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n720), .A2(new_n726), .ZN(G1336gat));
  NOR2_X1   g526(.A1(new_n406), .A2(G92gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n630), .B(new_n729), .C1(new_n723), .C2(new_n724), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(KEYINPUT52), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n657), .A2(new_n411), .A3(new_n659), .A4(new_n718), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT113), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G92gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(KEYINPUT113), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n732), .A2(new_n737), .A3(G92gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n732), .B2(G92gat), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n738), .A2(new_n739), .A3(new_n730), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n719), .B2(new_n642), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n723), .A2(new_n724), .ZN(new_n744));
  AOI211_X1 g543(.A(G99gat), .B(new_n630), .C1(new_n372), .C2(new_n369), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT114), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(G1338gat));
  NAND2_X1  g546(.A1(new_n409), .A2(G106gat), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n725), .A2(new_n409), .ZN(new_n749));
  OAI221_X1 g548(.A(KEYINPUT53), .B1(new_n719), .B2(new_n748), .C1(new_n749), .C2(G106gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n719), .A2(new_n748), .ZN(new_n752));
  AOI21_X1  g551(.A(G106gat), .B1(new_n725), .B2(new_n409), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(G1339gat));
  NAND4_X1  g554(.A1(new_n595), .A2(new_n598), .A3(new_n520), .A4(new_n630), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n615), .B2(new_n618), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n618), .B(new_n613), .C1(new_n608), .C2(new_n611), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n759), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n613), .B1(new_n608), .B2(new_n611), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n765), .A2(KEYINPUT54), .A3(new_n617), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(new_n767), .A3(new_n625), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n615), .A2(new_n760), .A3(new_n618), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n769), .B2(new_n626), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n758), .B(new_n764), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n628), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT54), .B1(new_n765), .B2(new_n617), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT55), .B1(new_n773), .B2(new_n762), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n767), .B1(new_n766), .B2(new_n625), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n769), .A2(KEYINPUT115), .A3(new_n626), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n758), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n514), .A2(new_n519), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n487), .A2(new_n489), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n488), .B1(new_n501), .B2(new_n486), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n509), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT117), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n768), .A2(new_n770), .B1(new_n762), .B2(new_n773), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n759), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n779), .A2(new_n594), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n629), .A2(new_n780), .A3(new_n784), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n520), .B1(new_n786), .B2(new_n759), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n779), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n791), .B2(new_n594), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n556), .B1(new_n792), .B2(KEYINPUT118), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n794), .B(new_n788), .C1(new_n791), .C2(new_n594), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n757), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n403), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n411), .A2(new_n345), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n691), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n629), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n556), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g604(.A1(new_n406), .A2(new_n695), .A3(new_n594), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(G134gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT56), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n299), .B1(new_n799), .B2(new_n594), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n809), .A2(new_n810), .ZN(G1343gat));
  NOR2_X1   g610(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT119), .B(new_n814), .C1(new_n796), .C2(new_n410), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n764), .B1(new_n768), .B2(new_n770), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n818));
  INV_X1    g617(.A(new_n628), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n777), .B2(new_n758), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n790), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n789), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n594), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n787), .A2(new_n594), .A3(new_n785), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n778), .A3(new_n772), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT118), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n795), .A3(new_n557), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n410), .B1(new_n827), .B2(new_n756), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n816), .B1(new_n828), .B2(KEYINPUT57), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n410), .A2(new_n814), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n792), .A2(new_n557), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n757), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n642), .A2(new_n798), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n691), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G141gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n520), .A2(G141gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n828), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n813), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n812), .B(new_n841), .C1(new_n836), .C2(G141gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n833), .A2(new_n835), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n630), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G148gat), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n756), .B(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n792), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n556), .B1(new_n792), .B2(new_n852), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n814), .B1(new_n855), .B2(new_n410), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n827), .A2(new_n756), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n830), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n834), .A2(new_n630), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n317), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n847), .A2(new_n849), .B1(new_n861), .B2(new_n848), .ZN(new_n862));
  INV_X1    g661(.A(new_n828), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n834), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n317), .A3(new_n629), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1345gat));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n320), .A3(new_n556), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n846), .A2(new_n557), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n320), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n846), .B2(new_n596), .ZN(new_n870));
  OR3_X1    g669(.A1(new_n806), .A2(G162gat), .A3(new_n446), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n863), .B2(new_n871), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n406), .A2(new_n695), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n373), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT124), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(KEYINPUT124), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(new_n409), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n857), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT125), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n880), .A3(new_n857), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(G169gat), .A3(new_n691), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n406), .A2(new_n403), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT123), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n857), .A2(new_n345), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n691), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n884), .A2(new_n888), .ZN(G1348gat));
  AND3_X1   g688(.A1(new_n883), .A2(G176gat), .A3(new_n629), .ZN(new_n890));
  AOI21_X1  g689(.A(G176gat), .B1(new_n887), .B2(new_n629), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT126), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(KEYINPUT126), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1349gat));
  OAI21_X1  g693(.A(G183gat), .B1(new_n882), .B2(new_n557), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n887), .A2(new_n215), .A3(new_n556), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n887), .A2(new_n216), .A3(new_n594), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n594), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(G190gat), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT61), .B(new_n216), .C1(new_n883), .C2(new_n594), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G1351gat));
  NAND3_X1  g703(.A1(new_n642), .A2(new_n409), .A3(new_n411), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n796), .A2(new_n695), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G197gat), .B1(new_n906), .B2(new_n691), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n642), .A2(new_n873), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n856), .B2(new_n858), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n691), .A2(G197gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(G1352gat));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n247), .A3(new_n629), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT62), .Z(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n629), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G204gat), .B1(new_n915), .B2(KEYINPUT127), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n913), .B1(new_n916), .B2(new_n918), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n906), .A2(new_n250), .A3(new_n556), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n909), .A2(new_n556), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  AOI21_X1  g723(.A(new_n251), .B1(new_n909), .B2(new_n594), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n906), .A2(new_n251), .A3(new_n594), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(new_n926), .ZN(G1355gat));
endmodule


