//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G140), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(new_n189), .B2(KEYINPUT81), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G125), .A3(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(new_n188), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n198), .B(new_n190), .C1(new_n195), .C2(new_n188), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT24), .B(G110), .Z(new_n201));
  XNOR2_X1  g015(.A(G119), .B(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT79), .B1(new_n208), .B2(G119), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT80), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n209), .B2(new_n210), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT80), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G110), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n200), .B(new_n203), .C1(new_n214), .C2(new_n218), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n213), .A2(G110), .B1(new_n202), .B2(new_n201), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT82), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n189), .A2(G140), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n191), .A2(G125), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n221), .B1(new_n228), .B2(new_n198), .ZN(new_n229));
  AOI211_X1 g043(.A(KEYINPUT83), .B(G146), .C1(new_n223), .C2(new_n227), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n197), .B(new_n220), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n219), .A2(new_n231), .A3(KEYINPUT84), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n236), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n187), .B1(new_n244), .B2(G902), .ZN(new_n245));
  INV_X1    g059(.A(G902), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n247));
  OAI211_X1 g061(.A(KEYINPUT25), .B(new_n246), .C1(new_n247), .C2(new_n238), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT78), .B(G217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n246), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n244), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(G902), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G137), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(G137), .ZN(new_n264));
  INV_X1    g078(.A(G137), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G134), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(G131), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n267), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n259), .A2(new_n257), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n264), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n269), .A2(KEYINPUT66), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(G131), .C1(new_n263), .C2(new_n268), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n198), .A2(G143), .ZN(new_n281));
  INV_X1    g095(.A(G143), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G146), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(KEYINPUT0), .B2(G128), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT0), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n208), .A3(KEYINPUT64), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n284), .A2(new_n285), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n281), .A2(new_n283), .A3(KEYINPUT0), .A4(G128), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n277), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n280), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT1), .B1(new_n282), .B2(G146), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n282), .A2(G146), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n198), .A2(G143), .ZN(new_n298));
  OAI211_X1 g112(.A(G128), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n281), .B(new_n283), .C1(KEYINPUT1), .C2(new_n208), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n266), .A2(new_n264), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G131), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n274), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G116), .B(G119), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT2), .B(G113), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n295), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n295), .A2(new_n304), .ZN(new_n311));
  INV_X1    g125(.A(new_n306), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n305), .ZN(new_n313));
  XOR2_X1   g127(.A(G116), .B(G119), .Z(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n306), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n308), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n310), .B1(new_n318), .B2(KEYINPUT28), .ZN(new_n319));
  NOR2_X1   g133(.A1(G237), .A2(G953), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G210), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT69), .Z(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G101), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n322), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G902), .B1(new_n319), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n275), .A2(new_n293), .A3(new_n277), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n304), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n333), .B2(new_n316), .ZN(new_n334));
  AOI211_X1 g148(.A(KEYINPUT72), .B(new_n307), .C1(new_n332), .C2(new_n304), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n309), .B1(new_n336), .B2(new_n308), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n337), .A2(new_n310), .A3(new_n327), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n328), .B1(new_n338), .B2(KEYINPUT75), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n316), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n333), .A2(new_n331), .A3(new_n316), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n308), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT28), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n308), .A2(new_n309), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(KEYINPUT75), .A3(new_n326), .A4(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n295), .A2(new_n304), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n295), .A2(KEYINPUT30), .A3(new_n304), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n307), .B1(new_n333), .B2(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n348), .A2(new_n307), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n347), .B1(new_n352), .B2(new_n326), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n308), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT76), .A3(new_n327), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n330), .B1(new_n339), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G472), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n308), .A2(KEYINPUT70), .A3(new_n326), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT70), .B1(new_n308), .B2(new_n326), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n354), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT71), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(new_n354), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(KEYINPUT31), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT31), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n368), .B(new_n354), .C1(new_n361), .C2(new_n362), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n327), .B1(new_n337), .B2(new_n310), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G472), .A2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(KEYINPUT32), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n360), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n359), .B1(new_n358), .B2(G472), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n373), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT74), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n373), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n367), .B2(new_n371), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT74), .B1(new_n384), .B2(new_n380), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n256), .B1(new_n377), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G214), .B1(G237), .B2(G902), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT88), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n320), .A2(G214), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n282), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n320), .A2(G143), .A3(G214), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n394), .A2(KEYINPUT17), .A3(G131), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n200), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n394), .B(G131), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(KEYINPUT17), .B2(new_n397), .ZN(new_n398));
  OAI22_X1  g212(.A1(new_n229), .A2(new_n230), .B1(new_n198), .B2(new_n195), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT18), .A2(G131), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n394), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(G104), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n398), .A2(new_n402), .A3(new_n406), .ZN(new_n409));
  AOI21_X1  g223(.A(G902), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT94), .B(G475), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n397), .A2(new_n197), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n228), .A2(KEYINPUT19), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n198), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n414), .A2(new_n417), .B1(new_n399), .B2(new_n401), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n409), .B1(new_n418), .B2(new_n406), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT20), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n413), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G478), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT15), .ZN(new_n428));
  INV_X1    g242(.A(G116), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT14), .A3(G122), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(G107), .B(new_n430), .C1(new_n434), .C2(KEYINPUT14), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n435), .A2(KEYINPUT99), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(KEYINPUT99), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT95), .ZN(new_n440));
  AOI21_X1  g254(.A(G107), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n436), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT96), .B1(new_n282), .B2(G128), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT96), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n208), .A3(G143), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n282), .A2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT98), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n449), .A2(G134), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G134), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n442), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  INV_X1    g269(.A(new_n441), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n439), .A2(new_n440), .A3(G107), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT97), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n447), .B(KEYINPUT13), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n446), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(G134), .ZN(new_n462));
  AOI211_X1 g276(.A(KEYINPUT97), .B(new_n258), .C1(new_n460), .C2(new_n446), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n455), .B(new_n458), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n250), .A2(new_n466), .A3(G953), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n454), .A2(new_n464), .A3(new_n467), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(KEYINPUT100), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(KEYINPUT100), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n428), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n428), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(G234), .A2(G237), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(G952), .A3(new_n234), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(G902), .A3(G953), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT101), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR4_X1   g298(.A1(new_n426), .A2(new_n474), .A3(new_n476), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G110), .B(G122), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT3), .B1(new_n405), .B2(G107), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT3), .ZN(new_n489));
  INV_X1    g303(.A(G107), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(G104), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n405), .A2(G107), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(G101), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(new_n307), .ZN(new_n497));
  INV_X1    g311(.A(G101), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n488), .A2(new_n491), .A3(new_n498), .A4(new_n492), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(G101), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT86), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND4_X1   g316(.A1(KEYINPUT86), .A2(new_n501), .A3(KEYINPUT4), .A4(new_n499), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT89), .B(new_n497), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n405), .A2(G107), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n490), .A2(G104), .ZN(new_n506));
  OAI21_X1  g320(.A(G101), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n205), .A3(G116), .ZN(new_n510));
  OAI211_X1 g324(.A(G113), .B(new_n510), .C1(new_n314), .C2(new_n509), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n313), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n316), .A2(new_n495), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n501), .A2(KEYINPUT4), .A3(new_n499), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n500), .A2(KEYINPUT86), .A3(new_n501), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT89), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n487), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n524), .A2(new_n486), .A3(new_n512), .A4(new_n504), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(KEYINPUT6), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n487), .C1(new_n513), .C2(new_n520), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n292), .A2(G125), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n299), .A2(new_n300), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n189), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G224), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n532), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n526), .A2(new_n528), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n511), .A2(new_n313), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n499), .A2(new_n507), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT91), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n486), .B(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n539), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n512), .ZN(new_n546));
  INV_X1    g360(.A(new_n534), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n532), .A2(KEYINPUT7), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n529), .A2(new_n531), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n543), .A2(new_n546), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n525), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n537), .B1(new_n552), .B2(new_n246), .ZN(new_n553));
  AOI211_X1 g367(.A(KEYINPUT92), .B(G902), .C1(new_n525), .C2(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n536), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G210), .B1(G237), .B2(G902), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT93), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n536), .B(new_n556), .C1(new_n553), .C2(new_n554), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n555), .A2(new_n561), .A3(new_n557), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G469), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n530), .A2(new_n539), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n299), .A2(new_n499), .A3(new_n507), .A4(new_n300), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n280), .A2(new_n294), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n278), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n568), .A2(new_n569), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT87), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n301), .A2(new_n508), .A3(new_n572), .A4(KEYINPUT10), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(KEYINPUT10), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n572), .A2(KEYINPUT10), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n566), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n496), .A2(new_n292), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n502), .B2(new_n503), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n277), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT67), .B1(new_n275), .B2(new_n277), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G140), .ZN(new_n585));
  INV_X1    g399(.A(G227), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G953), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n585), .B(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n571), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n573), .A2(new_n576), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n517), .A2(new_n518), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n280), .A2(new_n294), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n580), .A2(new_n583), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n564), .B(new_n246), .C1(new_n589), .C2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n588), .B1(new_n571), .B2(new_n584), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(new_n590), .A3(new_n596), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(G469), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(G469), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G221), .B1(new_n466), .B2(G902), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT85), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  AND4_X1   g421(.A1(new_n390), .A2(new_n485), .A3(new_n563), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n387), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  NAND2_X1  g424(.A1(new_n372), .A2(new_n246), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  INV_X1    g426(.A(new_n256), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n612), .A2(new_n378), .A3(new_n613), .A4(new_n607), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n389), .B1(new_n558), .B2(new_n560), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n427), .A2(new_n246), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n471), .B2(new_n427), .ZN(new_n617));
  INV_X1    g431(.A(new_n470), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n467), .B1(new_n454), .B2(new_n464), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n469), .A2(new_n621), .A3(new_n470), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n622), .A3(G478), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n425), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n483), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n615), .A2(KEYINPUT102), .A3(new_n483), .A4(new_n625), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n614), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n615), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n425), .B1(new_n474), .B2(new_n476), .ZN(new_n634));
  NOR4_X1   g448(.A1(new_n614), .A2(new_n484), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NAND3_X1  g451(.A1(new_n612), .A2(new_n378), .A3(new_n607), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n243), .A2(KEYINPUT36), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT103), .Z(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n242), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n240), .A3(new_n241), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n254), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n252), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n485), .A2(new_n563), .A3(new_n390), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n638), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT37), .B(G110), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  NAND2_X1  g464(.A1(new_n358), .A2(G472), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT77), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n360), .A2(new_n374), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n386), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n607), .A2(new_n646), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n481), .A2(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n478), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n425), .B(new_n657), .C1(new_n474), .C2(new_n476), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n655), .A2(new_n633), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n563), .B(KEYINPUT38), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n657), .B(KEYINPUT39), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n607), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n666));
  INV_X1    g480(.A(new_n646), .ZN(new_n667));
  INV_X1    g481(.A(new_n428), .ZN(new_n668));
  INV_X1    g482(.A(new_n473), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n471), .A2(KEYINPUT100), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n425), .B1(new_n671), .B2(new_n475), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n390), .A3(new_n672), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n662), .A2(new_n665), .A3(new_n666), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n318), .A2(new_n327), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n364), .A2(new_n366), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n675), .B1(new_n677), .B2(new_n246), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(KEYINPUT32), .B2(new_n384), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n379), .B1(new_n378), .B2(new_n381), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n380), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NAND2_X1  g498(.A1(new_n625), .A2(new_n657), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n655), .A2(new_n633), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n654), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  OAI21_X1  g502(.A(new_n246), .B1(new_n589), .B2(new_n597), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G469), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n690), .A2(new_n606), .A3(new_n598), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n628), .B2(new_n629), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n654), .A2(new_n613), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR4_X1   g510(.A1(new_n633), .A2(new_n692), .A3(new_n634), .A4(new_n484), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n654), .A2(new_n613), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  AND4_X1   g513(.A1(new_n485), .A2(new_n615), .A3(new_n646), .A4(new_n691), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n654), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n319), .A2(new_n326), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n367), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n369), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n703), .B1(new_n367), .B2(new_n704), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n373), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n256), .B(new_n709), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n483), .A2(new_n615), .A3(new_n672), .A4(new_n691), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n710), .A3(new_n711), .A4(new_n612), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n675), .B1(new_n372), .B2(new_n246), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n367), .A2(new_n704), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT104), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n369), .A3(new_n705), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n715), .B1(new_n718), .B2(new_n373), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(KEYINPUT106), .A3(new_n710), .A4(new_n711), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NAND2_X1  g536(.A1(new_n615), .A2(new_n691), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n685), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n612), .A2(new_n708), .A3(new_n646), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT107), .B(G125), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G27));
  AOI211_X1 g541(.A(KEYINPUT42), .B(new_n256), .C1(new_n377), .C2(new_n386), .ZN(new_n728));
  INV_X1    g542(.A(new_n685), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n560), .A2(new_n390), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n559), .A2(new_n730), .A3(new_n562), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n601), .A2(KEYINPUT108), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n599), .A2(new_n600), .A3(new_n734), .A4(G469), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n598), .A3(new_n602), .A4(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(KEYINPUT109), .A3(new_n606), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT109), .B1(new_n736), .B2(new_n606), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n559), .A2(new_n730), .A3(new_n740), .A4(new_n562), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n729), .A2(new_n732), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n384), .A2(KEYINPUT32), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n652), .A3(new_n374), .A4(new_n360), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n710), .A3(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n728), .A2(new_n742), .B1(new_n745), .B2(KEYINPUT42), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  INV_X1    g561(.A(new_n658), .ZN(new_n748));
  AND4_X1   g562(.A1(new_n748), .A2(new_n732), .A3(new_n739), .A4(new_n741), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n654), .A2(new_n749), .A3(new_n613), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND2_X1  g565(.A1(new_n599), .A2(new_n600), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n599), .A2(KEYINPUT45), .A3(new_n600), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(new_n602), .ZN(new_n757));
  OR3_X1    g571(.A1(new_n757), .A2(KEYINPUT111), .A3(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT111), .B1(new_n757), .B2(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(new_n598), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n606), .ZN(new_n762));
  INV_X1    g576(.A(new_n663), .ZN(new_n763));
  OR3_X1    g577(.A1(new_n762), .A2(KEYINPUT112), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT112), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n732), .A2(new_n741), .ZN(new_n766));
  INV_X1    g580(.A(new_n624), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n425), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT43), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n667), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n612), .A2(new_n378), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n766), .B1(new_n773), .B2(KEYINPUT44), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n764), .A2(new_n765), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT113), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n265), .ZN(G39));
  XNOR2_X1  g594(.A(new_n762), .B(KEYINPUT47), .ZN(new_n781));
  OR4_X1    g595(.A1(new_n654), .A2(new_n613), .A3(new_n685), .A4(new_n766), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n191), .ZN(G42));
  INV_X1    g598(.A(new_n682), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n768), .A2(new_n389), .A3(new_n605), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n690), .A2(new_n598), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n710), .A2(new_n786), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n785), .A2(new_n791), .A3(new_n662), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n744), .A2(new_n710), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n769), .A2(new_n478), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n766), .A2(new_n692), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(G952), .A3(new_n234), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n256), .A2(new_n478), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n785), .A2(new_n796), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n625), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n719), .A2(new_n710), .A3(new_n795), .ZN(new_n805));
  OAI221_X1 g619(.A(new_n804), .B1(new_n723), .B2(new_n805), .C1(new_n797), .C2(new_n799), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n788), .A2(new_n606), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n781), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n805), .A2(new_n766), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(KEYINPUT51), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n662), .A2(new_n389), .A3(new_n691), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n805), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT50), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n646), .A2(new_n796), .A3(new_n719), .A4(new_n795), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n426), .A2(new_n767), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n803), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n801), .B(new_n806), .C1(new_n812), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n809), .A2(new_n822), .A3(new_n810), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n815), .A2(KEYINPUT117), .A3(new_n818), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT117), .B1(new_n815), .B2(new_n818), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n820), .B1(new_n827), .B2(KEYINPUT51), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n742), .A2(new_n646), .A3(new_n719), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n607), .A2(new_n646), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n425), .A2(new_n657), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n474), .A3(new_n476), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n832), .A2(new_n732), .A3(new_n741), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n654), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n750), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n625), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n484), .B1(new_n838), .B2(new_n634), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n563), .A3(new_n390), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n614), .A2(new_n840), .B1(new_n638), .B2(new_n647), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n387), .B2(new_n608), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n615), .A2(new_n672), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n252), .A2(new_n645), .A3(new_n657), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n736), .A2(new_n606), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n251), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n245), .B2(new_n248), .ZN(new_n848));
  INV_X1    g662(.A(new_n645), .ZN(new_n849));
  INV_X1    g663(.A(new_n657), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n606), .A4(new_n736), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n843), .A2(new_n846), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(new_n682), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n680), .A2(new_n681), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n652), .A2(new_n374), .A3(new_n360), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n856), .A2(new_n857), .B1(new_n659), .B2(new_n686), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n719), .A2(new_n646), .A3(new_n724), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n746), .A2(new_n837), .A3(new_n842), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n694), .A2(new_n698), .A3(new_n701), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n682), .A2(new_n854), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT52), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n865), .A3(new_n721), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n830), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n387), .A2(new_n749), .B1(new_n654), .B2(new_n835), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n842), .A2(new_n868), .A3(new_n831), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n732), .A2(new_n739), .A3(new_n729), .A4(new_n741), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT42), .B1(new_n793), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT42), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n387), .A2(new_n872), .A3(new_n742), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n860), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n832), .A2(new_n615), .A3(new_n748), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n832), .A2(new_n615), .A3(new_n729), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n377), .A2(new_n386), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n725), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n876), .B1(new_n880), .B2(new_n863), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n721), .A2(new_n694), .A3(new_n698), .A4(new_n701), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n883), .A3(KEYINPUT53), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n867), .A2(new_n884), .A3(KEYINPUT54), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n867), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n829), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n861), .A2(new_n866), .A3(new_n830), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n875), .B2(new_n883), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n867), .A2(new_n884), .A3(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT115), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n828), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(G952), .A2(G953), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n792), .B1(new_n894), .B2(new_n895), .ZN(G75));
  OR2_X1    g710(.A1(new_n234), .A2(G952), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT120), .Z(new_n898));
  AOI21_X1  g712(.A(new_n246), .B1(new_n867), .B2(new_n884), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(G210), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n526), .A2(new_n528), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n535), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n898), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n899), .A2(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(KEYINPUT119), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n557), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n907), .B2(new_n909), .ZN(G51));
  INV_X1    g724(.A(new_n898), .ZN(new_n911));
  INV_X1    g725(.A(new_n756), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n912), .A3(new_n906), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n602), .B(KEYINPUT57), .Z(new_n914));
  NAND3_X1  g728(.A1(new_n891), .A2(new_n892), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n597), .B2(new_n589), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n911), .B1(new_n913), .B2(new_n916), .ZN(G54));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n905), .A2(new_n906), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n419), .ZN(new_n920));
  INV_X1    g734(.A(new_n419), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n905), .A2(new_n921), .A3(new_n906), .A4(new_n918), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n911), .B1(new_n920), .B2(new_n922), .ZN(G60));
  XNOR2_X1  g737(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(new_n616), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n887), .A2(new_n893), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n620), .A2(new_n622), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n891), .A2(new_n928), .A3(new_n892), .A4(new_n926), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n898), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n934), .A3(new_n898), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n930), .A2(new_n933), .A3(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(new_n867), .A2(new_n884), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT124), .ZN(new_n939));
  XNOR2_X1  g753(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n244), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n937), .A2(new_n644), .A3(new_n941), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n898), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G66));
  OAI21_X1  g761(.A(G953), .B1(new_n479), .B2(new_n533), .ZN(new_n948));
  INV_X1    g762(.A(new_n842), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n882), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n950), .B2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n901), .B1(G898), .B2(new_n234), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  NAND2_X1  g767(.A1(new_n683), .A2(new_n880), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  AOI211_X1 g769(.A(new_n664), .B(new_n766), .C1(new_n838), .C2(new_n634), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n387), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n779), .A2(new_n783), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(G953), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n333), .A2(new_n350), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n349), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n415), .A2(new_n416), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n783), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n764), .A2(new_n843), .A3(new_n765), .A4(new_n794), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n750), .A3(new_n880), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n746), .B1(new_n775), .B2(new_n778), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(G953), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(G900), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n963), .B1(new_n969), .B2(new_n234), .ZN(new_n970));
  OAI22_X1  g784(.A1(new_n959), .A2(new_n963), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(G953), .B1(new_n586), .B2(new_n969), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n974), .B(new_n976), .ZN(G72));
  XNOR2_X1  g791(.A(new_n355), .B(KEYINPUT127), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n955), .A2(new_n950), .A3(new_n958), .ZN(new_n980));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT63), .Z(new_n982));
  AOI211_X1 g796(.A(new_n327), .B(new_n979), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n982), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n966), .A2(new_n967), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n950), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n979), .A2(new_n327), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n898), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n364), .A2(new_n366), .A3(new_n353), .A4(new_n356), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n937), .A2(new_n982), .A3(new_n989), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n983), .A2(new_n988), .A3(new_n990), .ZN(G57));
endmodule


