//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n208), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n206), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(G50), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n212), .B1(KEYINPUT1), .B2(new_n219), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n238), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n239), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n220), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n206), .A2(G1), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G50), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n206), .B1(new_n201), .B2(new_n239), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT67), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n206), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n251), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n249), .B(new_n255), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G223), .A3(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G77), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n269), .B(new_n270), .C1(new_n271), .C2(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  AND2_X1   g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n220), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(KEYINPUT66), .A3(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(G274), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G226), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n266), .B1(new_n290), .B2(G169), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(G179), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n264), .A2(new_n265), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n255), .A2(new_n249), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n296), .A2(KEYINPUT9), .B1(new_n289), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n266), .A2(new_n299), .B1(new_n290), .B2(new_n300), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n298), .A2(KEYINPUT10), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n298), .B2(new_n301), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n293), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n259), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT15), .B(G87), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n261), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n265), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n247), .A2(KEYINPUT69), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT69), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n311), .A2(new_n205), .A3(G13), .A4(G20), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n251), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n313), .A2(G77), .A3(new_n254), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n312), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(G77), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n309), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n275), .A2(new_n278), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G107), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n319), .A2(new_n320), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n318), .B1(new_n327), .B2(KEYINPUT68), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT68), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n319), .A2(new_n320), .A3(new_n329), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G244), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n284), .A2(new_n286), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n285), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n317), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n334), .B1(new_n328), .B2(new_n330), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n339), .A2(KEYINPUT70), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT70), .B1(new_n339), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n317), .C1(new_n300), .C2(new_n339), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n304), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n322), .A2(new_n324), .A3(G226), .A4(new_n268), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n322), .A2(new_n324), .A3(G232), .A4(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n279), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n284), .A2(G238), .A3(new_n286), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n285), .A2(new_n352), .A3(KEYINPUT71), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT71), .B1(new_n285), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT13), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n351), .B(new_n358), .C1(new_n354), .C2(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G200), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(KEYINPUT72), .ZN(new_n362));
  INV_X1    g0162(.A(new_n355), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n353), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n358), .A4(new_n351), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n362), .A2(new_n366), .A3(new_n357), .A4(G190), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n241), .A2(G20), .ZN(new_n368));
  INV_X1    g0168(.A(new_n262), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n368), .B1(new_n260), .B2(new_n271), .C1(new_n369), .C2(new_n239), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n251), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT11), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT11), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n373), .A3(new_n251), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n313), .A2(G68), .A3(new_n254), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n310), .A2(new_n312), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n241), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n378), .A2(KEYINPUT12), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n205), .A2(G13), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n380), .A2(new_n368), .A3(KEYINPUT12), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n375), .B(new_n376), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n361), .A2(new_n367), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT73), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n361), .A2(new_n367), .A3(new_n383), .A4(KEYINPUT73), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n360), .A2(G169), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT14), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n362), .A2(new_n366), .A3(new_n357), .A4(G179), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n360), .A2(new_n392), .A3(G169), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n382), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n325), .B2(new_n206), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n398), .B(G20), .C1(new_n322), .C2(new_n324), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G58), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n241), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n201), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n262), .A2(G159), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n398), .B1(new_n267), .B2(G20), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n241), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n408), .B1(new_n411), .B2(new_n405), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(new_n412), .A3(new_n251), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n258), .A2(new_n253), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n252), .B1(new_n248), .B2(new_n258), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n284), .A2(G232), .A3(new_n286), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n285), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n322), .A2(new_n324), .A3(G223), .A4(new_n268), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n322), .A2(new_n324), .A3(G226), .A4(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G87), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n321), .C2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n422), .B2(new_n279), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G169), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n418), .A2(KEYINPUT74), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n285), .A2(new_n417), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(G179), .B1(new_n422), .B2(new_n279), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n416), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n416), .B2(new_n430), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n422), .A2(new_n279), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n297), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n425), .A2(new_n427), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n436), .A2(new_n437), .B1(new_n423), .B2(G200), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n413), .A3(new_n415), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n438), .A2(new_n413), .A3(KEYINPUT17), .A4(new_n415), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n346), .A2(new_n396), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n322), .A2(new_n324), .A3(G244), .A4(new_n268), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT4), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G250), .A2(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT4), .A2(G244), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G1698), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n267), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n279), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n282), .A2(G1), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G257), .A3(new_n284), .ZN(new_n462));
  INV_X1    g0262(.A(G274), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n276), .B2(new_n277), .ZN(new_n464));
  OR2_X1    g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n458), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n466), .A3(new_n457), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n456), .A2(new_n468), .A3(new_n340), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n318), .B1(new_n448), .B2(new_n454), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n462), .A2(new_n467), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n337), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n369), .A2(new_n271), .ZN(new_n474));
  XNOR2_X1  g0274(.A(G97), .B(G107), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n476), .A2(new_n478), .A3(G107), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n474), .B1(new_n481), .B2(G20), .ZN(new_n482));
  OAI21_X1  g0282(.A(G107), .B1(new_n397), .B2(new_n399), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(new_n251), .B1(new_n478), .B2(new_n248), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n205), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n247), .A2(new_n486), .A3(new_n220), .A4(new_n250), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G97), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n473), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT76), .ZN(new_n491));
  AOI21_X1  g0291(.A(G200), .B1(new_n456), .B2(new_n468), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n470), .A2(new_n471), .A3(G190), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n474), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n479), .B1(new_n475), .B2(new_n476), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n206), .ZN(new_n497));
  INV_X1    g0297(.A(G107), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n409), .B2(new_n410), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n251), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n248), .A2(new_n478), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n489), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n491), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n456), .A2(new_n468), .A3(new_n297), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n470), .A2(new_n471), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(G200), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n485), .A3(KEYINPUT76), .A4(new_n489), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n490), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT77), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n507), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n472), .A3(new_n469), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT77), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n322), .A2(new_n324), .A3(new_n206), .A4(G87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT22), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n267), .A2(new_n517), .A3(new_n206), .A4(G87), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT23), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n206), .B2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n498), .A2(KEYINPUT23), .A3(G20), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n321), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n521), .A2(new_n522), .B1(new_n524), .B2(new_n206), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT24), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n519), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n265), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n488), .A2(G107), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n248), .B(new_n498), .C1(KEYINPUT81), .C2(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n461), .A2(G264), .A3(new_n284), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G250), .A2(G1698), .ZN(new_n538));
  INV_X1    g0338(.A(G257), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(G1698), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n267), .B1(G33), .B2(G294), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n467), .B(new_n537), .C1(new_n541), .C2(new_n318), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT82), .B1(new_n543), .B2(G200), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n545), .A3(new_n300), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n542), .A2(G190), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n536), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n206), .B1(new_n349), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n421), .A2(new_n478), .A3(new_n498), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n322), .A2(new_n324), .A3(new_n206), .A4(G68), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n550), .B1(new_n260), .B2(new_n478), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n251), .B1(new_n377), .B2(new_n306), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n487), .A2(KEYINPUT75), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n487), .A2(KEYINPUT75), .ZN(new_n559));
  OAI21_X1  g0359(.A(G87), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G250), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n205), .B2(G45), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n464), .A2(new_n457), .B1(new_n284), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G238), .A2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n332), .B2(G1698), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n524), .B1(new_n566), .B2(new_n267), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n297), .C1(new_n567), .C2(new_n318), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n564), .B1(new_n567), .B2(new_n318), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n300), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n561), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(G169), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n564), .B(G179), .C1(new_n567), .C2(new_n318), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n307), .B1(new_n558), .B2(new_n559), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n572), .A2(new_n573), .B1(new_n557), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT78), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n284), .A2(G274), .A3(new_n457), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n563), .A2(new_n284), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n332), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G238), .B2(G1698), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n581), .A2(new_n325), .B1(new_n321), .B2(new_n523), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n279), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n573), .B1(new_n583), .B2(new_n337), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n557), .A2(new_n574), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT78), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n570), .A2(new_n568), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n561), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n542), .A2(new_n337), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n539), .A2(G1698), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(G250), .B2(G1698), .ZN(new_n592));
  INV_X1    g0392(.A(G294), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n592), .A2(new_n325), .B1(new_n321), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n279), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n595), .A2(new_n340), .A3(new_n467), .A4(new_n537), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n530), .B2(new_n535), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n549), .A2(new_n576), .A3(new_n589), .A4(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n315), .A2(G116), .A3(new_n265), .A4(new_n486), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n310), .A2(new_n523), .A3(new_n312), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n250), .A2(new_n220), .B1(G20), .B2(new_n523), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n449), .B(new_n206), .C1(G33), .C2(new_n478), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT20), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n600), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT79), .ZN(new_n607));
  INV_X1    g0407(.A(G303), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n325), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n268), .A2(G264), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G257), .A2(G1698), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n322), .B(new_n324), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n607), .B1(new_n613), .B2(new_n318), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n279), .A2(KEYINPUT79), .A3(new_n609), .A4(new_n612), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n461), .A2(G270), .A3(new_n284), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n467), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n606), .B1(new_n620), .B2(G200), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n297), .B2(new_n620), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n467), .A3(G179), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n616), .A2(new_n606), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT80), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n614), .B2(new_n615), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT80), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n606), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT21), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n620), .A2(new_n631), .A3(G169), .A4(new_n606), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n606), .A2(G169), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n618), .B1(new_n614), .B2(new_n615), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT21), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n622), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n599), .A2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n445), .A2(new_n509), .A3(new_n514), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n388), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n395), .B1(new_n640), .B2(new_n343), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n443), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n434), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n302), .A2(new_n303), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n293), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n636), .A2(new_n630), .A3(new_n598), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n584), .A2(KEYINPUT83), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT83), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n572), .A2(new_n648), .A3(new_n573), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n571), .B1(new_n650), .B2(new_n585), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n508), .A2(new_n646), .A3(new_n549), .A4(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n585), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n647), .B2(new_n649), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n654), .A2(new_n511), .A3(new_n571), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n576), .A2(new_n490), .A3(new_n589), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT26), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n652), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n445), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n645), .A2(new_n661), .ZN(G369));
  NAND2_X1  g0462(.A1(new_n636), .A2(new_n630), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  OAI21_X1  g0466(.A(G213), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G343), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n663), .A2(new_n606), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n606), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n622), .A2(new_n630), .A3(new_n636), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n549), .B(new_n598), .C1(new_n536), .C2(new_n669), .ZN(new_n677));
  INV_X1    g0477(.A(new_n598), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n670), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n670), .B1(new_n636), .B2(new_n630), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n549), .A3(new_n598), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n669), .B(KEYINPUT86), .Z(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n209), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n552), .A2(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n223), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n537), .B1(new_n541), .B2(new_n318), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n569), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n627), .A2(new_n505), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT88), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n505), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n583), .A2(G179), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n620), .A2(new_n704), .A3(new_n542), .A4(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n627), .A2(new_n698), .A3(KEYINPUT30), .A4(new_n505), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n703), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n696), .B1(new_n710), .B2(new_n669), .ZN(new_n711));
  INV_X1    g0511(.A(new_n684), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n699), .A2(new_n701), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n707), .A3(new_n706), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT87), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n712), .A2(KEYINPUT87), .A3(KEYINPUT31), .A4(new_n714), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n711), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n638), .A2(new_n514), .A3(new_n509), .A4(new_n684), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n695), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n660), .A2(new_n684), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n510), .A2(new_n651), .A3(new_n511), .A4(new_n549), .ZN(new_n725));
  INV_X1    g0525(.A(new_n646), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT90), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n654), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n651), .A2(new_n549), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT90), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n730), .A3(new_n508), .A4(new_n646), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n658), .A2(KEYINPUT89), .A3(new_n656), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n655), .A2(KEYINPUT26), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT89), .B1(new_n658), .B2(new_n656), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT29), .B(new_n669), .C1(new_n732), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n721), .B1(new_n724), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n694), .B1(new_n739), .B2(G1), .ZN(G364));
  INV_X1    g0540(.A(new_n676), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n206), .A2(G13), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n205), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n689), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n741), .B(new_n747), .C1(G330), .C2(new_n674), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n688), .A2(new_n325), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n749), .A2(G355), .B1(new_n523), .B2(new_n688), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n209), .A2(new_n325), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT91), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G45), .B2(new_n223), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n245), .A2(new_n282), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT92), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n220), .B1(G20), .B2(new_n337), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n747), .B1(new_n755), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  INV_X1    g0564(.A(new_n761), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n206), .A2(new_n340), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n767), .A2(new_n297), .A3(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G322), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n769), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n206), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n771), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n267), .B(new_n774), .C1(G329), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n766), .A2(new_n297), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G317), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n206), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n787), .A2(G294), .B1(new_n789), .B2(G303), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n775), .A2(new_n297), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G326), .A2(new_n792), .B1(new_n794), .B2(G283), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n778), .A2(new_n784), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT94), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT32), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n777), .B2(G159), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(G97), .C2(new_n787), .ZN(new_n803));
  INV_X1    g0603(.A(new_n768), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n267), .B1(new_n271), .B2(new_n773), .C1(new_n804), .C2(new_n401), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n791), .A2(new_n239), .B1(new_n788), .B2(new_n421), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n779), .A2(new_n241), .B1(new_n793), .B2(new_n498), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n796), .A2(new_n797), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n798), .A2(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n764), .B1(new_n765), .B2(new_n810), .C1(new_n674), .C2(new_n759), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n748), .A2(new_n811), .ZN(G396));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  INV_X1    g0613(.A(G150), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n791), .B1(new_n779), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT96), .Z(new_n816));
  INV_X1    g0616(.A(G143), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n817), .B2(new_n804), .C1(new_n799), .C2(new_n773), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n793), .A2(new_n241), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n267), .B1(new_n776), .B2(new_n823), .C1(new_n239), .C2(new_n788), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(G58), .C2(new_n787), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n820), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n804), .A2(new_n593), .B1(new_n478), .B2(new_n786), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT95), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n325), .B1(new_n776), .B2(new_n770), .C1(new_n773), .C2(new_n523), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n791), .A2(new_n608), .B1(new_n793), .B2(new_n421), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n779), .A2(new_n831), .B1(new_n788), .B2(new_n498), .ZN(new_n832));
  OR3_X1    g0632(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n826), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n761), .A2(new_n756), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n834), .A2(new_n761), .B1(new_n271), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n317), .A2(new_n669), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n343), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n343), .B(new_n345), .C1(new_n317), .C2(new_n669), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n836), .B1(new_n757), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n746), .ZN(new_n842));
  INV_X1    g0642(.A(new_n840), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n722), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n660), .A2(new_n684), .A3(new_n840), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT98), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n721), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n720), .A2(new_n711), .A3(new_n717), .A4(new_n718), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(G330), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n850), .A2(KEYINPUT98), .A3(new_n844), .A4(new_n845), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n848), .A2(new_n851), .B1(new_n847), .B2(new_n846), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n842), .B1(new_n852), .B2(new_n746), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT99), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n842), .B(new_n855), .C1(new_n746), .C2(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NAND2_X1  g0658(.A1(new_n416), .A2(new_n430), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT100), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n415), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n400), .A2(new_n406), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n265), .B1(new_n865), .B2(new_n408), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n866), .B2(new_n407), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n867), .B2(new_n438), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n416), .A2(new_n668), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n416), .A2(new_n430), .A3(KEYINPUT100), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n861), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n859), .A2(new_n869), .A3(new_n439), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n869), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n428), .A2(new_n429), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(G169), .B2(new_n423), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT18), .B1(new_n867), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n416), .A2(new_n430), .A3(new_n431), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n441), .A2(new_n442), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n874), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n874), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n382), .A2(new_n670), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n396), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n388), .A2(new_n395), .A3(new_n887), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n843), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n710), .A2(new_n669), .B1(KEYINPUT103), .B2(KEYINPUT31), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(new_n702), .A3(new_n707), .A4(new_n706), .ZN(new_n894));
  NOR2_X1   g0694(.A1(KEYINPUT103), .A2(KEYINPUT31), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n670), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n720), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n886), .A2(new_n891), .A3(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n889), .A2(new_n890), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n901), .A2(new_n898), .A3(new_n840), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n867), .A2(new_n877), .A3(new_n860), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT100), .B1(new_n416), .B2(new_n430), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n869), .A2(new_n439), .A3(new_n862), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n907), .A2(new_n908), .B1(new_n872), .B2(new_n863), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n869), .B1(new_n434), .B2(new_n443), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n903), .B1(new_n911), .B2(new_n885), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n899), .A2(new_n900), .B1(new_n902), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n445), .A2(new_n898), .ZN(new_n915));
  OAI21_X1  g0715(.A(G330), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n914), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT104), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n872), .A2(new_n863), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n871), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n923), .B2(new_n882), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n394), .A2(new_n382), .A3(new_n669), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n925), .B(new_n927), .C1(new_n886), .C2(new_n920), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n343), .A2(new_n670), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n845), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n886), .A2(new_n930), .A3(new_n901), .ZN(new_n931));
  INV_X1    g0731(.A(new_n668), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n880), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n928), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n445), .A2(new_n738), .A3(new_n724), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n645), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n919), .A2(new_n937), .B1(G1), .B2(new_n742), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n919), .B2(new_n937), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n523), .B(new_n222), .C1(new_n481), .C2(KEYINPUT35), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(KEYINPUT35), .B2(new_n481), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT36), .Z(new_n942));
  OR3_X1    g0742(.A1(new_n223), .A2(new_n271), .A3(new_n402), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n205), .B(G13), .C1(new_n943), .C2(new_n240), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n939), .A2(new_n945), .ZN(G367));
  INV_X1    g0746(.A(new_n752), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n762), .B1(new_n209), .B2(new_n306), .C1(new_n947), .C2(new_n234), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n746), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n804), .A2(new_n608), .B1(new_n791), .B2(new_n770), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT111), .ZN(new_n951));
  XOR2_X1   g0751(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n788), .B2(new_n523), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n950), .A2(KEYINPUT109), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n953), .A2(new_n951), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(KEYINPUT109), .C2(new_n950), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n325), .B1(new_n776), .B2(new_n781), .C1(new_n773), .C2(new_n831), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n788), .A2(new_n523), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(KEYINPUT46), .B2(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G294), .A2(new_n780), .B1(new_n794), .B2(G97), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n498), .C2(new_n786), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n786), .A2(new_n241), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G150), .B2(new_n768), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT112), .Z(new_n964));
  OAI221_X1 g0764(.A(new_n267), .B1(new_n776), .B2(new_n813), .C1(new_n773), .C2(new_n239), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n779), .A2(new_n799), .B1(new_n788), .B2(new_n401), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n791), .A2(new_n817), .B1(new_n793), .B2(new_n271), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n956), .A2(new_n961), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n949), .B1(new_n970), .B2(new_n761), .ZN(new_n971));
  INV_X1    g0771(.A(new_n561), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n651), .B1(new_n972), .B2(new_n669), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n654), .A2(new_n561), .A3(new_n670), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n973), .A2(new_n760), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n712), .A2(new_n502), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n508), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n511), .B1(new_n978), .B2(new_n598), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n981), .A2(new_n982), .A3(new_n712), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n712), .A2(new_n490), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n683), .B1(new_n978), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n973), .A2(new_n974), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n984), .A2(new_n987), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n978), .A2(new_n985), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n676), .A2(new_n680), .A3(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT106), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(KEYINPUT106), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(new_n993), .B2(new_n996), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n999), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(new_n989), .A3(new_n997), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n686), .A2(new_n991), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT45), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n686), .A2(new_n991), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT44), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n681), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1005), .A2(new_n681), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OR3_X1    g0812(.A1(new_n680), .A2(KEYINPUT108), .A3(new_n682), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT108), .B1(new_n680), .B2(new_n682), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n683), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n676), .B(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n739), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n739), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n689), .B(new_n1019), .Z(new_n1020));
  AOI21_X1  g0820(.A(new_n745), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n976), .B1(new_n1003), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT113), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n1016), .A2(new_n745), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n773), .A2(new_n241), .B1(new_n776), .B2(new_n814), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n325), .B(new_n1025), .C1(G50), .C2(new_n768), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n788), .A2(new_n271), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n307), .A2(new_n787), .B1(new_n780), .B2(new_n259), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G159), .A2(new_n792), .B1(new_n794), .B2(G97), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n768), .A2(G317), .B1(G303), .B2(new_n772), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT114), .B(G322), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n770), .B2(new_n779), .C1(new_n791), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT115), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n786), .A2(new_n831), .B1(new_n788), .B2(new_n593), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT49), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n267), .B1(new_n777), .B2(G326), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n523), .B2(new_n793), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT116), .Z(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1040), .A2(KEYINPUT49), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1031), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n761), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n691), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n749), .A2(new_n1049), .B1(new_n498), .B2(new_n688), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n231), .A2(new_n282), .ZN(new_n1051));
  AOI21_X1  g0851(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n259), .A2(KEYINPUT50), .A3(new_n239), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT50), .B1(new_n259), .B2(new_n239), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n691), .B(new_n1052), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n752), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1050), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n747), .B1(new_n1057), .B2(new_n762), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1048), .B(new_n1058), .C1(new_n680), .C2(new_n759), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1024), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1016), .A2(new_n739), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1017), .A2(new_n689), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  OAI221_X1 g0863(.A(new_n762), .B1(new_n478), .B2(new_n209), .C1(new_n947), .C2(new_n238), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n746), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n768), .A2(G159), .B1(new_n792), .B2(G150), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  OAI221_X1 g0867(.A(new_n267), .B1(new_n776), .B2(new_n817), .C1(new_n773), .C2(new_n258), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n786), .A2(new_n271), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n779), .A2(new_n239), .B1(new_n788), .B2(new_n241), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(G87), .C2(new_n794), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1067), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n768), .A2(G311), .B1(new_n792), .B2(G317), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n325), .B1(new_n776), .B2(new_n1033), .C1(new_n773), .C2(new_n593), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n779), .A2(new_n608), .B1(new_n793), .B2(new_n498), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n786), .A2(new_n523), .B1(new_n788), .B2(new_n831), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1065), .B1(new_n1080), .B2(new_n761), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n991), .B2(new_n759), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1011), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n681), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT117), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1010), .A2(new_n1086), .A3(new_n1011), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1087), .A3(new_n745), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n689), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1082), .B(new_n1088), .C1(new_n1089), .C2(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(new_n835), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G97), .A2(new_n772), .B1(new_n777), .B2(G294), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1093), .B(new_n325), .C1(new_n523), .C2(new_n804), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n822), .B(new_n1094), .C1(G87), .C2(new_n789), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n791), .A2(new_n831), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1096), .B(new_n1070), .C1(G107), .C2(new_n780), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n788), .A2(new_n814), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT53), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n804), .A2(new_n823), .B1(new_n773), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(G128), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n786), .A2(new_n799), .B1(new_n791), .B2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n779), .A2(new_n813), .B1(new_n793), .B2(new_n239), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n267), .B1(new_n776), .B2(new_n1105), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1095), .A2(new_n1097), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n746), .B1(new_n259), .B2(new_n1092), .C1(new_n1108), .C2(new_n765), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n925), .B1(new_n886), .B2(new_n920), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n756), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n849), .A2(new_n901), .A3(G330), .A4(new_n840), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n930), .A2(new_n901), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n926), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1113), .B1(new_n1115), .B2(new_n1110), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n669), .B(new_n840), .C1(new_n732), .C2(new_n737), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n929), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n901), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n927), .B1(new_n911), .B2(new_n885), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1121), .A3(KEYINPUT118), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT118), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n921), .A2(new_n883), .A3(new_n920), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT39), .B1(new_n911), .B2(new_n885), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n927), .B1(new_n930), .B2(new_n901), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1112), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1120), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1118), .B2(new_n901), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1123), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1115), .A2(new_n1110), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n898), .A2(G330), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n890), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n887), .B1(new_n388), .B2(new_n395), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1134), .A2(new_n1137), .A3(new_n843), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1122), .A2(new_n1131), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1111), .B1(new_n1139), .B2(new_n745), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n445), .A2(G330), .A3(new_n898), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n645), .A2(new_n935), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n901), .B1(new_n721), .B2(new_n840), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n930), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1137), .B1(new_n1134), .B2(new_n843), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(new_n929), .A3(new_n1117), .A4(new_n1112), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1142), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n689), .B1(new_n1139), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1132), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1138), .B1(new_n1149), .B2(new_n1130), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT118), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1128), .A2(new_n1130), .A3(new_n1123), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1147), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1140), .B1(new_n1148), .B2(new_n1154), .ZN(G378));
  INV_X1    g0955(.A(new_n293), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n644), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n296), .A2(new_n932), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n304), .B1(new_n296), .B2(new_n932), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n913), .B2(G330), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n901), .A2(new_n898), .A3(new_n840), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n921), .A2(new_n883), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n900), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n912), .A2(new_n898), .A3(new_n891), .ZN(new_n1171));
  AND4_X1   g0971(.A1(G330), .A2(new_n1170), .A3(new_n1166), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n934), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n913), .A2(G330), .A3(new_n1166), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1171), .A3(G330), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1166), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n934), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n756), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n746), .B1(G50), .B2(new_n1092), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n325), .A2(new_n281), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n239), .C1(G33), .C2(G41), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT119), .Z(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(G283), .B2(new_n777), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n306), .B2(new_n773), .C1(new_n804), .C2(new_n498), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G116), .A2(new_n792), .B1(new_n794), .B2(G58), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n478), .B2(new_n779), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1187), .A2(new_n1189), .A3(new_n962), .A4(new_n1027), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1185), .B1(new_n1190), .B2(KEYINPUT58), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n773), .A2(new_n813), .B1(new_n779), .B2(new_n823), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT120), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n804), .A2(new_n1102), .B1(new_n814), .B2(new_n786), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n791), .A2(new_n1105), .B1(new_n788), .B2(new_n1100), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n794), .A2(G159), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n777), .C2(G124), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1191), .B1(KEYINPUT58), .B2(new_n1190), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1182), .B1(new_n1203), .B2(new_n761), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1180), .A2(new_n745), .B1(new_n1181), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1142), .B1(new_n1139), .B2(new_n1147), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1167), .A2(new_n1172), .A3(new_n934), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1178), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n689), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1142), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1153), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1180), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1205), .B1(new_n1210), .B2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n745), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n786), .A2(new_n239), .B1(new_n791), .B2(new_n823), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G159), .B2(new_n789), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n325), .B1(new_n777), .B2(G128), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n768), .A2(G137), .B1(G150), .B2(new_n772), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1100), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n780), .A2(new_n1221), .B1(new_n794), .B2(G58), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n804), .A2(new_n831), .B1(new_n773), .B2(new_n498), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n307), .B2(new_n787), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n325), .B1(new_n793), .B2(new_n271), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1226), .A2(KEYINPUT121), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(KEYINPUT121), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G116), .A2(new_n780), .B1(new_n792), .B2(G294), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n788), .A2(new_n478), .B1(new_n776), .B2(new_n608), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1223), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n765), .B1(new_n1233), .B2(KEYINPUT123), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(KEYINPUT123), .B2(new_n1233), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n747), .B1(new_n241), .B2(new_n835), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n901), .C2(new_n757), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1216), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1147), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1144), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1020), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(G381));
  OR2_X1    g1043(.A1(new_n1062), .A2(new_n1061), .ZN(new_n1244));
  INV_X1    g1044(.A(G396), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1060), .ZN(new_n1246));
  OR4_X1    g1046(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1246), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(G387), .A2(new_n1247), .A3(G378), .A4(G375), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT124), .ZN(G407));
  OR2_X1    g1049(.A1(G378), .A2(G343), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G375), .C2(new_n1250), .ZN(G409));
  OAI211_X1 g1051(.A(G378), .B(new_n1205), .C1(new_n1210), .C2(new_n1213), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1150), .B(new_n745), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1111), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n690), .B1(new_n1256), .B2(new_n1240), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1257), .B2(new_n1153), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1020), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1206), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1180), .A2(new_n745), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1181), .A2(new_n1204), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1252), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n1142), .A4(new_n1146), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1270), .A2(new_n689), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1241), .B1(new_n1147), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1239), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n857), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G384), .A2(new_n1239), .A3(new_n1274), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1266), .A2(new_n1269), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1245), .B1(new_n1244), .B2(new_n1060), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  OAI21_X1  g1083(.A(G390), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT113), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G393), .A2(G396), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1246), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1287), .B2(G390), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1022), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1284), .B(new_n1022), .C1(G390), .C2(new_n1287), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1268), .B(new_n1278), .C1(new_n1252), .C2(new_n1265), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1281), .B(new_n1292), .C1(new_n1293), .C2(KEYINPUT63), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1268), .B1(new_n1252), .B2(new_n1265), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1268), .A2(G2897), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1275), .A2(new_n857), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1274), .A2(new_n1239), .B1(new_n854), .B2(new_n856), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1298), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1276), .A2(new_n1277), .A3(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1295), .B1(new_n1296), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT125), .B1(new_n1294), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1296), .B2(new_n1280), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1266), .A2(new_n1269), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1279), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1306), .A2(new_n1308), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1305), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1304), .A2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(KEYINPUT126), .B(new_n1295), .C1(new_n1296), .C2(new_n1303), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1293), .A2(new_n1318), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1307), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1313), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1313), .A2(new_n1321), .A3(KEYINPUT127), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(G405));
  XNOR2_X1  g1126(.A(G375), .B(G378), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1278), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1327), .B(new_n1328), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1292), .ZN(G402));
endmodule


