

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597;

  XOR2_X2 U326 ( .A(n458), .B(n457), .Z(n575) );
  XOR2_X1 U327 ( .A(KEYINPUT124), .B(n574), .Z(n294) );
  XOR2_X1 U328 ( .A(G176GAT), .B(G71GAT), .Z(n295) );
  AND2_X1 U329 ( .A1(n582), .A2(n546), .ZN(n518) );
  OR2_X1 U330 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U331 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U332 ( .A(n588), .B(KEYINPUT41), .Z(n546) );
  XOR2_X1 U333 ( .A(n412), .B(KEYINPUT28), .Z(n531) );
  XOR2_X1 U334 ( .A(KEYINPUT6), .B(G1GAT), .Z(n297) );
  XNOR2_X1 U335 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n296) );
  XNOR2_X1 U336 ( .A(n297), .B(n296), .ZN(n316) );
  XOR2_X1 U337 ( .A(G141GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U338 ( .A(G29GAT), .B(G85GAT), .ZN(n298) );
  XNOR2_X1 U339 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U340 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n301) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(G120GAT), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U343 ( .A(n303), .B(n302), .Z(n309) );
  XNOR2_X1 U344 ( .A(G127GAT), .B(KEYINPUT80), .ZN(n304) );
  XNOR2_X1 U345 ( .A(n304), .B(KEYINPUT0), .ZN(n383) );
  XOR2_X1 U346 ( .A(G134GAT), .B(n383), .Z(n306) );
  NAND2_X1 U347 ( .A1(G225GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U348 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U349 ( .A(G162GAT), .B(n307), .ZN(n308) );
  XNOR2_X1 U350 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U351 ( .A(n310), .B(KEYINPUT93), .Z(n314) );
  XOR2_X1 U352 ( .A(G155GAT), .B(KEYINPUT2), .Z(n312) );
  XNOR2_X1 U353 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n311) );
  XNOR2_X1 U354 ( .A(n312), .B(n311), .ZN(n363) );
  XNOR2_X1 U355 ( .A(n363), .B(KEYINPUT94), .ZN(n313) );
  XNOR2_X1 U356 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U357 ( .A(n316), .B(n315), .ZN(n561) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(G43GAT), .ZN(n317) );
  XNOR2_X1 U359 ( .A(n317), .B(G15GAT), .ZN(n379) );
  XOR2_X1 U360 ( .A(G141GAT), .B(G22GAT), .Z(n358) );
  XOR2_X1 U361 ( .A(n379), .B(n358), .Z(n319) );
  NAND2_X1 U362 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U363 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U364 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n321) );
  XNOR2_X1 U365 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U367 ( .A(n323), .B(n322), .Z(n336) );
  INV_X1 U368 ( .A(G29GAT), .ZN(n331) );
  INV_X1 U369 ( .A(KEYINPUT7), .ZN(n324) );
  NAND2_X1 U370 ( .A1(G50GAT), .A2(n324), .ZN(n327) );
  INV_X1 U371 ( .A(G50GAT), .ZN(n325) );
  NAND2_X1 U372 ( .A1(n325), .A2(KEYINPUT7), .ZN(n326) );
  NAND2_X1 U373 ( .A1(n327), .A2(n326), .ZN(n329) );
  XNOR2_X1 U374 ( .A(KEYINPUT8), .B(G36GAT), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U376 ( .A(n331), .B(n330), .ZN(n438) );
  XOR2_X1 U377 ( .A(KEYINPUT30), .B(G169GAT), .Z(n333) );
  XNOR2_X1 U378 ( .A(G1GAT), .B(G197GAT), .ZN(n332) );
  XNOR2_X1 U379 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U380 ( .A(n438), .B(n334), .ZN(n335) );
  XOR2_X1 U381 ( .A(n336), .B(n335), .Z(n582) );
  XNOR2_X1 U382 ( .A(KEYINPUT69), .B(n582), .ZN(n566) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(G99GAT), .ZN(n337) );
  XNOR2_X1 U384 ( .A(n295), .B(n337), .ZN(n380) );
  XNOR2_X1 U385 ( .A(n380), .B(KEYINPUT74), .ZN(n339) );
  AND2_X1 U386 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U387 ( .A(n339), .B(n338), .ZN(n344) );
  XNOR2_X1 U388 ( .A(G78GAT), .B(KEYINPUT71), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n340), .B(KEYINPUT72), .ZN(n341) );
  XOR2_X1 U390 ( .A(n341), .B(G204GAT), .Z(n343) );
  XNOR2_X1 U391 ( .A(G148GAT), .B(G106GAT), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n369) );
  XNOR2_X1 U393 ( .A(n344), .B(n369), .ZN(n352) );
  XOR2_X1 U394 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n346) );
  XNOR2_X1 U395 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U397 ( .A(G92GAT), .B(G64GAT), .Z(n392) );
  XOR2_X1 U398 ( .A(n347), .B(n392), .Z(n350) );
  XOR2_X1 U399 ( .A(G85GAT), .B(KEYINPUT73), .Z(n441) );
  XNOR2_X1 U400 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n348), .B(KEYINPUT13), .ZN(n430) );
  XNOR2_X1 U402 ( .A(n441), .B(n430), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n588) );
  NOR2_X1 U405 ( .A1(n566), .A2(n588), .ZN(n480) );
  INV_X1 U406 ( .A(n561), .ZN(n492) );
  XOR2_X1 U407 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n354) );
  NAND2_X1 U408 ( .A1(G228GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U410 ( .A(KEYINPUT92), .B(n355), .ZN(n367) );
  XOR2_X1 U411 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n357) );
  XNOR2_X1 U412 ( .A(KEYINPUT91), .B(KEYINPUT22), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n359) );
  XOR2_X1 U414 ( .A(n359), .B(n358), .Z(n361) );
  XNOR2_X1 U415 ( .A(G50GAT), .B(G211GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U417 ( .A(KEYINPUT21), .B(G197GAT), .Z(n401) );
  XOR2_X1 U418 ( .A(n362), .B(n401), .Z(n365) );
  XOR2_X1 U419 ( .A(G162GAT), .B(G218GAT), .Z(n455) );
  XNOR2_X1 U420 ( .A(n363), .B(n455), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U423 ( .A(n369), .B(n368), .Z(n562) );
  XOR2_X1 U424 ( .A(KEYINPUT85), .B(KEYINPUT81), .Z(n371) );
  XNOR2_X1 U425 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n378) );
  XOR2_X1 U427 ( .A(G134GAT), .B(G190GAT), .Z(n437) );
  XOR2_X1 U428 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n373) );
  XNOR2_X1 U429 ( .A(G183GAT), .B(KEYINPUT86), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U431 ( .A(n437), .B(n374), .Z(n376) );
  NAND2_X1 U432 ( .A1(G227GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n387) );
  XOR2_X1 U435 ( .A(n380), .B(n379), .Z(n385) );
  XOR2_X1 U436 ( .A(G169GAT), .B(KEYINPUT19), .Z(n382) );
  XNOR2_X1 U437 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n397) );
  XNOR2_X1 U439 ( .A(n383), .B(n397), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U441 ( .A(n387), .B(n386), .Z(n564) );
  NOR2_X1 U442 ( .A1(n562), .A2(n564), .ZN(n389) );
  XNOR2_X1 U443 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n580) );
  XOR2_X1 U445 ( .A(KEYINPUT95), .B(G176GAT), .Z(n391) );
  XNOR2_X1 U446 ( .A(G36GAT), .B(G204GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n395) );
  XNOR2_X1 U448 ( .A(G218GAT), .B(G190GAT), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U450 ( .A(n395), .B(n394), .Z(n399) );
  XNOR2_X1 U451 ( .A(G211GAT), .B(G183GAT), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n396), .B(G8GAT), .ZN(n429) );
  XNOR2_X1 U453 ( .A(n429), .B(n397), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U455 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n495) );
  XOR2_X1 U458 ( .A(n495), .B(KEYINPUT27), .Z(n414) );
  NOR2_X1 U459 ( .A1(n580), .A2(n414), .ZN(n404) );
  XNOR2_X1 U460 ( .A(KEYINPUT98), .B(n404), .ZN(n409) );
  INV_X1 U461 ( .A(n562), .ZN(n412) );
  INV_X1 U462 ( .A(n495), .ZN(n558) );
  INV_X1 U463 ( .A(n564), .ZN(n530) );
  NOR2_X1 U464 ( .A1(n558), .A2(n530), .ZN(n405) );
  XOR2_X1 U465 ( .A(KEYINPUT99), .B(n405), .Z(n406) );
  NOR2_X1 U466 ( .A1(n412), .A2(n406), .ZN(n407) );
  XOR2_X1 U467 ( .A(KEYINPUT25), .B(n407), .Z(n408) );
  NOR2_X1 U468 ( .A1(n409), .A2(n408), .ZN(n410) );
  NOR2_X1 U469 ( .A1(n492), .A2(n410), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n411), .B(KEYINPUT100), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(n530), .Z(n413) );
  NAND2_X1 U472 ( .A1(n413), .A2(n531), .ZN(n416) );
  OR2_X1 U473 ( .A1(n414), .A2(n561), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n415), .B(KEYINPUT96), .ZN(n528) );
  NOR2_X1 U475 ( .A1(n416), .A2(n528), .ZN(n417) );
  NOR2_X1 U476 ( .A1(n418), .A2(n417), .ZN(n473) );
  XOR2_X1 U477 ( .A(G71GAT), .B(G15GAT), .Z(n420) );
  XNOR2_X1 U478 ( .A(G127GAT), .B(G22GAT), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U480 ( .A(G155GAT), .B(G78GAT), .Z(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n434) );
  XOR2_X1 U482 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n424) );
  XNOR2_X1 U483 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n426) );
  XNOR2_X1 U486 ( .A(G1GAT), .B(G64GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U488 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n436) );
  NAND2_X1 U492 ( .A1(G231GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n591) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n440) );
  XNOR2_X1 U496 ( .A(KEYINPUT11), .B(KEYINPUT76), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U498 ( .A(n442), .B(n441), .Z(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n447) );
  XOR2_X1 U500 ( .A(G92GAT), .B(G43GAT), .Z(n446) );
  NAND2_X1 U501 ( .A1(G232GAT), .A2(G233GAT), .ZN(n445) );
  XOR2_X1 U502 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U503 ( .A1(n447), .A2(n448), .ZN(n452) );
  INV_X1 U504 ( .A(n447), .ZN(n450) );
  INV_X1 U505 ( .A(n448), .ZN(n449) );
  NAND2_X1 U506 ( .A1(n450), .A2(n449), .ZN(n451) );
  NAND2_X1 U507 ( .A1(n452), .A2(n451), .ZN(n458) );
  XOR2_X1 U508 ( .A(G99GAT), .B(G106GAT), .Z(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n591), .A2(n575), .ZN(n459) );
  XNOR2_X1 U513 ( .A(KEYINPUT16), .B(n459), .ZN(n460) );
  NOR2_X1 U514 ( .A1(n473), .A2(n460), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT101), .B(n461), .Z(n490) );
  NAND2_X1 U516 ( .A1(n480), .A2(n490), .ZN(n470) );
  NOR2_X1 U517 ( .A1(n561), .A2(n470), .ZN(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U520 ( .A(G1GAT), .B(n464), .Z(G1324GAT) );
  NOR2_X1 U521 ( .A1(n558), .A2(n470), .ZN(n466) );
  XNOR2_X1 U522 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(G1325GAT) );
  NOR2_X1 U524 ( .A1(n530), .A2(n470), .ZN(n468) );
  XNOR2_X1 U525 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U527 ( .A(G15GAT), .B(n469), .ZN(G1326GAT) );
  NOR2_X1 U528 ( .A1(n531), .A2(n470), .ZN(n472) );
  XNOR2_X1 U529 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(G1327GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT38), .B(KEYINPUT107), .Z(n482) );
  NOR2_X1 U532 ( .A1(n591), .A2(n473), .ZN(n474) );
  XNOR2_X1 U533 ( .A(KEYINPUT106), .B(n474), .ZN(n478) );
  INV_X1 U534 ( .A(KEYINPUT36), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n475), .A2(n575), .ZN(n477) );
  INV_X1 U536 ( .A(n575), .ZN(n554) );
  NAND2_X1 U537 ( .A1(KEYINPUT36), .A2(n554), .ZN(n476) );
  NAND2_X1 U538 ( .A1(n477), .A2(n476), .ZN(n595) );
  NAND2_X1 U539 ( .A1(n478), .A2(n595), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT37), .ZN(n504) );
  NAND2_X1 U541 ( .A1(n480), .A2(n504), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n488) );
  NOR2_X1 U543 ( .A1(n561), .A2(n488), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n483), .B(KEYINPUT39), .ZN(n484) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(n484), .ZN(G1328GAT) );
  NOR2_X1 U546 ( .A1(n558), .A2(n488), .ZN(n485) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n485), .Z(G1329GAT) );
  NOR2_X1 U548 ( .A1(n530), .A2(n488), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT40), .B(n486), .Z(n487) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n487), .ZN(G1330GAT) );
  NOR2_X1 U551 ( .A1(n488), .A2(n531), .ZN(n489) );
  XOR2_X1 U552 ( .A(G50GAT), .B(n489), .Z(G1331GAT) );
  XNOR2_X1 U553 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n494) );
  INV_X1 U554 ( .A(n546), .ZN(n568) );
  NOR2_X1 U555 ( .A1(n582), .A2(n568), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n490), .A2(n503), .ZN(n491) );
  XOR2_X1 U557 ( .A(KEYINPUT108), .B(n491), .Z(n498) );
  NAND2_X1 U558 ( .A1(n492), .A2(n498), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(G1332GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n495), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U562 ( .A1(n498), .A2(n564), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n497), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n501) );
  INV_X1 U565 ( .A(n531), .ZN(n499) );
  NAND2_X1 U566 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U568 ( .A(G78GAT), .B(n502), .Z(G1335GAT) );
  NAND2_X1 U569 ( .A1(n504), .A2(n503), .ZN(n509) );
  NOR2_X1 U570 ( .A1(n561), .A2(n509), .ZN(n505) );
  XOR2_X1 U571 ( .A(G85GAT), .B(n505), .Z(n506) );
  XNOR2_X1 U572 ( .A(KEYINPUT110), .B(n506), .ZN(G1336GAT) );
  NOR2_X1 U573 ( .A1(n558), .A2(n509), .ZN(n507) );
  XOR2_X1 U574 ( .A(G92GAT), .B(n507), .Z(G1337GAT) );
  NOR2_X1 U575 ( .A1(n530), .A2(n509), .ZN(n508) );
  XOR2_X1 U576 ( .A(G99GAT), .B(n508), .Z(G1338GAT) );
  NOR2_X1 U577 ( .A1(n531), .A2(n509), .ZN(n510) );
  XOR2_X1 U578 ( .A(KEYINPUT44), .B(n510), .Z(n511) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(n511), .ZN(G1339GAT) );
  INV_X1 U580 ( .A(KEYINPUT115), .ZN(n515) );
  NAND2_X1 U581 ( .A1(n591), .A2(n595), .ZN(n512) );
  XNOR2_X1 U582 ( .A(KEYINPUT45), .B(n512), .ZN(n513) );
  NOR2_X1 U583 ( .A1(n513), .A2(n588), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U585 ( .A1(n516), .A2(n566), .ZN(n525) );
  XNOR2_X1 U586 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n591), .B(KEYINPUT111), .ZN(n573) );
  NAND2_X1 U589 ( .A1(n573), .A2(n575), .ZN(n519) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U593 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n526), .B(KEYINPUT48), .ZN(n527) );
  XOR2_X1 U595 ( .A(KEYINPUT64), .B(n527), .Z(n557) );
  NOR2_X1 U596 ( .A1(n528), .A2(n557), .ZN(n529) );
  XOR2_X1 U597 ( .A(KEYINPUT116), .B(n529), .Z(n543) );
  NOR2_X1 U598 ( .A1(n530), .A2(n543), .ZN(n532) );
  NAND2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n566), .A2(n538), .ZN(n533) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  NOR2_X1 U602 ( .A1(n568), .A2(n538), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n573), .A2(n538), .ZN(n536) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n536), .Z(n537) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  NOR2_X1 U608 ( .A1(n538), .A2(n575), .ZN(n542) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n540) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT117), .ZN(n539) );
  XNOR2_X1 U611 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U612 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  XOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT119), .Z(n545) );
  NOR2_X1 U614 ( .A1(n580), .A2(n543), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n555), .A2(n582), .ZN(n544) );
  XNOR2_X1 U616 ( .A(n545), .B(n544), .ZN(G1344GAT) );
  XNOR2_X1 U617 ( .A(KEYINPUT52), .B(KEYINPUT120), .ZN(n550) );
  XOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .Z(n548) );
  NAND2_X1 U619 ( .A1(n555), .A2(n546), .ZN(n547) );
  XNOR2_X1 U620 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U621 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n552) );
  NAND2_X1 U623 ( .A1(n555), .A2(n591), .ZN(n551) );
  XNOR2_X1 U624 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U627 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U628 ( .A(KEYINPUT54), .B(n559), .ZN(n560) );
  AND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n579) );
  NAND2_X1 U630 ( .A1(n562), .A2(n579), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT55), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n576) );
  NOR2_X1 U633 ( .A1(n566), .A2(n576), .ZN(n567) );
  XOR2_X1 U634 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  NOR2_X1 U635 ( .A1(n576), .A2(n568), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n570) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NOR2_X1 U640 ( .A1(n573), .A2(n576), .ZN(n574) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(n294), .ZN(G1350GAT) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G190GAT), .B(n577), .Z(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT58), .B(n578), .ZN(G1351GAT) );
  INV_X1 U645 ( .A(n579), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n594) );
  AND2_X1 U647 ( .A1(n582), .A2(n594), .ZN(n587) );
  XOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(KEYINPUT59), .B(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .Z(n590) );
  NAND2_X1 U654 ( .A1(n594), .A2(n588), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  XOR2_X1 U656 ( .A(G211GAT), .B(KEYINPUT127), .Z(n593) );
  NAND2_X1 U657 ( .A1(n594), .A2(n591), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1354GAT) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(KEYINPUT62), .ZN(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

