//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n193), .A2(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n196), .A3(KEYINPUT16), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(G146), .A3(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G128), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT24), .B(G110), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n204), .B(new_n210), .C1(new_n211), .C2(KEYINPUT23), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n212), .B2(G110), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT72), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n214), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n202), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n207), .A2(new_n208), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(G110), .B2(new_n212), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n194), .A2(G146), .A3(new_n197), .ZN(new_n221));
  AOI21_X1  g035(.A(G146), .B1(new_n194), .B2(new_n197), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n191), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n217), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n198), .B(new_n201), .C1(new_n226), .C2(new_n215), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n223), .A3(new_n190), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G217), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(G234), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G902), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT75), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n225), .A2(new_n228), .A3(new_n232), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT73), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n229), .A2(new_n241), .A3(KEYINPUT25), .A4(new_n232), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT74), .B1(new_n237), .B2(new_n238), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT73), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n237), .A2(new_n244), .A3(new_n238), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n242), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n236), .B1(new_n246), .B2(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(KEYINPUT32), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT11), .B1(new_n252), .B2(G137), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT65), .B1(new_n255), .B2(G134), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n252), .A3(G137), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n257), .A2(new_n258), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n255), .A2(G134), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n252), .A2(G137), .ZN(new_n264));
  OAI21_X1  g078(.A(G131), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n200), .A2(G143), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G146), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n269), .A2(KEYINPUT64), .A3(G146), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT64), .B1(new_n269), .B2(G146), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT1), .B1(new_n269), .B2(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G128), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n271), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT66), .B1(new_n266), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n268), .A2(new_n270), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n274), .A2(new_n282), .B1(new_n284), .B2(new_n280), .ZN(new_n285));
  INV_X1    g099(.A(new_n262), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n259), .A2(new_n261), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n258), .B1(new_n287), .B2(new_n257), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT2), .B(G113), .ZN(new_n290));
  INV_X1    g104(.A(G116), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(G119), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n203), .A2(G116), .ZN(new_n293));
  OR3_X1    g107(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(G116), .B(G119), .Z(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n290), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n269), .A2(G146), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT64), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n200), .B2(G143), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n269), .A2(KEYINPUT64), .A3(G146), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n205), .B1(new_n268), .B2(KEYINPUT1), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n265), .A4(new_n262), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n278), .A2(new_n289), .A3(new_n298), .A4(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G237), .A2(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G210), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT27), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(G101), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n306), .A2(new_n265), .A3(new_n262), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n289), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n278), .A2(new_n289), .A3(new_n308), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(KEYINPUT30), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n251), .B(new_n316), .C1(new_n321), .C2(new_n298), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n289), .A2(new_n298), .A3(new_n318), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n289), .A2(new_n318), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n297), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n325), .B(new_n327), .C1(new_n324), .C2(new_n309), .ZN(new_n328));
  INV_X1    g142(.A(new_n314), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n320), .A2(KEYINPUT30), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n289), .A2(new_n317), .A3(new_n318), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n298), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT31), .B1(new_n334), .B2(new_n315), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT67), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(KEYINPUT31), .C1(new_n334), .C2(new_n315), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n331), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(G472), .A2(G902), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n250), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n322), .A2(new_n330), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n316), .B1(new_n321), .B2(new_n298), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n337), .B1(new_n344), .B2(KEYINPUT31), .ZN(new_n345));
  INV_X1    g159(.A(new_n338), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT32), .A3(new_n340), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G472), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n332), .A2(new_n333), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n297), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n314), .B1(new_n352), .B2(new_n309), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT69), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n328), .B2(new_n329), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n325), .A2(new_n327), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n309), .A2(new_n324), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n360), .B2(new_n314), .ZN(new_n361));
  INV_X1    g175(.A(new_n309), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n329), .B1(new_n334), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT69), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n320), .A2(new_n297), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT70), .A3(new_n309), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT70), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n320), .A2(new_n368), .A3(new_n297), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(KEYINPUT28), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT29), .A3(new_n314), .A4(new_n325), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(new_n232), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n350), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT71), .B1(new_n349), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n354), .B1(new_n353), .B2(new_n356), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n361), .A2(KEYINPUT69), .A3(new_n363), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G472), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT71), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n348), .A4(new_n342), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n248), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G104), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n385), .A3(G104), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n387), .A2(new_n390), .A3(new_n385), .A4(G104), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n384), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n383), .A2(new_n392), .B1(new_n294), .B2(new_n296), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G107), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n395), .A2(KEYINPUT76), .A3(G107), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(new_n390), .ZN(new_n398));
  INV_X1    g212(.A(new_n391), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n394), .B(G101), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n401), .A2(new_n384), .A3(new_n391), .A4(new_n396), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n392), .A2(new_n394), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n393), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G122), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n395), .A2(G107), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n408), .B2(new_n386), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G113), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n292), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n295), .B2(new_n413), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n294), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n393), .B(new_n417), .C1(new_n403), .C2(new_n404), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n406), .A2(new_n407), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n418), .A2(new_n416), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n422), .A2(KEYINPUT85), .A3(new_n407), .A4(new_n406), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n406), .ZN(new_n426));
  INV_X1    g240(.A(new_n407), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n418), .A2(new_n416), .ZN(new_n430));
  OAI21_X1  g244(.A(G101), .B1(new_n398), .B2(new_n399), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n400), .A4(new_n402), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n417), .B1(new_n433), .B2(new_n393), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n425), .B(new_n427), .C1(new_n430), .C2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n280), .A2(new_n281), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n304), .A2(new_n436), .B1(new_n283), .B2(new_n279), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G125), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(G125), .B2(new_n306), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n188), .A2(G224), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n429), .A2(new_n435), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(KEYINPUT7), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n439), .B(new_n444), .Z(new_n445));
  XNOR2_X1  g259(.A(new_n407), .B(KEYINPUT8), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n415), .A2(new_n294), .A3(new_n410), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n414), .B1(new_n448), .B2(new_n295), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n449), .A2(new_n294), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n446), .B(new_n447), .C1(new_n450), .C2(new_n410), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G902), .B1(new_n424), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G210), .B1(G237), .B2(G902), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n443), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n443), .B2(new_n453), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n382), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n382), .ZN(new_n461));
  INV_X1    g275(.A(new_n454), .ZN(new_n462));
  INV_X1    g276(.A(new_n435), .ZN(new_n463));
  AOI211_X1 g277(.A(new_n441), .B(new_n463), .C1(new_n424), .C2(new_n428), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n424), .A2(new_n452), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n232), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n461), .B1(new_n467), .B2(new_n455), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT86), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT9), .B(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(G221), .B1(new_n470), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n291), .A2(G122), .ZN(new_n473));
  INV_X1    g287(.A(G122), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT92), .B1(new_n474), .B2(G116), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n291), .A3(G122), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n385), .ZN(new_n479));
  XNOR2_X1  g293(.A(G128), .B(G143), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(new_n252), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n477), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n483), .A2(new_n484), .A3(new_n473), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n479), .B(new_n481), .C1(new_n485), .C2(new_n385), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n269), .A2(KEYINPUT13), .A3(G128), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n487), .B(KEYINPUT93), .C1(G128), .C2(new_n269), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT13), .B1(new_n269), .B2(G128), .ZN(new_n489));
  OAI221_X1 g303(.A(G134), .B1(KEYINPUT93), .B2(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n480), .A2(new_n252), .ZN(new_n491));
  INV_X1    g305(.A(new_n479), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n478), .A2(new_n385), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n490), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n470), .A2(new_n231), .A3(G953), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n486), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n486), .B2(new_n494), .ZN(new_n497));
  OAI211_X1 g311(.A(KEYINPUT94), .B(new_n232), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G478), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n500), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n188), .A2(G952), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(G234), .B2(G237), .ZN(new_n505));
  AOI211_X1 g319(.A(new_n232), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT21), .B(G898), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n221), .A2(new_n222), .ZN(new_n510));
  INV_X1    g324(.A(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n188), .A3(G214), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n269), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n310), .A2(G143), .A3(G214), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n258), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n515), .A2(KEYINPUT88), .A3(KEYINPUT17), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT88), .B1(new_n515), .B2(KEYINPUT17), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n519));
  INV_X1    g333(.A(new_n514), .ZN(new_n520));
  AOI21_X1  g334(.A(G143), .B1(new_n310), .B2(G214), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n513), .A2(new_n258), .A3(new_n514), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n510), .B(new_n528), .C1(new_n516), .C2(new_n517), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n199), .B(new_n200), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT18), .B(G131), .C1(new_n520), .C2(new_n521), .ZN(new_n532));
  NAND2_X1  g346(.A1(KEYINPUT18), .A2(G131), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n513), .A2(new_n514), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G113), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT87), .B(G104), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n536), .B(new_n537), .Z(new_n538));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n522), .A2(new_n524), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n199), .B(KEYINPUT19), .Z(new_n541));
  OAI211_X1 g355(.A(new_n198), .B(new_n540), .C1(new_n541), .C2(G146), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(new_n535), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G475), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(KEYINPUT20), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT20), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n546), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n530), .A2(new_n535), .A3(new_n538), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n538), .B1(new_n530), .B2(new_n535), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n232), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n549), .A2(new_n550), .B1(new_n553), .B2(G475), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n509), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G140), .ZN(new_n556));
  INV_X1    g370(.A(G227), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G953), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n286), .A2(new_n288), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n275), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n268), .A2(KEYINPUT78), .A3(KEYINPUT1), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(G128), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n271), .B1(new_n564), .B2(new_n283), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(new_n410), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n306), .B1(new_n402), .B2(new_n409), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT12), .B(new_n560), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n410), .A2(new_n277), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n410), .B2(new_n565), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT79), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT12), .A4(new_n560), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n560), .B1(new_n566), .B2(new_n567), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n437), .B1(new_n383), .B2(new_n392), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n403), .B2(new_n404), .ZN(new_n579));
  INV_X1    g393(.A(new_n560), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n565), .B2(new_n410), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n411), .A2(KEYINPUT10), .A3(new_n306), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n579), .A2(new_n580), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n577), .A2(KEYINPUT80), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT80), .B1(new_n577), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n559), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n559), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n560), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n587), .A2(G469), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(G469), .A2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n588), .B1(new_n592), .B2(new_n584), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT81), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n569), .A2(new_n576), .A3(new_n600), .A4(new_n573), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n601), .A3(new_n590), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n598), .B1(new_n602), .B2(KEYINPUT82), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n589), .B1(new_n577), .B2(KEYINPUT81), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT82), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n601), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n232), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n472), .B(new_n555), .C1(new_n597), .C2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n381), .A2(new_n460), .A3(new_n469), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AOI211_X1 g426(.A(G469), .B(G902), .C1(new_n603), .C2(new_n606), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n471), .B1(new_n613), .B2(new_n596), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n339), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n347), .A2(new_n340), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n247), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n549), .A2(new_n550), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n553), .A2(G475), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n619), .A2(new_n548), .A3(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n499), .B(new_n232), .C1(new_n496), .C2(new_n497), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n499), .A2(new_n232), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT33), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n486), .A2(new_n494), .ZN(new_n628));
  INV_X1    g442(.A(new_n495), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n486), .A2(new_n494), .A3(new_n495), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n625), .B1(new_n633), .B2(G478), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n621), .A2(new_n508), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n468), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n618), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(new_n508), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n550), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n503), .A2(new_n620), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n468), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n618), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NAND2_X1  g463(.A1(new_n227), .A2(new_n223), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n235), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n246), .B2(new_n233), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n656), .A2(new_n616), .A3(new_n615), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n610), .A2(new_n460), .A3(new_n469), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT95), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n506), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n505), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n643), .A2(new_n644), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n656), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n374), .B2(new_n380), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n614), .A2(new_n458), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT96), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  NAND3_X1  g490(.A1(new_n619), .A2(new_n548), .A3(new_n620), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n503), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n678), .A2(new_n656), .A3(new_n461), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n352), .A2(new_n309), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n314), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n367), .A2(new_n369), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n329), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(KEYINPUT97), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n232), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT97), .B1(new_n681), .B2(new_n683), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n348), .A3(new_n342), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n679), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n472), .B1(new_n597), .B2(new_n609), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n665), .B(KEYINPUT39), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n692), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT40), .B1(new_n614), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n467), .A2(new_n455), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT38), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n467), .A2(KEYINPUT38), .A3(new_n455), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n689), .A2(new_n693), .A3(new_n695), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  NAND4_X1  g516(.A1(new_n656), .A2(new_n677), .A3(new_n634), .A4(new_n665), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n374), .B2(new_n380), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n670), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT98), .B(G146), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G48));
  AND3_X1   g521(.A1(new_n604), .A2(new_n605), .A3(new_n601), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n605), .B1(new_n604), .B2(new_n601), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n598), .ZN(new_n710));
  OAI21_X1  g524(.A(G469), .B1(new_n710), .B2(G902), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n471), .A3(new_n609), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n381), .A2(new_n637), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND2_X1  g530(.A1(new_n374), .A2(new_n380), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n646), .A3(new_n247), .A4(new_n713), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NOR2_X1   g533(.A1(new_n712), .A2(new_n458), .ZN(new_n720));
  INV_X1    g534(.A(new_n555), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n717), .A3(new_n721), .A4(new_n656), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT99), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n655), .B1(new_n374), .B2(new_n380), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT99), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n720), .A4(new_n721), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NAND2_X1  g542(.A1(new_n246), .A2(new_n233), .ZN(new_n729));
  INV_X1    g543(.A(new_n236), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT101), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT101), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n732), .B(new_n236), .C1(new_n246), .C2(new_n233), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n314), .B1(new_n370), .B2(new_n325), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n335), .A2(new_n322), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n340), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n615), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n458), .A2(new_n508), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT102), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n678), .B(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n742), .A3(new_n713), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT103), .B(G122), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G24));
  NOR2_X1   g561(.A1(new_n621), .A2(new_n635), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n665), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n656), .A2(new_n738), .A3(new_n615), .A4(new_n739), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n720), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  NAND3_X1  g567(.A1(new_n467), .A2(new_n382), .A3(new_n455), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n614), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n731), .A2(new_n733), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT32), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n616), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n378), .A2(new_n759), .A3(new_n348), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n756), .A2(new_n761), .A3(new_n762), .A4(new_n749), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n749), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n717), .A2(new_n755), .A3(new_n247), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n766), .A2(new_n767), .A3(new_n762), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n766), .B2(new_n762), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND3_X1  g585(.A1(new_n381), .A2(new_n667), .A3(new_n755), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND3_X1  g587(.A1(new_n587), .A2(KEYINPUT45), .A3(new_n593), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  INV_X1    g591(.A(new_n586), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n577), .A2(KEYINPUT80), .A3(new_n584), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n588), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n593), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n587), .A2(KEYINPUT105), .A3(KEYINPUT45), .A4(new_n593), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n776), .A2(G469), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n595), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n613), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(KEYINPUT106), .A3(KEYINPUT46), .A4(new_n595), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n595), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT106), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n619), .A2(new_n634), .A3(new_n548), .A4(new_n620), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT43), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(KEYINPUT107), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n554), .A2(new_n548), .A3(new_n634), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n655), .B1(new_n615), .B2(new_n616), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n801), .A2(KEYINPUT44), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT44), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n803), .A2(new_n804), .A3(new_n754), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n792), .A2(new_n805), .A3(new_n471), .A4(new_n692), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  NOR4_X1   g621(.A1(new_n717), .A2(new_n247), .A3(new_n749), .A4(new_n754), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n471), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT47), .B1(new_n792), .B2(new_n471), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT108), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  AND3_X1   g630(.A1(new_n714), .A2(new_n718), .A3(new_n745), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n677), .B1(new_n501), .B2(new_n502), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n641), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n618), .A2(new_n460), .A3(new_n469), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT111), .B1(new_n820), .B2(new_n658), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n820), .A2(new_n658), .A3(KEYINPUT111), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n727), .B(new_n817), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT110), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n618), .A2(new_n460), .A3(new_n469), .A4(new_n636), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n611), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n611), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n704), .A2(new_n670), .B1(new_n720), .B2(new_n751), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n656), .A2(new_n666), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n670), .A2(new_n744), .A3(new_n688), .A4(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n669), .A2(new_n673), .A3(new_n670), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n673), .B1(new_n669), .B2(new_n670), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n830), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n675), .A2(KEYINPUT52), .A3(new_n830), .A4(new_n832), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n620), .A2(new_n501), .A3(new_n502), .A4(new_n665), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n643), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n751), .B1(new_n724), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n772), .B1(new_n842), .B2(new_n756), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n766), .A2(new_n762), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT104), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n766), .A2(new_n767), .A3(new_n762), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n843), .B1(new_n847), .B2(new_n764), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n839), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT112), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n611), .A2(new_n825), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT110), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n611), .A2(new_n824), .A3(new_n825), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n714), .A2(new_n718), .A3(new_n745), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n726), .B2(new_n723), .ZN(new_n856));
  INV_X1    g670(.A(new_n821), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n820), .A2(new_n658), .A3(KEYINPUT111), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n843), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n770), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT53), .A4(new_n839), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n829), .A2(new_n839), .A3(new_n848), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n850), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT54), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n871), .A3(new_n849), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n712), .A2(new_n754), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n664), .B1(new_n797), .B2(new_n800), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n761), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(KEYINPUT115), .A3(KEYINPUT48), .ZN(new_n877));
  XOR2_X1   g691(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n875), .B2(new_n761), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n688), .A2(new_n248), .A3(new_n664), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n748), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n741), .A2(new_n874), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n504), .B1(new_n883), .B2(new_n720), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n877), .A2(new_n879), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n712), .A2(new_n734), .A3(new_n740), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n382), .B1(new_n698), .B2(new_n699), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n874), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT50), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n886), .A2(KEYINPUT50), .A3(new_n874), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT113), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n875), .A2(new_n750), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n677), .A2(new_n634), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n881), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n897), .A3(new_n891), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n809), .A2(new_n810), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n608), .B1(new_n607), .B2(new_n232), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n613), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n472), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n754), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n883), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n899), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n885), .B1(new_n908), .B2(KEYINPUT51), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n896), .A2(KEYINPUT51), .A3(new_n892), .ZN(new_n910));
  INV_X1    g724(.A(new_n904), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n906), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT114), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT114), .B(new_n910), .C1(new_n911), .C2(new_n906), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n909), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n870), .A2(new_n872), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT116), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n870), .A2(new_n916), .A3(new_n919), .A4(new_n872), .ZN(new_n920));
  OR2_X1    g734(.A1(G952), .A2(G953), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n734), .A2(new_n461), .A3(new_n472), .A4(new_n793), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT109), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n902), .B(KEYINPUT49), .Z(new_n925));
  OR4_X1    g739(.A1(new_n700), .A2(new_n924), .A3(new_n688), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(G75));
  NOR2_X1   g741(.A1(new_n188), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n232), .B1(new_n868), .B2(new_n849), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT56), .B1(new_n930), .B2(G210), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n429), .A2(new_n435), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n441), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n443), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n931), .B2(new_n936), .ZN(G51));
  NAND2_X1  g752(.A1(new_n868), .A2(new_n849), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n871), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n595), .B(KEYINPUT57), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n607), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n784), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n930), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT117), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n928), .B1(new_n942), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  INV_X1    g761(.A(new_n545), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n928), .ZN(G60));
  INV_X1    g765(.A(new_n633), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n623), .B(KEYINPUT59), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n929), .B1(new_n940), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n870), .A2(new_n872), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n956), .B2(new_n953), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(G63));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(KEYINPUT118), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n928), .B1(KEYINPUT118), .B2(new_n959), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n939), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n962), .B1(new_n965), .B2(new_n653), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n230), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n970), .A2(new_n966), .A3(new_n960), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(G66));
  INV_X1    g786(.A(G224), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n507), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT119), .B1(new_n823), .B2(new_n828), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT119), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n854), .A2(new_n856), .A3(new_n859), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n974), .B1(new_n978), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n932), .B1(G898), .B2(new_n188), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  XNOR2_X1  g795(.A(new_n678), .B(KEYINPUT102), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n761), .A2(new_n982), .A3(new_n458), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n792), .A2(new_n983), .A3(new_n471), .A4(new_n692), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n806), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n772), .B(new_n830), .C1(new_n833), .C2(new_n834), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n770), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n814), .B2(new_n812), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n188), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n321), .B(KEYINPUT120), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(new_n541), .Z(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(G900), .B2(G953), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n992), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n701), .B(new_n830), .C1(new_n833), .C2(new_n834), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n748), .A2(new_n818), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n754), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n381), .A2(new_n999), .A3(new_n690), .A4(new_n692), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n806), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n675), .A2(new_n1002), .A3(new_n701), .A4(new_n830), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n997), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n815), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n995), .B1(new_n1005), .B2(new_n188), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n557), .B2(new_n662), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT121), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT122), .Z(new_n1009));
  NOR3_X1   g823(.A1(new_n994), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n990), .A2(new_n993), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1013), .A2(KEYINPUT123), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT123), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n990), .B2(new_n993), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1014), .A2(new_n1006), .A3(new_n1016), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1011), .B(new_n1012), .C1(new_n1017), .C2(new_n1008), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n994), .A2(new_n1015), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1006), .B1(new_n1013), .B2(KEYINPUT123), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1008), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT124), .B1(new_n1021), .B2(new_n1010), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1018), .A2(new_n1022), .ZN(G72));
  NOR2_X1   g837(.A1(new_n680), .A2(new_n314), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  AND3_X1   g841(.A1(new_n1025), .A2(new_n681), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1027), .B(KEYINPUT125), .Z(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n975), .A2(new_n977), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n1005), .ZN(new_n1032));
  INV_X1    g846(.A(new_n681), .ZN(new_n1033));
  AOI22_X1  g847(.A1(new_n869), .A2(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n763), .B1(new_n845), .B2(new_n846), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n806), .A2(new_n984), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1035), .A2(new_n986), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n810), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n471), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n813), .B1(new_n1040), .B2(new_n808), .ZN(new_n1041));
  INV_X1    g855(.A(new_n814), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1030), .B1(new_n1031), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(new_n1024), .ZN(new_n1045));
  AOI21_X1  g859(.A(KEYINPUT126), .B1(new_n1045), .B2(new_n929), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1029), .B1(new_n989), .B2(new_n978), .ZN(new_n1047));
  OAI211_X1 g861(.A(KEYINPUT126), .B(new_n929), .C1(new_n1047), .C2(new_n1025), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1034), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT127), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g866(.A(KEYINPUT127), .B(new_n1034), .C1(new_n1046), .C2(new_n1049), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(G57));
endmodule


