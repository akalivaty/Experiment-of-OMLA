//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n201), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n202), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n213), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n207), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(new_n203), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(G20), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n207), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n225), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G226), .B(G232), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT69), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n250), .B(new_n254), .Z(G351));
  NAND2_X1  g0055(.A1(new_n204), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT8), .A2(G58), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT70), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n256), .B1(new_n257), .B2(new_n259), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n229), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n267), .A2(new_n269), .B1(new_n201), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(new_n270), .B2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT9), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n282), .B1(G222), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n286), .B(new_n287), .C1(G77), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n287), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n290), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n289), .B(new_n293), .C1(new_n209), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n277), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT71), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT10), .A4(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n277), .A2(new_n301), .A3(new_n297), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n296), .A2(G179), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n296), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n276), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G97), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n215), .A2(G1698), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G226), .B2(G1698), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n314), .B2(new_n282), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n292), .B1(new_n315), .B2(new_n287), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n211), .B2(new_n295), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT14), .ZN(new_n320));
  INV_X1    g0120(.A(new_n318), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G179), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(new_n323), .A3(G169), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n210), .A2(G20), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n326), .B1(new_n201), .B2(new_n259), .C1(new_n327), .C2(new_n266), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n269), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT11), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT12), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n271), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n274), .A2(new_n331), .ZN(new_n333));
  INV_X1    g0133(.A(new_n326), .ZN(new_n334));
  INV_X1    g0134(.A(G13), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n331), .A2(new_n335), .A3(G1), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n333), .A2(G68), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n325), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n321), .A2(G190), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n318), .A2(G200), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n282), .B1(G232), .B2(new_n283), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n211), .B2(new_n283), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n287), .C1(G107), .C2(new_n288), .ZN(new_n346));
  INV_X1    g0146(.A(G244), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n346), .B(new_n293), .C1(new_n347), .C2(new_n295), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n348), .A2(G179), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT8), .B(G58), .Z(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n258), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n351), .B1(new_n265), .B2(new_n327), .C1(new_n266), .C2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n269), .B1(new_n327), .B2(new_n272), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n274), .A2(G77), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n348), .A2(new_n308), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n349), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OR4_X1    g0158(.A1(new_n311), .A2(new_n340), .A3(new_n343), .A4(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(KEYINPUT70), .A2(G58), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT70), .A2(G58), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n260), .B1(new_n362), .B2(KEYINPUT8), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n270), .A2(G20), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n269), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(KEYINPUT73), .A3(new_n364), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n271), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n264), .A2(new_n272), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n258), .A2(G159), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT65), .A2(G68), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT65), .A2(G68), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n362), .B1(new_n202), .B2(new_n203), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n373), .B1(new_n377), .B2(new_n265), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT72), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n278), .B2(G33), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n279), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n278), .A3(G33), .ZN(new_n382));
  AOI21_X1  g0182(.A(G20), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT72), .B1(new_n280), .B2(KEYINPUT3), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n265), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n203), .B1(new_n389), .B2(KEYINPUT7), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n368), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n288), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n265), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n210), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n393), .B1(new_n378), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n372), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n285), .A2(new_n283), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n382), .B(new_n400), .C1(new_n386), .C2(new_n387), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n283), .A2(G226), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT74), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT74), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n399), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n287), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n295), .A2(new_n215), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n292), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(G190), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n409), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G200), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n226), .B1(new_n210), .B2(new_n262), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n383), .B2(new_n384), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n389), .A2(KEYINPUT7), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n269), .B(new_n397), .C1(new_n418), .C2(new_n393), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n370), .A2(new_n371), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n412), .A2(new_n419), .A3(new_n420), .A4(new_n410), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G179), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n407), .A2(new_n425), .A3(new_n409), .ZN(new_n426));
  AOI21_X1  g0226(.A(G169), .B1(new_n407), .B2(new_n409), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT75), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n411), .A2(new_n308), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n407), .A2(new_n425), .A3(new_n409), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n398), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(KEYINPUT18), .A3(new_n434), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n424), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n348), .A2(G200), .ZN(new_n440));
  INV_X1    g0240(.A(new_n356), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n441), .C1(new_n300), .C2(new_n348), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n359), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT24), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n216), .A2(G20), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT22), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n279), .A3(new_n281), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT83), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n288), .A2(KEYINPUT83), .A3(new_n447), .A4(new_n446), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n265), .B(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT22), .B1(new_n453), .B2(new_n216), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(KEYINPUT78), .A2(G116), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT78), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n265), .A3(G33), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G20), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT23), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AND4_X1   g0263(.A1(new_n445), .A2(new_n455), .A3(new_n459), .A4(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n452), .B2(new_n454), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n445), .B1(new_n465), .B2(new_n459), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n269), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  XOR2_X1   g0267(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n468));
  NOR2_X1   g0268(.A1(new_n271), .A2(G107), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n270), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n271), .A2(new_n471), .A3(new_n229), .A4(new_n268), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G264), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n270), .A2(G45), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT5), .B(G41), .ZN(new_n478));
  AOI211_X1 g0278(.A(new_n475), .B(new_n287), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G294), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n217), .A2(new_n283), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n381), .A2(new_n382), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n283), .A2(G257), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n479), .B1(new_n484), .B2(new_n287), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n477), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G274), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(G190), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n488), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G200), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n467), .A2(new_n474), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(G169), .B1(new_n485), .B2(new_n488), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n280), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n279), .B2(new_n380), .ZN(new_n496));
  INV_X1    g0296(.A(new_n483), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n481), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n294), .B1(new_n498), .B2(new_n480), .ZN(new_n499));
  INV_X1    g0299(.A(new_n488), .ZN(new_n500));
  NOR4_X1   g0300(.A1(new_n499), .A2(new_n500), .A3(new_n479), .A4(G179), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n455), .A2(new_n459), .A3(new_n463), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT24), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n465), .A2(new_n445), .A3(new_n459), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n368), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n474), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n467), .A2(new_n474), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n502), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n493), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n496), .A2(new_n514), .A3(G257), .A4(new_n283), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n475), .A2(new_n283), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n382), .B(new_n516), .C1(new_n386), .C2(new_n387), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n282), .A2(G303), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G257), .B(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT81), .B1(new_n520), .B2(G1698), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n287), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n486), .A2(new_n294), .A3(G270), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n488), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(G20), .B1(new_n456), .B2(new_n457), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n265), .C1(G33), .C2(new_n221), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n269), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n527), .A2(KEYINPUT20), .A3(new_n269), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n272), .B1(new_n457), .B2(new_n456), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n472), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AND4_X1   g0338(.A1(KEYINPUT82), .A2(new_n534), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n532), .B2(new_n533), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT82), .B1(new_n540), .B2(new_n535), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n526), .B(G169), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(KEYINPUT82), .A3(new_n535), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n549), .A2(G179), .A3(new_n525), .A4(new_n523), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n526), .A2(G200), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n539), .A2(new_n541), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n523), .A2(G190), .A3(new_n525), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n549), .A2(KEYINPUT21), .A3(G169), .A4(new_n526), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n544), .A2(new_n550), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n288), .B2(G250), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n528), .C1(new_n559), .C2(new_n283), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT4), .B1(new_n496), .B2(G244), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n287), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n486), .A2(new_n294), .A3(G257), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n488), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT4), .B1(new_n282), .B2(new_n217), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G1698), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n558), .B1(new_n388), .B2(new_n347), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n557), .A4(new_n528), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n500), .B1(new_n569), .B2(new_n287), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(G190), .A3(new_n563), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n271), .A2(G97), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n288), .A2(new_n384), .A3(G20), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT7), .B1(new_n282), .B2(new_n265), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n258), .A2(KEYINPUT76), .A3(G77), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT76), .B1(new_n258), .B2(G77), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n460), .A2(KEYINPUT6), .A3(G97), .ZN(new_n578));
  AND2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n581), .B2(KEYINPUT6), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n577), .B1(new_n582), .B2(G20), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n575), .A2(new_n576), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n572), .B1(new_n584), .B2(new_n269), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n472), .A2(new_n221), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n565), .A2(new_n571), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n564), .A2(new_n308), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n570), .A2(new_n425), .A3(new_n563), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n269), .ZN(new_n591));
  INV_X1    g0391(.A(new_n572), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n587), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT80), .ZN(new_n595));
  INV_X1    g0395(.A(G200), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n458), .A2(G33), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n211), .A2(new_n283), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n382), .B(new_n598), .C1(new_n386), .C2(new_n387), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n283), .A2(G244), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n287), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT77), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n291), .B1(new_n603), .B2(new_n217), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n477), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n476), .A2(new_n603), .A3(G250), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n287), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n596), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n216), .A2(new_n221), .A3(new_n460), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n312), .A2(new_n265), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n312), .A2(KEYINPUT19), .A3(G20), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n453), .A2(new_n203), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n269), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n352), .A2(new_n272), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n472), .A2(new_n216), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n595), .B1(new_n609), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n602), .A2(G190), .A3(new_n608), .ZN(new_n621));
  INV_X1    g0421(.A(new_n600), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n381), .A2(new_n382), .A3(new_n622), .A4(new_n598), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n294), .B1(new_n623), .B2(new_n597), .ZN(new_n624));
  OAI21_X1  g0424(.A(G200), .B1(new_n624), .B2(new_n607), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n615), .A2(new_n269), .B1(new_n272), .B2(new_n352), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(KEYINPUT80), .A3(new_n626), .A4(new_n618), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n602), .A2(new_n425), .A3(new_n608), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT79), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n624), .A2(new_n607), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(KEYINPUT79), .A3(new_n425), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n308), .B1(new_n624), .B2(new_n607), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n472), .A2(new_n352), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n616), .A2(new_n617), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n631), .A2(new_n633), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n588), .A2(new_n594), .A3(new_n628), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n556), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n444), .A2(new_n513), .A3(new_n639), .ZN(G372));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n629), .A3(new_n634), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n621), .A2(new_n625), .A3(new_n626), .A4(new_n618), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n641), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n492), .A2(new_n594), .A3(new_n588), .A4(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n508), .A2(new_n544), .A3(new_n550), .A4(new_n555), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n628), .A2(new_n637), .ZN(new_n648));
  INV_X1    g0448(.A(new_n594), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(KEYINPUT86), .A3(KEYINPUT26), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n562), .A2(new_n488), .A3(new_n563), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n425), .B1(new_n585), .B2(new_n587), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n644), .A3(new_n589), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n628), .A2(new_n637), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n657), .A2(new_n655), .A3(new_n594), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n650), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n647), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n444), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n310), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n437), .A2(new_n438), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n341), .A2(new_n339), .A3(new_n342), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n340), .B1(new_n664), .B2(new_n358), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n665), .B2(new_n424), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n302), .A2(new_n306), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n544), .A2(new_n550), .A3(new_n555), .ZN(new_n670));
  XNOR2_X1  g0470(.A(KEYINPUT87), .B(KEYINPUT27), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n335), .A2(G20), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n671), .A2(new_n673), .A3(G1), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n671), .B1(new_n673), .B2(G1), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n552), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n670), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n556), .B2(new_n680), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n511), .B1(new_n510), .B2(new_n502), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n492), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n679), .B1(new_n467), .B2(new_n474), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n508), .B2(new_n679), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n670), .A2(new_n679), .ZN(new_n690));
  INV_X1    g0490(.A(new_n508), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n690), .A2(new_n513), .B1(new_n691), .B2(new_n679), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  NOR2_X1   g0493(.A1(new_n611), .A2(G116), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT88), .ZN(new_n695));
  INV_X1    g0495(.A(new_n232), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n695), .A2(new_n270), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n228), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND3_X1  g0500(.A1(new_n513), .A2(new_n639), .A3(new_n679), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n570), .A2(new_n485), .A3(new_n563), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n523), .A2(G179), .A3(new_n632), .A4(new_n525), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  OR3_X1    g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n632), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n564), .A2(new_n425), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n526), .A2(new_n490), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT89), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n704), .B1(new_n702), .B2(new_n703), .ZN(new_n710));
  AOI21_X1  g0510(.A(G179), .B1(new_n570), .B2(new_n563), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n523), .A2(new_n525), .B1(new_n485), .B2(new_n488), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT89), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .A4(new_n706), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n705), .A2(new_n709), .A3(new_n710), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n678), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n705), .B(new_n710), .C1(new_n707), .C2(new_n708), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n701), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n678), .B1(new_n647), .B2(new_n659), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(KEYINPUT90), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT90), .ZN(new_n725));
  AOI211_X1 g0525(.A(new_n725), .B(new_n678), .C1(new_n647), .C2(new_n659), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n724), .A2(new_n726), .A3(KEYINPUT29), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n657), .A2(new_n594), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n642), .B1(new_n730), .B2(new_n655), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n670), .B1(new_n509), .B2(new_n512), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n588), .A2(new_n594), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n492), .A3(new_n644), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n729), .B(new_n731), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n679), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT91), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT91), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n738), .A3(new_n679), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n728), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n722), .B1(new_n727), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n700), .B1(new_n742), .B2(G1), .ZN(G364));
  AOI21_X1  g0543(.A(new_n270), .B1(new_n672), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n697), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n683), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n682), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n250), .A2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT92), .ZN(new_n750));
  INV_X1    g0550(.A(G45), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n228), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n496), .A2(new_n696), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(new_n750), .C2(new_n749), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n288), .A2(G355), .A3(new_n232), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(G116), .C2(new_n232), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n229), .B1(G20), .B2(new_n308), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n746), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n265), .A2(G179), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n216), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n764), .A2(new_n300), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n282), .B(new_n766), .C1(G107), .C2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT96), .Z(new_n770));
  INV_X1    g0570(.A(KEYINPUT93), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n265), .B2(new_n425), .ZN(new_n772));
  NAND3_X1  g0572(.A1(KEYINPUT93), .A2(G20), .A3(G179), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G190), .A2(G200), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT94), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G77), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n764), .A2(new_n774), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  NAND3_X1  g0584(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n300), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(G190), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G50), .A2(new_n787), .B1(new_n788), .B2(G68), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n300), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n425), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n221), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n772), .A2(new_n790), .A3(new_n773), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n794), .B1(new_n362), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n780), .A2(new_n784), .A3(new_n789), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n767), .A2(new_n799), .B1(new_n781), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n775), .B1(new_n795), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n804), .C1(G294), .C2(new_n792), .ZN(new_n805));
  INV_X1    g0605(.A(G303), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n282), .B1(new_n765), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT97), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n787), .A2(G326), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n788), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI211_X1 g0611(.A(new_n805), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n807), .A2(new_n808), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n770), .A2(new_n798), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n763), .B1(new_n814), .B2(new_n760), .ZN(new_n815));
  INV_X1    g0615(.A(new_n759), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n762), .B(new_n815), .C1(new_n682), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n748), .A2(new_n817), .ZN(G396));
  OR2_X1    g0618(.A1(new_n723), .A2(KEYINPUT90), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n723), .A2(KEYINPUT90), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n356), .A2(new_n678), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n442), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n349), .A2(new_n356), .A3(new_n357), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n358), .A2(new_n679), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n819), .A2(new_n820), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n826), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n723), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n722), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n763), .ZN(new_n833));
  INV_X1    g0633(.A(new_n760), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n793), .A2(new_n262), .B1(new_n767), .B2(new_n203), .ZN(new_n835));
  INV_X1    g0635(.A(new_n781), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n388), .B(new_n835), .C1(G132), .C2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G137), .A2(new_n787), .B1(new_n788), .B2(G150), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  INV_X1    g0639(.A(G143), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n840), .B2(new_n795), .C1(new_n782), .C2(new_n778), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n841), .A2(KEYINPUT34), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(KEYINPUT34), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n837), .B1(new_n201), .B2(new_n765), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n787), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n799), .A2(new_n810), .B1(new_n845), .B2(new_n806), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n794), .ZN(new_n847));
  INV_X1    g0647(.A(new_n765), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G107), .B1(new_n768), .B2(G87), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n802), .B2(new_n781), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G294), .B2(new_n796), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n779), .A2(new_n458), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n847), .A2(new_n851), .A3(new_n282), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n834), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n763), .B(new_n854), .C1(new_n757), .C2(new_n826), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n760), .A2(new_n757), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(G77), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n833), .A2(new_n858), .ZN(G384));
  OAI211_X1 g0659(.A(G20), .B(new_n230), .C1(new_n582), .C2(KEYINPUT35), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n536), .B(new_n860), .C1(KEYINPUT35), .C2(new_n582), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT36), .Z(new_n862));
  NAND2_X1  g0662(.A1(G50), .A2(G58), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n270), .B1(new_n863), .B2(new_n203), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n327), .B1(new_n376), .B2(new_n362), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n335), .B(new_n864), .C1(new_n865), .C2(new_n201), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT99), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n340), .A2(new_n679), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT102), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT39), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  INV_X1    g0674(.A(new_n676), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n434), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n435), .A2(new_n874), .A3(new_n421), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n269), .B1(new_n418), .B2(new_n393), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n391), .A2(KEYINPUT16), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n420), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n875), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n421), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n418), .A2(new_n393), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n372), .B1(new_n392), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n428), .B2(new_n432), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n421), .A2(new_n422), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n421), .A2(new_n422), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n436), .B(new_n398), .C1(new_n428), .C2(new_n432), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT18), .B1(new_n433), .B2(new_n434), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n881), .ZN(new_n893));
  AOI221_X4 g0693(.A(new_n873), .B1(new_n877), .B2(new_n886), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n877), .A2(new_n886), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT103), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n424), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n413), .A2(new_n423), .A3(KEYINPUT103), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n900), .B(new_n901), .C1(new_n891), .C2(new_n890), .ZN(new_n902));
  INV_X1    g0702(.A(new_n876), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n435), .A2(new_n421), .A3(new_n876), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n902), .A2(new_n903), .B1(new_n877), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT104), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n872), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n901), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT103), .B1(new_n413), .B2(new_n423), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n876), .B1(new_n911), .B2(new_n663), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n905), .A2(new_n877), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n873), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n915));
  NOR2_X1   g0715(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n871), .B1(new_n908), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n338), .A2(new_n678), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n664), .B(new_n919), .C1(new_n325), .C2(new_n339), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n338), .B(new_n678), .C1(new_n343), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n678), .B(new_n826), .C1(new_n647), .C2(new_n659), .ZN(new_n925));
  INV_X1    g0725(.A(new_n825), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT100), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT100), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n829), .A2(new_n928), .A3(new_n825), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n924), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT101), .B1(new_n894), .B2(new_n897), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n896), .B1(new_n439), .B2(new_n881), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n873), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT101), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n915), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n437), .A2(new_n438), .A3(new_n676), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n918), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n819), .A2(new_n728), .A3(new_n820), .ZN(new_n939));
  INV_X1    g0739(.A(new_n739), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n738), .B1(new_n735), .B2(new_n679), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT29), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n444), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n668), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n938), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n923), .A2(new_n828), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n701), .A2(new_n718), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT105), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT105), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n701), .A2(new_n718), .A3(new_n950), .A4(new_n947), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n946), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n931), .A2(new_n952), .A3(new_n935), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n914), .B2(new_n915), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n953), .A2(new_n954), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n949), .A2(new_n951), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n444), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(G330), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n945), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n672), .A2(new_n270), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n868), .B1(new_n961), .B2(new_n962), .ZN(G367));
  NAND2_X1  g0763(.A1(new_n593), .A2(new_n678), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n733), .A2(new_n509), .A3(new_n512), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n678), .B1(new_n965), .B2(new_n594), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n690), .A2(new_n513), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n733), .A2(new_n964), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT42), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT109), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n619), .A2(new_n678), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n644), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n641), .A2(new_n976), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT106), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT43), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n974), .A2(new_n975), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT109), .B1(new_n973), .B2(new_n983), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n973), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n649), .A2(new_n678), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n968), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n683), .A2(new_n688), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT108), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n985), .A2(new_n986), .A3(new_n993), .A4(new_n988), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT111), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n689), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT44), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n692), .B2(new_n991), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n691), .A2(new_n679), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n670), .A2(new_n679), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n686), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n991), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(KEYINPUT44), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1001), .A2(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n683), .A2(KEYINPUT111), .A3(new_n688), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n999), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1014));
  AND4_X1   g0814(.A1(new_n999), .A2(new_n1013), .A3(new_n1014), .A4(new_n1011), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n967), .B1(new_n688), .B2(new_n690), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(new_n683), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n742), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT112), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n697), .B(new_n1021), .Z(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1024), .A2(new_n998), .A3(new_n689), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1010), .A2(new_n999), .A3(new_n1011), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1018), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n741), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1022), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT112), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1023), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n997), .B1(new_n1032), .B2(new_n744), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n848), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n768), .A2(G97), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n460), .B2(new_n793), .C1(new_n845), .C2(new_n802), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(G294), .C2(new_n788), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT46), .B1(new_n848), .B2(new_n458), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n496), .B(new_n1038), .C1(G303), .C2(new_n796), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(new_n799), .C2(new_n778), .ZN(new_n1040));
  INV_X1    g0840(.A(G317), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n781), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(G137), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n781), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n793), .A2(new_n203), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n795), .A2(new_n257), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n767), .A2(new_n327), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n288), .B1(new_n765), .B2(new_n262), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G143), .A2(new_n787), .B1(new_n788), .B2(G159), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n201), .C2(new_n778), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1040), .A2(new_n1042), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT47), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n763), .B1(new_n1053), .B2(new_n760), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n753), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n761), .B1(new_n232), .B2(new_n352), .C1(new_n1055), .C2(new_n245), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n982), .A2(new_n816), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT113), .B1(new_n1033), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n745), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1058), .C1(new_n1062), .C2(new_n997), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(G387));
  AOI22_X1  g0864(.A1(G311), .A2(new_n788), .B1(new_n787), .B2(G322), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n1041), .B2(new_n795), .C1(new_n806), .C2(new_n778), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n848), .A2(G294), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n792), .A2(G283), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n836), .A2(G326), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n496), .B1(new_n458), .B2(new_n768), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n775), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G50), .A2(new_n796), .B1(new_n1079), .B2(G68), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n352), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n792), .A2(new_n1081), .ZN(new_n1082));
  AND4_X1   g0882(.A1(new_n496), .A2(new_n1080), .A3(new_n1035), .A4(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G159), .A2(new_n787), .B1(new_n788), .B2(new_n363), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n765), .A2(new_n327), .B1(new_n781), .B2(new_n257), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT114), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1078), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n763), .B1(new_n1088), .B2(new_n760), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n350), .A2(new_n201), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT50), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n203), .A2(new_n327), .ZN(new_n1092));
  NOR4_X1   g0892(.A1(new_n1091), .A2(G45), .A3(new_n695), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n753), .B1(new_n242), .B2(new_n751), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n695), .A2(new_n232), .A3(new_n288), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n232), .A2(G107), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n761), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1089), .B(new_n1098), .C1(new_n688), .C2(new_n816), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT117), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n697), .B1(new_n742), .B2(new_n1028), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n741), .A2(new_n1018), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1100), .B1(new_n744), .B2(new_n1018), .C1(new_n1101), .C2(new_n1102), .ZN(G393));
  NOR2_X1   g0903(.A1(new_n810), .A2(new_n806), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G283), .A2(new_n848), .B1(new_n792), .B2(new_n458), .ZN(new_n1105));
  INV_X1    g0905(.A(G294), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n775), .C1(new_n803), .C2(new_n781), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT52), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n845), .A2(new_n1041), .B1(new_n802), .B2(new_n795), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1104), .B(new_n1107), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n288), .B1(new_n768), .B2(G107), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT119), .Z(new_n1113));
  AOI22_X1  g0913(.A1(new_n779), .A2(new_n350), .B1(G50), .B2(new_n788), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n327), .B2(new_n793), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT118), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n787), .A2(G150), .B1(new_n796), .B2(G159), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n496), .B1(new_n216), .B2(new_n767), .C1(new_n840), .C2(new_n781), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1116), .B(new_n1121), .C1(new_n210), .C2(new_n765), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n763), .B1(new_n1123), .B2(new_n760), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n761), .B1(new_n221), .B2(new_n232), .C1(new_n254), .C2(new_n1055), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n816), .C2(new_n991), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1016), .B2(new_n744), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n697), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1102), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n1016), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1102), .A2(new_n1027), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1127), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G390));
  NAND3_X1  g0933(.A1(new_n444), .A2(G330), .A3(new_n957), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n943), .A2(new_n1134), .A3(new_n668), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n824), .A2(new_n825), .A3(G330), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n949), .B2(new_n951), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n923), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n721), .A2(new_n1136), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n924), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n927), .A2(new_n929), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1138), .A2(new_n923), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1140), .A2(new_n924), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n737), .A2(new_n739), .A3(new_n825), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n824), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1135), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT104), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n902), .A2(new_n903), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n905), .A2(new_n877), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n1154), .B2(new_n873), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n933), .A2(new_n915), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT39), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n930), .C2(new_n871), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1147), .A2(new_n824), .A3(new_n923), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n914), .A2(new_n915), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n870), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1159), .A2(new_n1162), .A3(new_n1146), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1139), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1150), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1165), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1135), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1159), .A2(new_n1162), .A3(new_n1146), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1166), .A2(new_n1172), .A3(new_n697), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n745), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1157), .A2(new_n757), .A3(new_n1158), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n787), .A2(G128), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n282), .B1(new_n792), .B2(G159), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n201), .C2(new_n767), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G137), .B2(new_n788), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n836), .A2(G125), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT54), .B(G143), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n779), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n848), .A2(G150), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1184), .A2(KEYINPUT53), .B1(new_n796), .B2(G132), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1184), .A2(KEYINPUT53), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G68), .A2(new_n768), .B1(new_n792), .B2(G77), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n796), .A2(G116), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n836), .A2(G294), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1188), .A2(new_n282), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G107), .A2(new_n788), .B1(new_n787), .B2(G283), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n216), .B2(new_n765), .C1(new_n221), .C2(new_n778), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1186), .A2(new_n1187), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT120), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n763), .B1(new_n1195), .B2(new_n760), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1176), .B(new_n1196), .C1(new_n363), .C2(new_n857), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1173), .A2(new_n1175), .A3(new_n1197), .ZN(G378));
  NAND2_X1  g0998(.A1(new_n953), .A2(new_n954), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n955), .A2(new_n952), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n311), .B(KEYINPUT55), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n276), .A2(new_n875), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT56), .Z(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AND4_X1   g1008(.A1(G330), .A2(new_n1199), .A3(new_n1200), .A4(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n956), .B2(G330), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n938), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1199), .A2(G330), .A3(new_n1200), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1208), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n918), .A2(new_n936), .A3(new_n937), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n956), .A2(G330), .A3(new_n1208), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT123), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1211), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1220));
  OAI211_X1 g1020(.A(KEYINPUT123), .B(new_n938), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1169), .A2(new_n1166), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1128), .B1(new_n1225), .B2(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1219), .A2(new_n1221), .A3(new_n745), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1205), .A2(new_n757), .A3(new_n1206), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n768), .A2(new_n362), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n327), .B2(new_n765), .C1(new_n799), .C2(new_n781), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1231), .A2(G41), .A3(new_n496), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT121), .Z(new_n1233));
  OAI22_X1  g1033(.A1(new_n221), .A2(new_n810), .B1(new_n845), .B2(new_n536), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1045), .B(new_n1234), .C1(new_n1081), .C2(new_n1079), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(new_n460), .C2(new_n795), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT58), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n792), .A2(G150), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G125), .A2(new_n787), .B1(new_n788), .B2(G132), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1079), .A2(G137), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n796), .A2(G128), .B1(new_n848), .B2(new_n1182), .ZN(new_n1241));
  AND4_X1   g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT59), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G41), .B1(new_n768), .B2(G159), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G33), .B1(new_n836), .B2(G124), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G41), .B1(new_n496), .B2(G33), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1237), .B(new_n1246), .C1(G50), .C2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n763), .B1(new_n1248), .B2(new_n760), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1229), .B(new_n1249), .C1(G50), .C2(new_n857), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1228), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1227), .A2(new_n1251), .ZN(G375));
  NAND3_X1  g1052(.A1(new_n1135), .A2(new_n1144), .A3(new_n1149), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1170), .A2(new_n1022), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n856), .A2(new_n203), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n845), .A2(new_n1106), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1047), .B(new_n1256), .C1(new_n458), .C2(new_n788), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1082), .B1(new_n221), .B2(new_n765), .C1(new_n806), .C2(new_n781), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G283), .B2(new_n796), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n779), .A2(G107), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1257), .A2(new_n282), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n788), .A2(new_n1182), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n1230), .C1(new_n782), .C2(new_n765), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G132), .B2(new_n787), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n496), .B1(new_n795), .B2(new_n1043), .C1(new_n257), .C2(new_n775), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G128), .B2(new_n836), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(new_n201), .C2(new_n793), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n834), .B1(new_n1261), .B2(new_n1267), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n763), .B(new_n1268), .C1(new_n924), .C2(new_n757), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1168), .A2(new_n745), .B1(new_n1255), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1254), .A2(new_n1270), .ZN(G381));
  NOR2_X1   g1071(.A1(G375), .A2(G378), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(G381), .A2(G384), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1060), .A2(new_n1063), .A3(new_n1132), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1274), .A2(G396), .A3(G393), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1275), .ZN(G407));
  AOI21_X1  g1076(.A(new_n677), .B1(new_n1275), .B2(new_n1273), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1272), .ZN(new_n1278));
  OAI21_X1  g1078(.A(G213), .B1(new_n1277), .B2(new_n1278), .ZN(G409));
  NAND3_X1  g1079(.A1(new_n1227), .A2(G378), .A3(new_n1251), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1211), .A2(new_n1217), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n745), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1250), .B(new_n1282), .C1(new_n1222), .C2(new_n1030), .ZN(new_n1283));
  INV_X1    g1083(.A(G378), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1280), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(G213), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(G343), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(G2897), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT124), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1135), .A2(new_n1144), .A3(KEYINPUT60), .A4(new_n1149), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1170), .A2(new_n1294), .A3(new_n697), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1253), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1270), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G384), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1293), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1253), .A2(new_n1296), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1301), .A2(new_n697), .A3(new_n1170), .A4(new_n1294), .ZN(new_n1302));
  AOI211_X1 g1102(.A(KEYINPUT124), .B(G384), .C1(new_n1302), .C2(new_n1270), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(G384), .A3(new_n1270), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1292), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1305), .ZN(new_n1307));
  NOR4_X1   g1107(.A1(new_n1300), .A2(new_n1303), .A3(new_n1307), .A4(new_n1291), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1288), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1311), .B(new_n1313), .C1(new_n1314), .C2(KEYINPUT63), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1286), .A2(new_n1289), .A3(new_n1313), .ZN(new_n1316));
  XOR2_X1   g1116(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1310), .A2(new_n1315), .A3(new_n1318), .ZN(new_n1319));
  XOR2_X1   g1119(.A(G393), .B(G396), .Z(new_n1320));
  OAI21_X1  g1120(.A(G390), .B1(new_n1033), .B2(new_n1059), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1058), .B(new_n1132), .C1(new_n1062), .C2(new_n997), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1274), .A2(new_n1321), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1320), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  AOI211_X1 g1127(.A(KEYINPUT126), .B(new_n1320), .C1(new_n1274), .C2(new_n1321), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1323), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  AND4_X1   g1130(.A1(new_n1330), .A2(new_n1286), .A3(new_n1289), .A4(new_n1313), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1334), .B1(new_n1311), .B2(new_n1335), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1336), .A2(new_n1329), .ZN(new_n1337));
  AOI22_X1  g1137(.A1(new_n1319), .A2(new_n1329), .B1(new_n1333), .B2(new_n1337), .ZN(G405));
  INV_X1    g1138(.A(new_n1280), .ZN(new_n1339));
  AOI21_X1  g1139(.A(G378), .B1(new_n1227), .B2(new_n1251), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1313), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1340), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1342), .A2(new_n1280), .A3(new_n1312), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(new_n1329), .ZN(G402));
endmodule


