//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT95), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(new_n204), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(G43gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(G43gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n213), .B(KEYINPUT93), .Z(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT94), .B(G50gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G43gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G29gat), .A2(G36gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT14), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n220), .A2(KEYINPUT14), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT92), .B(G29gat), .ZN(new_n223));
  AOI211_X1 g022(.A(new_n221), .B(new_n222), .C1(G36gat), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n214), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n214), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n210), .A2(new_n227), .ZN(new_n228));
  OR3_X1    g027(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT17), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n210), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT96), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(G169gat), .B(G197gat), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT12), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n232), .A2(KEYINPUT18), .A3(new_n235), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n210), .B(new_n227), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n234), .B(KEYINPUT13), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT98), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT98), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n244), .A4(new_n238), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT97), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n246), .A2(KEYINPUT97), .A3(new_n249), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n238), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n244), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n251), .A2(new_n254), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT35), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g061(.A1(G211gat), .A2(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G197gat), .A2(G204gat), .ZN(new_n266));
  AND2_X1   g065(.A1(G197gat), .A2(G204gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(KEYINPUT77), .A3(new_n263), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273));
  AND2_X1   g072(.A1(G211gat), .A2(G218gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(G211gat), .A2(G218gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n268), .A2(new_n272), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n268), .A2(new_n272), .A3(new_n276), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n274), .A2(new_n275), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT78), .B1(new_n268), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n262), .B1(new_n282), .B2(KEYINPUT29), .ZN(new_n283));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  INV_X1    g083(.A(G155gat), .ZN(new_n285));
  INV_X1    g084(.A(G162gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G141gat), .B(G148gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n284), .B(new_n287), .C1(new_n288), .C2(KEYINPUT2), .ZN(new_n289));
  INV_X1    g088(.A(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G148gat), .ZN(new_n291));
  INV_X1    g090(.A(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G141gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n284), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n284), .A2(KEYINPUT2), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n289), .A2(new_n262), .A3(new_n297), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(KEYINPUT83), .A3(new_n301), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n282), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G228gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n282), .ZN(new_n310));
  OAI221_X1 g109(.A(new_n265), .B1(new_n274), .B2(new_n275), .C1(new_n266), .C2(new_n267), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n268), .A2(new_n280), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT29), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n298), .B1(new_n313), .B2(KEYINPUT3), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n308), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT82), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317));
  AOI211_X1 g116(.A(new_n317), .B(new_n308), .C1(new_n310), .C2(new_n314), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n309), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G22gat), .ZN(new_n320));
  INV_X1    g119(.A(G22gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n321), .B(new_n309), .C1(new_n316), .C2(new_n318), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT31), .B(G50gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  AND2_X1   g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n319), .B2(G22gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n315), .B(KEYINPUT82), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n329), .A2(KEYINPUT84), .A3(new_n321), .A4(new_n309), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n328), .A2(new_n330), .A3(new_n332), .A4(KEYINPUT85), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n327), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G113gat), .ZN(new_n338));
  INV_X1    g137(.A(G120gat), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT1), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n338), .B2(new_n339), .ZN(new_n341));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344));
  AND2_X1   g143(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n340), .B(new_n344), .C1(new_n347), .C2(new_n338), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(KEYINPUT23), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n353), .A2(G169gat), .A3(G176gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT65), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT64), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT64), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(G183gat), .ZN(new_n362));
  INV_X1    g161(.A(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n357), .A2(new_n359), .A3(new_n361), .A4(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT23), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT65), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n353), .B1(G169gat), .B2(G176gat), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n350), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n355), .A2(new_n365), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n350), .A3(new_n369), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n358), .A2(KEYINPUT67), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT67), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n356), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(KEYINPUT69), .A2(G190gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(KEYINPUT69), .A2(G190gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n382), .A2(new_n385), .B1(new_n377), .B2(new_n356), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n372), .B1(new_n379), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n371), .B1(new_n387), .B2(new_n366), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n351), .A2(KEYINPUT26), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(new_n362), .B2(new_n363), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n350), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n351), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT27), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT70), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n399), .A3(G183gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT68), .B(G183gat), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n400), .B(new_n382), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT28), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT27), .B(G183gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n405), .A3(KEYINPUT28), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n395), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n349), .B1(new_n388), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G227gat), .ZN(new_n409));
  INV_X1    g208(.A(G233gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT69), .B(G190gat), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(KEYINPUT27), .B2(new_n385), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT28), .B1(new_n413), .B2(new_n400), .ZN(new_n414));
  INV_X1    g213(.A(new_n406), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n394), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n343), .A2(new_n348), .ZN(new_n417));
  INV_X1    g216(.A(new_n372), .ZN(new_n418));
  OAI22_X1  g217(.A1(new_n412), .A2(new_n401), .B1(new_n357), .B2(KEYINPUT66), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n373), .B(new_n375), .C1(new_n377), .C2(new_n356), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT25), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n416), .A2(new_n417), .A3(new_n422), .A4(new_n371), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n411), .A3(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G71gat), .B(G99gat), .Z(new_n425));
  XNOR2_X1  g224(.A(G15gat), .B(G43gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT33), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT72), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(KEYINPUT32), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n408), .A2(new_n423), .A3(new_n411), .A4(new_n427), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n432), .B2(new_n428), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n411), .B1(new_n408), .B2(new_n423), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT34), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI211_X1 g237(.A(KEYINPUT34), .B(new_n411), .C1(new_n408), .C2(new_n423), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT74), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n435), .A2(new_n442), .A3(new_n440), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n435), .B2(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n337), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n343), .A2(new_n348), .A3(new_n289), .A4(new_n297), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n348), .A2(new_n343), .B1(new_n289), .B2(new_n297), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n289), .A4(new_n297), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n300), .A3(new_n417), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n454), .A2(new_n456), .A3(new_n447), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT0), .ZN(new_n462));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT4), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n465), .A2(KEYINPUT5), .A3(new_n447), .A4(new_n456), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n460), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n460), .B2(new_n466), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT6), .ZN(new_n469));
  AND4_X1   g268(.A1(KEYINPUT6), .A2(new_n460), .A3(new_n464), .A4(new_n466), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT79), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n301), .B1(new_n388), .B2(new_n407), .ZN(new_n473));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n355), .A2(new_n370), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n365), .A2(new_n366), .ZN(new_n477));
  AOI22_X1  g276(.A1(KEYINPUT25), .A2(new_n421), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n478), .B2(new_n416), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n472), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT79), .B1(new_n473), .B2(new_n474), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n282), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT29), .B1(new_n478), .B2(new_n416), .ZN(new_n484));
  INV_X1    g283(.A(new_n474), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT80), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n473), .A2(new_n487), .A3(new_n474), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n479), .A2(new_n282), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT81), .A4(new_n488), .ZN(new_n493));
  XNOR2_X1  g292(.A(G8gat), .B(G36gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(G64gat), .B(G92gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n494), .B(new_n495), .Z(new_n496));
  NAND4_X1  g295(.A1(new_n483), .A2(new_n492), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n492), .A3(new_n493), .ZN(new_n500));
  INV_X1    g299(.A(new_n496), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n498), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n483), .A2(new_n492), .A3(new_n493), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT86), .A4(new_n504), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n471), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n261), .B(new_n446), .C1(new_n509), .C2(KEYINPUT89), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n435), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n440), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT73), .B(new_n431), .C1(new_n433), .C2(new_n434), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n444), .B2(new_n443), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n337), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n505), .A2(new_n471), .ZN(new_n519));
  AOI211_X1 g318(.A(KEYINPUT90), .B(new_n261), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n335), .A2(new_n336), .ZN(new_n522));
  INV_X1    g321(.A(new_n327), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n525));
  INV_X1    g324(.A(new_n471), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n435), .A2(new_n440), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n435), .A2(new_n442), .A3(new_n440), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n440), .B1(new_n435), .B2(new_n512), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n515), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n521), .B1(new_n532), .B2(KEYINPUT35), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n510), .A2(new_n511), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n524), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n445), .A2(KEYINPUT76), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n516), .B(KEYINPUT36), .C1(new_n444), .C2(new_n443), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n445), .A2(new_n537), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n535), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n471), .A2(new_n497), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n501), .A2(KEYINPUT37), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n502), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n486), .A2(new_n488), .ZN(new_n550));
  INV_X1    g349(.A(new_n282), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n479), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n481), .B2(new_n482), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT38), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n546), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n500), .A2(KEYINPUT37), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n501), .B1(new_n500), .B2(KEYINPUT37), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT38), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n337), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n464), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n465), .A2(new_n456), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n448), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n563), .B2(KEYINPUT39), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n450), .A2(new_n451), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT39), .B1(new_n565), .B2(new_n448), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n562), .B2(new_n448), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT87), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(KEYINPUT40), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n467), .B1(new_n568), .B2(KEYINPUT40), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n507), .A2(new_n571), .A3(new_n508), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT88), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n560), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n560), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n545), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n260), .B1(new_n534), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT21), .ZN(new_n578));
  XOR2_X1   g377(.A(G57gat), .B(G64gat), .Z(new_n579));
  INV_X1    g378(.A(KEYINPUT9), .ZN(new_n580));
  INV_X1    g379(.A(G71gat), .ZN(new_n581));
  INV_X1    g380(.A(G78gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(KEYINPUT99), .A3(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n210), .B1(new_n578), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT101), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G127gat), .B(G155gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n588), .A2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n595), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n231), .A2(new_n229), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n615), .B(new_n617), .C1(new_n227), .C2(new_n614), .ZN(new_n618));
  XOR2_X1   g417(.A(G190gat), .B(G218gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n613), .B(new_n586), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR3_X1    g429(.A1(new_n614), .A2(new_n629), .A3(new_n586), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n628), .B2(new_n633), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n604), .A2(new_n627), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n577), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n526), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT102), .B(G1gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1324gat));
  NAND2_X1  g448(.A1(new_n507), .A2(new_n508), .ZN(new_n650));
  OAI21_X1  g449(.A(G8gat), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n507), .A2(new_n508), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT16), .B(G8gat), .Z(new_n654));
  NAND4_X1  g453(.A1(new_n577), .A2(new_n653), .A3(new_n645), .A4(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n655), .A2(KEYINPUT103), .A3(new_n652), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT103), .B1(new_n655), .B2(new_n652), .ZN(new_n657));
  OAI221_X1 g456(.A(new_n651), .B1(new_n652), .B2(new_n655), .C1(new_n656), .C2(new_n657), .ZN(G1325gat));
  AOI21_X1  g457(.A(KEYINPUT76), .B1(new_n445), .B2(new_n537), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT104), .B1(new_n540), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n544), .A2(new_n661), .A3(new_n539), .A4(new_n538), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G15gat), .B1(new_n646), .B2(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n445), .A2(G15gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n646), .B2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n646), .A2(new_n524), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n604), .A2(new_n642), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n627), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n577), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(new_n526), .A3(new_n223), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n671), .A2(new_n260), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n534), .A2(new_n576), .ZN(new_n679));
  INV_X1    g478(.A(new_n627), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n560), .A2(new_n572), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n560), .A2(new_n572), .A3(new_n573), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n535), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n663), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n534), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n627), .A2(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n678), .B1(new_n682), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n223), .B1(new_n693), .B2(new_n526), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n694), .ZN(G1328gat));
  INV_X1    g494(.A(new_n673), .ZN(new_n696));
  AOI21_X1  g495(.A(G36gat), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n653), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G36gat), .B1(new_n693), .B2(new_n650), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n663), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G43gat), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n445), .A2(G43gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n577), .A2(new_n672), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n706), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n705), .B(new_n712), .C1(new_n708), .C2(G43gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(G1330gat));
  INV_X1    g515(.A(new_n217), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n673), .A2(new_n524), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n679), .B2(new_n680), .ZN(new_n720));
  INV_X1    g519(.A(new_n690), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n688), .B2(new_n534), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n337), .B(new_n677), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n718), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n724), .A2(KEYINPUT108), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n724), .B2(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1331gat));
  INV_X1    g528(.A(new_n260), .ZN(new_n730));
  INV_X1    g529(.A(new_n604), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n730), .A2(new_n731), .A3(new_n680), .A4(new_n643), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n689), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n471), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g535(.A(new_n650), .B(KEYINPUT110), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  NOR3_X1   g542(.A1(new_n733), .A2(G71gat), .A3(new_n445), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n707), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(G71gat), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n733), .A2(new_n524), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n582), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n730), .A2(new_n604), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n642), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n682), .B2(new_n691), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n608), .B1(new_n752), .B2(new_n471), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n535), .B1(new_n684), .B2(new_n685), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT89), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n653), .B2(new_n471), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n757), .A2(new_n261), .A3(new_n758), .A4(new_n446), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT90), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n532), .A2(new_n521), .A3(KEYINPUT35), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n755), .A2(new_n663), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n750), .A2(new_n680), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n754), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n765), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n689), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n643), .A2(G85gat), .A3(new_n526), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n753), .A2(new_n771), .A3(KEYINPUT111), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT111), .B1(new_n753), .B2(new_n771), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1336gat));
  INV_X1    g573(.A(new_n751), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n653), .B(new_n775), .C1(new_n720), .C2(new_n722), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n776), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT112), .B1(new_n776), .B2(G92gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n765), .B1(new_n688), .B2(new_n534), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n754), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n764), .C2(new_n765), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n738), .A2(G92gat), .A3(new_n643), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n777), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(new_n769), .B2(new_n783), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n737), .B(new_n775), .C1(new_n720), .C2(new_n722), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G92gat), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n787), .B2(new_n790), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n785), .A2(new_n786), .B1(new_n791), .B2(new_n792), .ZN(G1337gat));
  NAND2_X1  g592(.A1(new_n752), .A2(new_n707), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G99gat), .ZN(new_n795));
  INV_X1    g594(.A(new_n769), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n643), .A2(new_n445), .A3(G99gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT115), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(G1338gat));
  NAND2_X1  g598(.A1(new_n752), .A2(new_n337), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n524), .A2(new_n643), .A3(G106gat), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT116), .Z(new_n803));
  AOI21_X1  g602(.A(KEYINPUT53), .B1(new_n769), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n781), .A2(new_n782), .ZN(new_n806));
  AOI22_X1  g605(.A1(G106gat), .A2(new_n800), .B1(new_n806), .B2(new_n803), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G1339gat));
  OAI21_X1  g608(.A(new_n639), .B1(new_n634), .B2(KEYINPUT54), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n632), .A2(KEYINPUT117), .A3(new_n633), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT117), .B1(new_n632), .B2(new_n633), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n630), .A2(new_n631), .B1(G230gat), .B2(G233gat), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n810), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT55), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n640), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n254), .A2(new_n251), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n817), .A2(KEYINPUT55), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n247), .A2(new_n248), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT118), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n232), .A2(new_n235), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n243), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n604), .B1(new_n826), .B2(new_n680), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(new_n642), .A3(new_n825), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n819), .A2(new_n821), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n627), .B(new_n828), .C1(new_n829), .C2(new_n260), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n827), .A2(new_n830), .B1(new_n260), .B2(new_n645), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n337), .A3(new_n445), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n738), .A2(new_n471), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(new_n338), .A3(new_n260), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n831), .A2(new_n526), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n518), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n737), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n730), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n338), .B2(new_n840), .ZN(G1340gat));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n347), .A3(new_n642), .ZN(new_n842));
  OAI21_X1  g641(.A(G120gat), .B1(new_n835), .B2(new_n643), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n845), .A3(new_n604), .ZN(new_n846));
  OAI21_X1  g645(.A(G127gat), .B1(new_n835), .B2(new_n731), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  NAND2_X1  g647(.A1(new_n680), .A2(new_n650), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n838), .A2(G134gat), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n835), .B2(new_n627), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n707), .A2(new_n524), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n737), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n290), .A3(new_n730), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n827), .A2(new_n830), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n645), .A2(new_n260), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n337), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT57), .B1(new_n831), .B2(new_n524), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n833), .A2(new_n707), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n864), .A2(new_n260), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n857), .B1(new_n290), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1344gat));
  NAND3_X1  g669(.A1(new_n856), .A2(new_n292), .A3(new_n642), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  OR3_X1    g671(.A1(new_n524), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n860), .A2(new_n873), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n874), .A2(new_n642), .A3(new_n865), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n872), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n864), .A2(new_n643), .A3(new_n866), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(KEYINPUT59), .A3(new_n292), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n871), .B1(new_n878), .B2(new_n880), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n856), .A2(new_n285), .A3(new_n604), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n864), .A2(new_n731), .A3(new_n866), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n285), .ZN(G1346gat));
  OR3_X1    g683(.A1(new_n855), .A2(G162gat), .A3(new_n849), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n864), .A2(new_n627), .A3(new_n866), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n286), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT121), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n650), .A2(new_n471), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n832), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n260), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT124), .Z(new_n892));
  OR3_X1    g691(.A1(new_n831), .A2(KEYINPUT122), .A3(new_n471), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT122), .B1(new_n831), .B2(new_n471), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n738), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n518), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT123), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n898), .A3(new_n518), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n260), .A2(G169gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n892), .A2(new_n901), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n643), .A2(G176gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G176gat), .B1(new_n890), .B2(new_n643), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1349gat));
  OAI21_X1  g705(.A(KEYINPUT125), .B1(new_n890), .B2(new_n731), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n832), .A2(new_n908), .A3(new_n604), .A4(new_n889), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n401), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n405), .A3(new_n518), .A4(new_n604), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1350gat));
  NAND4_X1  g716(.A1(new_n897), .A2(new_n382), .A3(new_n680), .A4(new_n899), .ZN(new_n918));
  OAI21_X1  g717(.A(G190gat), .B1(new_n890), .B2(new_n627), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1351gat));
  INV_X1    g720(.A(new_n874), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n663), .A2(new_n889), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n922), .A2(new_n875), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(G197gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n260), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n895), .A2(new_n730), .A3(new_n854), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n924), .A2(new_n926), .B1(new_n927), .B2(new_n925), .ZN(G1352gat));
  INV_X1    g727(.A(G204gat), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n895), .A2(new_n929), .A3(new_n642), .A4(new_n854), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n922), .A2(new_n643), .A3(new_n875), .A4(new_n923), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n931), .B(new_n932), .C1(new_n929), .C2(new_n933), .ZN(G1353gat));
  INV_X1    g733(.A(new_n923), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n874), .A2(new_n604), .A3(new_n876), .A4(new_n935), .ZN(new_n936));
  AND2_X1   g735(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n937));
  OAI21_X1  g736(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n936), .B2(new_n939), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n895), .A2(new_n854), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n604), .A2(new_n269), .ZN(new_n943));
  OAI22_X1  g742(.A1(new_n940), .A2(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1354gat));
  NOR4_X1   g743(.A1(new_n922), .A2(new_n627), .A3(new_n875), .A4(new_n923), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n680), .A2(new_n270), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n945), .A2(new_n270), .B1(new_n942), .B2(new_n946), .ZN(G1355gat));
endmodule


