

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XOR2_X1 U318 ( .A(n318), .B(n317), .Z(n286) );
  NOR2_X1 U319 ( .A1(n574), .A2(n386), .ZN(n387) );
  XNOR2_X1 U320 ( .A(n310), .B(KEYINPUT73), .ZN(n311) );
  XNOR2_X1 U321 ( .A(n322), .B(n311), .ZN(n312) );
  XNOR2_X1 U322 ( .A(n319), .B(n286), .ZN(n320) );
  XNOR2_X1 U323 ( .A(n321), .B(n320), .ZN(n571) );
  NOR2_X1 U324 ( .A1(n532), .A2(n446), .ZN(n562) );
  XNOR2_X1 U325 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U326 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  NAND2_X1 U327 ( .A1(G227GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U328 ( .A(G176GAT), .B(G99GAT), .Z(n288) );
  XNOR2_X1 U329 ( .A(G169GAT), .B(G15GAT), .ZN(n287) );
  XNOR2_X1 U330 ( .A(n288), .B(n287), .ZN(n290) );
  XOR2_X1 U331 ( .A(G43GAT), .B(G134GAT), .Z(n289) );
  XNOR2_X1 U332 ( .A(n290), .B(n289), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n305) );
  XOR2_X1 U334 ( .A(KEYINPUT20), .B(G71GAT), .Z(n294) );
  XNOR2_X1 U335 ( .A(G113GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n303) );
  XOR2_X1 U337 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n301) );
  XOR2_X1 U338 ( .A(KEYINPUT17), .B(G190GAT), .Z(n296) );
  XNOR2_X1 U339 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U341 ( .A(KEYINPUT19), .B(n297), .Z(n402) );
  XOR2_X1 U342 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n299) );
  XNOR2_X1 U343 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n428) );
  XNOR2_X1 U345 ( .A(n402), .B(n428), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(n303), .B(n302), .Z(n304) );
  XNOR2_X1 U348 ( .A(n305), .B(n304), .ZN(n532) );
  XNOR2_X1 U349 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n391) );
  XOR2_X1 U350 ( .A(KEYINPUT74), .B(G204GAT), .Z(n307) );
  XOR2_X1 U351 ( .A(G120GAT), .B(G57GAT), .Z(n419) );
  XOR2_X1 U352 ( .A(G106GAT), .B(G78GAT), .Z(n440) );
  XNOR2_X1 U353 ( .A(n419), .B(n440), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(n308), .B(KEYINPUT33), .Z(n314) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G85GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n309), .B(KEYINPUT75), .ZN(n322) );
  AND2_X1 U358 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(G148GAT), .B(n312), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n321) );
  XNOR2_X1 U361 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n315), .B(KEYINPUT13), .ZN(n345) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(G92GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n316), .B(G64GAT), .ZN(n392) );
  XNOR2_X1 U365 ( .A(n345), .B(n392), .ZN(n319) );
  XOR2_X1 U366 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n318) );
  XNOR2_X1 U367 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n317) );
  XOR2_X1 U368 ( .A(n322), .B(KEYINPUT9), .Z(n324) );
  XOR2_X1 U369 ( .A(G134GAT), .B(KEYINPUT80), .Z(n420) );
  XNOR2_X1 U370 ( .A(n420), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n324), .B(n323), .ZN(n337) );
  XOR2_X1 U372 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n326) );
  XNOR2_X1 U373 ( .A(KEYINPUT78), .B(KEYINPUT10), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U375 ( .A(G106GAT), .B(KEYINPUT81), .Z(n328) );
  XNOR2_X1 U376 ( .A(G162GAT), .B(KEYINPUT79), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U378 ( .A(n330), .B(n329), .Z(n335) );
  XOR2_X1 U379 ( .A(G190GAT), .B(G92GAT), .Z(n332) );
  NAND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U382 ( .A(G36GAT), .B(n333), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U384 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U385 ( .A(KEYINPUT8), .B(G50GAT), .Z(n339) );
  XNOR2_X1 U386 ( .A(G43GAT), .B(G29GAT), .ZN(n338) );
  XNOR2_X1 U387 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U388 ( .A(KEYINPUT7), .B(n340), .ZN(n374) );
  XNOR2_X1 U389 ( .A(n341), .B(n374), .ZN(n557) );
  XNOR2_X1 U390 ( .A(KEYINPUT36), .B(n557), .ZN(n578) );
  XOR2_X1 U391 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n343) );
  XNOR2_X1 U392 ( .A(KEYINPUT14), .B(KEYINPUT84), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n360) );
  XNOR2_X1 U394 ( .A(G15GAT), .B(KEYINPUT69), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n344), .B(G22GAT), .ZN(n369) );
  XNOR2_X1 U396 ( .A(n369), .B(n345), .ZN(n358) );
  XOR2_X1 U397 ( .A(G211GAT), .B(G64GAT), .Z(n347) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U400 ( .A(KEYINPUT12), .B(G78GAT), .Z(n349) );
  XNOR2_X1 U401 ( .A(G1GAT), .B(G57GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U403 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U404 ( .A(G155GAT), .B(KEYINPUT15), .Z(n353) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U407 ( .A(G127GAT), .B(n354), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U410 ( .A(n360), .B(n359), .ZN(n553) );
  NOR2_X1 U411 ( .A1(n578), .A2(n553), .ZN(n361) );
  XNOR2_X1 U412 ( .A(KEYINPUT45), .B(n361), .ZN(n376) );
  XOR2_X1 U413 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n363) );
  XNOR2_X1 U414 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n373) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(G141GAT), .ZN(n364) );
  XOR2_X1 U417 ( .A(n364), .B(G113GAT), .Z(n429) );
  XNOR2_X1 U418 ( .A(KEYINPUT68), .B(n429), .ZN(n366) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U421 ( .A(n367), .B(G197GAT), .Z(n371) );
  XNOR2_X1 U422 ( .A(G169GAT), .B(G36GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n368), .B(G8GAT), .ZN(n403) );
  XNOR2_X1 U424 ( .A(n403), .B(n369), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n375) );
  XNOR2_X1 U427 ( .A(n375), .B(n374), .ZN(n545) );
  XOR2_X1 U428 ( .A(KEYINPUT70), .B(n545), .Z(n559) );
  INV_X1 U429 ( .A(n559), .ZN(n453) );
  NAND2_X1 U430 ( .A1(n376), .A2(n453), .ZN(n377) );
  NOR2_X1 U431 ( .A1(n571), .A2(n377), .ZN(n378) );
  XOR2_X1 U432 ( .A(KEYINPUT116), .B(n378), .Z(n389) );
  INV_X1 U433 ( .A(n553), .ZN(n574) );
  INV_X1 U434 ( .A(n545), .ZN(n566) );
  XNOR2_X1 U435 ( .A(KEYINPUT41), .B(n571), .ZN(n547) );
  INV_X1 U436 ( .A(n547), .ZN(n379) );
  NAND2_X1 U437 ( .A1(n566), .A2(n379), .ZN(n380) );
  NAND2_X1 U438 ( .A1(n380), .A2(KEYINPUT46), .ZN(n384) );
  INV_X1 U439 ( .A(n380), .ZN(n382) );
  INV_X1 U440 ( .A(KEYINPUT46), .ZN(n381) );
  NAND2_X1 U441 ( .A1(n382), .A2(n381), .ZN(n383) );
  NAND2_X1 U442 ( .A1(n384), .A2(n383), .ZN(n385) );
  NAND2_X1 U443 ( .A1(n385), .A2(n557), .ZN(n386) );
  XNOR2_X1 U444 ( .A(KEYINPUT47), .B(n387), .ZN(n388) );
  NAND2_X1 U445 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n527) );
  XOR2_X1 U447 ( .A(KEYINPUT98), .B(n392), .Z(n394) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n401) );
  XOR2_X1 U450 ( .A(KEYINPUT21), .B(G204GAT), .Z(n396) );
  XNOR2_X1 U451 ( .A(G197GAT), .B(G211GAT), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U453 ( .A(KEYINPUT91), .B(KEYINPUT89), .Z(n398) );
  XNOR2_X1 U454 ( .A(G218GAT), .B(KEYINPUT90), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U456 ( .A(n400), .B(n399), .Z(n439) );
  XOR2_X1 U457 ( .A(n401), .B(n439), .Z(n405) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(n405), .B(n404), .Z(n518) );
  XNOR2_X1 U460 ( .A(KEYINPUT123), .B(n518), .ZN(n406) );
  NOR2_X1 U461 ( .A1(n527), .A2(n406), .ZN(n407) );
  XNOR2_X1 U462 ( .A(KEYINPUT54), .B(n407), .ZN(n431) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n409) );
  XNOR2_X1 U464 ( .A(KEYINPUT92), .B(KEYINPUT94), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U466 ( .A(KEYINPUT6), .B(n410), .Z(n412) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U469 ( .A(n413), .B(KEYINPUT4), .Z(n418) );
  XOR2_X1 U470 ( .A(G148GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U473 ( .A(G155GAT), .B(n416), .ZN(n443) );
  XOR2_X1 U474 ( .A(n443), .B(KEYINPUT93), .Z(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n424) );
  XOR2_X1 U476 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n422) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U479 ( .A(n424), .B(n423), .Z(n426) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G85GAT), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n467) );
  XNOR2_X1 U484 ( .A(KEYINPUT97), .B(n467), .ZN(n457) );
  NAND2_X1 U485 ( .A1(n431), .A2(n457), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n432), .B(KEYINPUT64), .ZN(n565) );
  XOR2_X1 U487 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n434) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U490 ( .A(KEYINPUT23), .B(G141GAT), .Z(n436) );
  XNOR2_X1 U491 ( .A(G50GAT), .B(G22GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U493 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n461) );
  NOR2_X1 U497 ( .A1(n565), .A2(n461), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n562), .A2(n379), .ZN(n449) );
  XOR2_X1 U500 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n447) );
  XNOR2_X1 U501 ( .A(n447), .B(G176GAT), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  INV_X1 U503 ( .A(n557), .ZN(n539) );
  NAND2_X1 U504 ( .A1(n562), .A2(n539), .ZN(n452) );
  XOR2_X1 U505 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n450) );
  INV_X1 U506 ( .A(n457), .ZN(n515) );
  NOR2_X1 U507 ( .A1(n571), .A2(n453), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(KEYINPUT77), .ZN(n485) );
  NOR2_X1 U509 ( .A1(n539), .A2(n553), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n455), .B(KEYINPUT16), .ZN(n472) );
  XOR2_X1 U511 ( .A(n518), .B(KEYINPUT99), .Z(n456) );
  XOR2_X1 U512 ( .A(n456), .B(KEYINPUT27), .Z(n464) );
  OR2_X1 U513 ( .A1(n464), .A2(n457), .ZN(n528) );
  XOR2_X1 U514 ( .A(n461), .B(KEYINPUT28), .Z(n530) );
  NAND2_X1 U515 ( .A1(n532), .A2(n530), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n528), .A2(n458), .ZN(n470) );
  INV_X1 U517 ( .A(n532), .ZN(n521) );
  AND2_X1 U518 ( .A1(n521), .A2(n518), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n461), .A2(n459), .ZN(n460) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n460), .Z(n466) );
  NAND2_X1 U521 ( .A1(n461), .A2(n532), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT100), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT26), .B(n463), .ZN(n564) );
  NOR2_X1 U524 ( .A1(n564), .A2(n464), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n482) );
  INV_X1 U528 ( .A(n482), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n502) );
  NOR2_X1 U530 ( .A1(n485), .A2(n502), .ZN(n479) );
  NAND2_X1 U531 ( .A1(n515), .A2(n479), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n518), .A2(n479), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U537 ( .A1(n479), .A2(n521), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  INV_X1 U540 ( .A(n530), .ZN(n524) );
  NAND2_X1 U541 ( .A1(n524), .A2(n479), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(KEYINPUT102), .ZN(n481) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XNOR2_X1 U544 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n491) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT105), .Z(n489) );
  NOR2_X1 U546 ( .A1(n578), .A2(n482), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n483), .A2(n553), .ZN(n484) );
  XOR2_X1 U548 ( .A(KEYINPUT37), .B(n484), .Z(n513) );
  NOR2_X1 U549 ( .A1(n513), .A2(n485), .ZN(n487) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n497) );
  NAND2_X1 U552 ( .A1(n497), .A2(n515), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n518), .A2(n497), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(KEYINPUT106), .ZN(n493) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n495) );
  NAND2_X1 U559 ( .A1(n497), .A2(n521), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n499) );
  NAND2_X1 U563 ( .A1(n497), .A2(n524), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  NAND2_X1 U567 ( .A1(n545), .A2(n379), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(KEYINPUT110), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n514), .A2(n502), .ZN(n508) );
  NAND2_X1 U570 ( .A1(n508), .A2(n515), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  XOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT111), .Z(n506) );
  NAND2_X1 U573 ( .A1(n508), .A2(n518), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n521), .A2(n508), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U578 ( .A1(n508), .A2(n524), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n510), .B(n509), .ZN(n512) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT113), .Z(n511) );
  XNOR2_X1 U581 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n523), .A2(n515), .ZN(n516) );
  XNOR2_X1 U584 ( .A(KEYINPUT114), .B(n516), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT115), .Z(n520) );
  NAND2_X1 U587 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n521), .A2(n523), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(KEYINPUT118), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n530), .A2(n543), .ZN(n531) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n540), .A2(n559), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U601 ( .A1(n540), .A2(n379), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n537) );
  NAND2_X1 U604 ( .A1(n540), .A2(n574), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  INV_X1 U610 ( .A(n564), .ZN(n544) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n545), .A2(n556), .ZN(n546) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n556), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(KEYINPUT120), .B(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n556), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT122), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n574), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(KEYINPUT126), .B(KEYINPUT59), .ZN(n570) );
  XOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT60), .Z(n568) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n576), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n576), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U641 ( .A(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

