//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G221), .A2(G218), .A3(G220), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n456), .A2(KEYINPUT67), .A3(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n452), .ZN(new_n459));
  AOI21_X1  g034(.A(KEYINPUT67), .B1(new_n456), .B2(G2106), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n466), .A2(new_n469), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n464), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT68), .B(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n476), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n470), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g059(.A1(G124), .A2(new_n482), .B1(new_n484), .B2(G136), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n470), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n492), .A2(new_n496), .B1(new_n480), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G138), .C1(new_n462), .C2(new_n463), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n502), .B2(new_n476), .ZN(new_n503));
  INV_X1    g078(.A(new_n500), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n469), .A2(new_n480), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n498), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n515), .A2(G62), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n515), .A2(G88), .A3(new_n517), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G50), .A3(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n516), .B1(new_n511), .B2(new_n514), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G62), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n531), .B2(new_n519), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT72), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n528), .A2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT73), .ZN(new_n536));
  XOR2_X1   g111(.A(new_n536), .B(KEYINPUT7), .Z(new_n537));
  NAND2_X1  g112(.A1(new_n522), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G51), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n530), .A2(new_n522), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n537), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n529), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  INV_X1    g123(.A(G52), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n543), .A2(new_n548), .B1(new_n549), .B2(new_n538), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n547), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n543), .A2(new_n553), .B1(new_n554), .B2(new_n538), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT74), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n529), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g137(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n563));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT76), .B1(new_n538), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n522), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  OAI211_X1 g147(.A(KEYINPUT76), .B(new_n572), .C1(new_n538), .C2(new_n567), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n575), .A2(new_n529), .B1(new_n576), .B2(new_n543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  AND3_X1   g156(.A1(new_n530), .A2(G87), .A3(new_n522), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n530), .A2(G74), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G49), .B2(new_n539), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n530), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G48), .B2(new_n539), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n530), .A2(G86), .A3(new_n522), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(G305));
  INV_X1    g170(.A(new_n543), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G85), .B1(G47), .B2(new_n539), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n598), .A2(KEYINPUT79), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n598), .B2(KEYINPUT79), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(KEYINPUT80), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n543), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n543), .B2(new_n606), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n538), .B2(KEYINPUT82), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT82), .B2(new_n538), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n530), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n529), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n605), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n605), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n578), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n578), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g202(.A1(G123), .A2(new_n482), .B1(new_n484), .B2(G135), .ZN(new_n628));
  OAI221_X1 g203(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n480), .A2(new_n471), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT84), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT85), .Z(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  INV_X1    g238(.A(new_n660), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n664), .B2(new_n658), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n658), .B(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n667), .B2(new_n664), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n664), .A3(new_n661), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2100), .Z(new_n671));
  XOR2_X1   g246(.A(KEYINPUT87), .B(G2096), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  INV_X1    g256(.A(new_n676), .ZN(new_n682));
  INV_X1    g257(.A(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n681), .B(new_n685), .C1(new_n682), .C2(new_n684), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G6), .ZN(new_n696));
  INV_X1    g271(.A(G305), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT90), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G23), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT91), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G288), .B2(new_n695), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT33), .B(G1976), .Z(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G22), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G166), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1971), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n701), .A2(new_n702), .A3(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G24), .B(G290), .S(G16), .Z(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G1986), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(G1986), .ZN(new_n715));
  AOI22_X1  g290(.A1(G119), .A2(new_n482), .B1(new_n484), .B2(G131), .ZN(new_n716));
  OAI221_X1 g291(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n718), .S(G29), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  XOR2_X1   g295(.A(new_n719), .B(new_n720), .Z(new_n721));
  NOR3_X1   g296(.A1(new_n714), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n712), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n702), .B1(new_n701), .B2(new_n711), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT36), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n726), .A2(new_n727), .A3(new_n712), .A4(new_n722), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G35), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n730), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT102), .B(G2090), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n730), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n730), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT100), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2078), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G171), .A2(new_n695), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G5), .B2(new_n695), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n745), .B2(G34), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G34), .B2(new_n745), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n730), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n743), .A2(new_n744), .B1(G2084), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n695), .A2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G168), .B2(new_n695), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT98), .B(G1966), .Z(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n560), .A2(new_n695), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n695), .B2(G19), .ZN(new_n756));
  INV_X1    g331(.A(G1341), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n750), .B1(new_n752), .B2(new_n754), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT26), .Z(new_n760));
  INV_X1    g335(.A(G129), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n481), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n471), .A2(G105), .ZN(new_n763));
  INV_X1    g338(.A(G141), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n483), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(new_n730), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n730), .B2(G32), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n632), .B2(new_n730), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n730), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n482), .A2(G128), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n484), .A2(G140), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT93), .B1(G104), .B2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(KEYINPUT93), .A2(G104), .A3(G2105), .ZN(new_n779));
  OAI221_X1 g354(.A(G2104), .B1(new_n778), .B2(new_n779), .C1(new_n469), .C2(G116), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n775), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n774), .B1(new_n781), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G28), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT30), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n787));
  OR2_X1    g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  NAND2_X1  g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n768), .B2(new_n769), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n771), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n752), .A2(new_n754), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(new_n744), .C2(new_n743), .ZN(new_n794));
  NOR2_X1   g369(.A1(G4), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n616), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT92), .B(G1348), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n741), .A2(new_n758), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n749), .A2(G2084), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n484), .A2(G139), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n804), .B(new_n805), .C1(new_n469), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  MUX2_X1   g383(.A(G33), .B(new_n808), .S(G29), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G2072), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n801), .B(new_n810), .C1(new_n757), .C2(new_n756), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n695), .A2(G20), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT23), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n578), .B2(new_n695), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT104), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT103), .ZN(new_n816));
  INV_X1    g391(.A(G1956), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n799), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n729), .A2(new_n819), .ZN(G150));
  NOR2_X1   g395(.A1(G150), .A2(KEYINPUT105), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT105), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n729), .B2(new_n819), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n616), .A2(G559), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT38), .Z(new_n826));
  AOI22_X1  g401(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n529), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n543), .A2(new_n829), .B1(new_n830), .B2(new_n538), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n559), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n556), .A2(new_n558), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n826), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n832), .A2(new_n839), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n632), .B(new_n478), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n487), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT106), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n503), .A2(new_n847), .A3(new_n507), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n503), .B2(new_n507), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n498), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n781), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n808), .B(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n766), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n766), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n718), .B(KEYINPUT108), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n636), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n482), .A2(G130), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT107), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n484), .A2(G142), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n469), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n857), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n855), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n853), .A2(new_n864), .A3(new_n854), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT109), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n855), .A2(new_n864), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n846), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n846), .B(KEYINPUT110), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n866), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n876), .B2(new_n871), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT40), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n846), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n865), .A2(new_n868), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n870), .A2(new_n871), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n883), .A2(new_n884), .A3(new_n877), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n879), .A2(new_n885), .ZN(G395));
  INV_X1    g461(.A(KEYINPUT113), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT112), .ZN(new_n888));
  NAND2_X1  g463(.A1(G290), .A2(new_n697), .ZN(new_n889));
  INV_X1    g464(.A(G288), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n528), .A2(new_n533), .A3(KEYINPUT111), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT111), .B1(new_n528), .B2(new_n533), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n602), .A2(G305), .A3(new_n603), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n889), .A2(new_n893), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n894), .A2(new_n889), .B1(new_n893), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n888), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n893), .A2(new_n895), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT112), .A3(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n836), .B(new_n624), .Z(new_n906));
  XNOR2_X1  g481(.A(G299), .B(new_n616), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n907), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n908), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT42), .B1(new_n902), .B2(new_n896), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n905), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(new_n899), .B2(new_n903), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n911), .A2(new_n906), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n917), .A2(new_n913), .B1(new_n908), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(G868), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n832), .A2(G868), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n887), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AOI211_X1 g499(.A(KEYINPUT113), .B(new_n922), .C1(new_n920), .C2(G868), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(G295));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n923), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT114), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(KEYINPUT114), .A2(KEYINPUT44), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n899), .A2(new_n903), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n834), .A2(G301), .A3(new_n835), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G301), .B1(new_n834), .B2(new_n835), .ZN(new_n935));
  OAI21_X1  g510(.A(G286), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(G168), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n907), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n910), .A2(new_n938), .A3(new_n936), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n932), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n904), .A2(new_n940), .A3(new_n941), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n930), .B(new_n931), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n928), .A3(new_n929), .A4(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n948), .A2(new_n952), .ZN(G397));
  XOR2_X1   g528(.A(KEYINPUT115), .B(G1384), .Z(new_n954));
  AOI21_X1  g529(.A(KEYINPUT45), .B1(new_n850), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n472), .A2(G40), .A3(new_n477), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n781), .B(new_n783), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n766), .B(G1996), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT116), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n718), .B(new_n720), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g539(.A1(G290), .A2(G1986), .ZN(new_n965));
  NAND2_X1  g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n528), .A2(new_n533), .A3(G8), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n972));
  INV_X1    g547(.A(new_n498), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n503), .A2(new_n507), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT106), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n503), .A2(new_n847), .A3(new_n507), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n508), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n957), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n972), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1971), .ZN(new_n986));
  INV_X1    g561(.A(new_n978), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n850), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n956), .B1(new_n981), .B2(new_n982), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(KEYINPUT117), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n985), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT50), .B1(new_n977), .B2(G1384), .ZN(new_n992));
  INV_X1    g567(.A(G2090), .ZN(new_n993));
  INV_X1    g568(.A(new_n981), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n956), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n971), .B1(new_n998), .B2(G8), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n850), .A2(new_n995), .A3(new_n980), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n956), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n993), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n1000), .B(new_n970), .C1(new_n991), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n850), .A2(new_n980), .A3(new_n957), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n591), .A2(new_n1008), .A3(new_n593), .A4(new_n594), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n539), .A2(G48), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n530), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n529), .ZN(new_n1012));
  INV_X1    g587(.A(new_n592), .ZN(new_n1013));
  OAI21_X1  g588(.A(G1981), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1009), .A2(KEYINPUT49), .A3(new_n1014), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1009), .A2(KEYINPUT118), .A3(new_n1014), .A4(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n890), .B2(G1976), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1006), .B(G8), .C1(G288), .C2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(KEYINPUT52), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n999), .A2(new_n1005), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n982), .B1(new_n977), .B2(G1384), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n957), .B1(new_n981), .B2(new_n982), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n754), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2084), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1001), .A2(new_n1036), .A3(new_n1002), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n537), .B2(new_n544), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1042), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1001), .A2(new_n1036), .A3(new_n1002), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n850), .A2(new_n980), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1033), .B1(new_n1048), .B2(new_n982), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1049), .B2(new_n754), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1042), .B1(new_n1050), .B2(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1044), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G2078), .ZN(new_n1055));
  INV_X1    g630(.A(new_n990), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT117), .B1(new_n988), .B2(new_n989), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1055), .A2(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1049), .A2(new_n1062), .B1(new_n1063), .B2(new_n744), .ZN(new_n1064));
  AOI21_X1  g639(.A(G301), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1044), .B(KEYINPUT62), .C1(new_n1046), .C2(new_n1051), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1031), .A2(new_n1054), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1023), .A2(new_n1026), .A3(new_n890), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1007), .B1(new_n1068), .B2(new_n1009), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1030), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1005), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n577), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n573), .A4(new_n571), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT57), .B1(new_n574), .B2(new_n577), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1956), .B1(new_n992), .B2(new_n996), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n988), .A2(new_n989), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n995), .B1(new_n850), .B2(new_n980), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n957), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n817), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1076), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n988), .A2(new_n989), .A3(new_n1078), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1348), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1006), .A2(G2067), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n616), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1080), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1996), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n988), .A2(new_n1092), .A3(new_n989), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1006), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT58), .B(G1341), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n560), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT59), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n560), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT119), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT121), .A4(new_n1085), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1080), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1086), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1102), .A2(new_n1103), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1088), .A2(new_n1089), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n616), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1109), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n616), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1114), .B2(new_n1110), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1091), .B1(new_n1108), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1052), .ZN(new_n1120));
  INV_X1    g695(.A(new_n999), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1005), .A2(new_n1030), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G301), .B(KEYINPUT54), .ZN(new_n1123));
  AOI21_X1  g698(.A(G2078), .B1(new_n985), .B2(new_n990), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1064), .B(new_n1123), .C1(new_n1124), .C2(new_n1059), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n988), .A2(new_n957), .A3(new_n1062), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1003), .A2(G1961), .B1(new_n955), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(new_n1123), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1067), .B(new_n1071), .C1(new_n1119), .C2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1050), .A2(G8), .A3(G168), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1031), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n991), .A2(new_n1004), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n971), .B1(new_n1136), .B2(G8), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1137), .A2(new_n1135), .A3(new_n1132), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1134), .A2(new_n1135), .B1(new_n1122), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n968), .B1(new_n1131), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n958), .B1(new_n766), .B2(new_n959), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n955), .A2(new_n957), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(KEYINPUT46), .A3(new_n1092), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1143), .A2(KEYINPUT126), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(KEYINPUT126), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT46), .B1(new_n1142), .B2(new_n1092), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT125), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(KEYINPUT47), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(KEYINPUT47), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n965), .A2(new_n958), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT48), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1150), .A2(new_n1151), .B1(new_n964), .B2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n716), .A2(new_n717), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n962), .A2(new_n720), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n781), .A2(G2067), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n958), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1154), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1140), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT127), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1140), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g742(.A(G319), .B1(new_n655), .B2(new_n654), .ZN(new_n1169));
  NOR3_X1   g743(.A1(G229), .A2(G227), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n1170), .B1(new_n883), .B2(new_n877), .ZN(new_n1171));
  NOR2_X1   g745(.A1(new_n946), .A2(new_n947), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1171), .A2(new_n1172), .ZN(G308));
  OR2_X1    g747(.A1(new_n1171), .A2(new_n1172), .ZN(G225));
endmodule


