//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND3_X1  g0012(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n212), .B1(new_n214), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G226), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G13), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n243), .A2(G1), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G1), .B2(new_n207), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G20), .A2(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT15), .B(G87), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n207), .A2(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT8), .B(G58), .Z(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n248), .B1(new_n247), .B2(new_n253), .C1(new_n260), .C2(new_n252), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G238), .ZN(new_n266));
  INV_X1    g0066(.A(G107), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n262), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n266), .B1(new_n267), .B2(new_n268), .C1(new_n229), .C2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n250), .B1(G33), .B2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n275), .B1(new_n279), .B2(G244), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n272), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n272), .B(new_n285), .C1(new_n281), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n290), .A3(new_n286), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n261), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(G179), .B1(new_n284), .B2(new_n286), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT69), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n284), .A2(new_n296), .A3(new_n286), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n261), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n293), .A2(new_n294), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n292), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT72), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n265), .A2(new_n302), .A3(G232), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n268), .A2(G226), .A3(new_n262), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n265), .B2(G232), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n271), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT13), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n275), .B1(new_n279), .B2(G238), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n308), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n288), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(new_n310), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n290), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n258), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n256), .A2(new_n247), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n251), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT74), .ZN(new_n325));
  XOR2_X1   g0125(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n326));
  XNOR2_X1  g0126(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n253), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G68), .ZN(new_n329));
  INV_X1    g0129(.A(G68), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n244), .A2(G20), .A3(new_n330), .ZN(new_n331));
  OR3_X1    g0131(.A1(new_n331), .A2(KEYINPUT75), .A3(KEYINPUT12), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT75), .B1(new_n331), .B2(KEYINPUT12), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(KEYINPUT12), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n327), .A2(new_n329), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n320), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n313), .A2(new_n339), .A3(G179), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT76), .B1(new_n318), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(G169), .B1(new_n311), .B2(new_n312), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(KEYINPUT14), .B(G169), .C1(new_n311), .C2(new_n312), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n340), .A2(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n301), .B(new_n338), .C1(new_n337), .C2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(KEYINPUT8), .A2(G58), .ZN(new_n349));
  INV_X1    g0149(.A(G58), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT65), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT65), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G58), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n349), .B1(new_n354), .B2(KEYINPUT8), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n246), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n355), .B2(new_n253), .ZN(new_n357));
  INV_X1    g0157(.A(G159), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n321), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n201), .B1(new_n354), .B2(G68), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n207), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n263), .A2(new_n207), .A3(new_n264), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n264), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n330), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n362), .A2(new_n367), .A3(KEYINPUT16), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  AND2_X1   g0169(.A1(KEYINPUT3), .A2(G33), .ZN(new_n370));
  NOR2_X1   g0170(.A1(KEYINPUT3), .A2(G33), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n372), .B2(new_n207), .ZN(new_n373));
  INV_X1    g0173(.A(new_n366), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT65), .B(G58), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n215), .B1(new_n376), .B2(new_n330), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n359), .B1(new_n377), .B2(G20), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n369), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n251), .B1(new_n368), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n357), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n275), .B1(new_n279), .B2(G232), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  INV_X1    g0184(.A(G33), .ZN(new_n385));
  INV_X1    g0185(.A(G87), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n265), .B2(G226), .ZN(new_n388));
  OAI211_X1 g0188(.A(G223), .B(new_n262), .C1(new_n370), .C2(new_n371), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(G226), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n391));
  INV_X1    g0191(.A(new_n387), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n389), .A2(new_n391), .A3(new_n384), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n271), .ZN(new_n394));
  OAI211_X1 g0194(.A(G190), .B(new_n383), .C1(new_n390), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT78), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(new_n393), .A3(new_n271), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n290), .B1(new_n399), .B2(new_n383), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT79), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT16), .B1(new_n362), .B2(new_n367), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n375), .A2(new_n378), .A3(new_n369), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n252), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT77), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT79), .ZN(new_n406));
  INV_X1    g0206(.A(new_n383), .ZN(new_n407));
  INV_X1    g0207(.A(new_n394), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n398), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(new_n395), .C1(new_n409), .C2(new_n290), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n382), .A2(new_n401), .A3(new_n405), .A4(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n357), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n404), .B2(KEYINPUT77), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n381), .B(new_n252), .C1(new_n402), .C2(new_n403), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n417), .A2(KEYINPUT17), .A3(new_n410), .A4(new_n401), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(G169), .B1(new_n399), .B2(new_n383), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n341), .B2(new_n409), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n415), .B2(new_n416), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT18), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n421), .C1(new_n415), .C2(new_n416), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT71), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n275), .B1(new_n279), .B2(G226), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n265), .A2(G223), .ZN(new_n431));
  INV_X1    g0231(.A(G222), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n431), .B1(new_n247), .B2(new_n268), .C1(new_n432), .C2(new_n269), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(new_n271), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT70), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(G200), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT70), .B1(new_n434), .B2(new_n290), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n355), .A2(new_n207), .A3(G33), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n252), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n246), .A2(G50), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n253), .B2(G50), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT9), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT9), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n442), .B2(new_n444), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n448), .C1(new_n288), .C2(new_n435), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n439), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT10), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n428), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n439), .A2(new_n449), .A3(KEYINPUT71), .A4(KEYINPUT10), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(new_n451), .B2(new_n450), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n445), .B1(new_n435), .B2(new_n296), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n434), .A2(new_n341), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n348), .A2(new_n427), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n206), .B(G45), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(G1), .B(G13), .C1(new_n385), .C2(new_n276), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G270), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n466), .A2(new_n274), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(G257), .B(new_n262), .C1(new_n370), .C2(new_n371), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n263), .A2(G303), .A3(new_n264), .ZN(new_n473));
  OAI211_X1 g0273(.A(G264), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(KEYINPUT81), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n265), .B2(G264), .ZN(new_n477));
  OAI211_X1 g0277(.A(KEYINPUT82), .B(new_n271), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n268), .A2(new_n476), .A3(G264), .A4(G1698), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n472), .A4(new_n473), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT82), .B1(new_n482), .B2(new_n271), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n471), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT83), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n471), .B(new_n486), .C1(new_n479), .C2(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n385), .A2(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  AOI21_X1  g0289(.A(G20), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G116), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n207), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n251), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g0293(.A(new_n493), .B(KEYINPUT20), .Z(new_n494));
  NAND2_X1  g0294(.A1(new_n245), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n206), .A2(G33), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n252), .A2(new_n245), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(new_n491), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n296), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n485), .A2(new_n487), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n485), .A2(KEYINPUT21), .A3(new_n487), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n494), .A2(new_n499), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n471), .B(G179), .C1(new_n479), .C2(new_n483), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n485), .A2(new_n290), .A3(new_n487), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G190), .B1(new_n485), .B2(new_n487), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n267), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  XOR2_X1   g0315(.A(G97), .B(G107), .Z(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(G20), .B1(G77), .B2(new_n258), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n373), .B2(new_n374), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n252), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n246), .A2(G97), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n497), .B2(G97), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G244), .B1(new_n370), .B2(new_n371), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(G1698), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n268), .A2(G244), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n528), .A3(new_n489), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n268), .A2(G250), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n262), .B1(new_n530), .B2(KEYINPUT4), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n271), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n466), .A2(G257), .A3(new_n467), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n470), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n532), .A2(new_n534), .A3(new_n288), .ZN(new_n535));
  AOI21_X1  g0335(.A(G200), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n523), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n532), .A2(new_n534), .A3(G179), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n296), .B1(new_n532), .B2(new_n534), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(new_n520), .B2(new_n522), .ZN(new_n540));
  INV_X1    g0340(.A(G250), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n206), .B2(G45), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n467), .A2(new_n542), .B1(KEYINPUT80), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n467), .A2(new_n542), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(KEYINPUT80), .ZN(new_n546));
  OAI211_X1 g0346(.A(G238), .B(new_n262), .C1(new_n370), .C2(new_n371), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(new_n524), .C2(new_n262), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n271), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n296), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n268), .A2(new_n207), .A3(G68), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n207), .B1(new_n304), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n386), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(G107), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n554), .B1(new_n304), .B2(G20), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n553), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n251), .B1(new_n246), .B2(new_n255), .ZN(new_n561));
  INV_X1    g0361(.A(new_n255), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n498), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n552), .B(new_n564), .C1(G179), .C2(new_n551), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n551), .A2(G200), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n498), .A2(G87), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n546), .A2(new_n550), .A3(G190), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n561), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n537), .A2(new_n540), .A3(new_n565), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n468), .A2(G264), .ZN(new_n571));
  OAI211_X1 g0371(.A(G250), .B(new_n262), .C1(new_n370), .C2(new_n371), .ZN(new_n572));
  OAI211_X1 g0372(.A(G257), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G294), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n575), .A2(KEYINPUT85), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT85), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n572), .A2(new_n573), .A3(new_n577), .A4(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n271), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n470), .B(new_n571), .C1(new_n576), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G169), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n575), .A2(KEYINPUT85), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n271), .A3(new_n578), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n583), .A2(G179), .A3(new_n470), .A4(new_n571), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n244), .A2(G20), .A3(new_n267), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n586), .B(KEYINPUT25), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(G107), .B2(new_n498), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n268), .A2(new_n207), .A3(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n268), .A2(new_n591), .A3(new_n207), .A4(G87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n267), .A2(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT84), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT23), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(KEYINPUT23), .C2(new_n594), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n594), .B2(KEYINPUT23), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n600), .A3(KEYINPUT24), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n251), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT24), .B1(new_n593), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n588), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n585), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n580), .A2(G190), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n580), .A2(new_n290), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n570), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n510), .A2(new_n514), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n462), .A2(new_n611), .ZN(G372));
  INV_X1    g0412(.A(new_n459), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n347), .A2(new_n337), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n297), .B(new_n261), .C1(new_n293), .C2(new_n294), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n293), .A2(new_n294), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n419), .A2(new_n338), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n426), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n613), .B1(new_n620), .B2(new_n454), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  INV_X1    g0422(.A(new_n551), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n623), .A2(new_n341), .B1(new_n561), .B2(new_n563), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n549), .A2(new_n626), .A3(new_n271), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n546), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n296), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(G200), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n568), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n561), .A2(KEYINPUT87), .A3(new_n567), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT87), .B1(new_n561), .B2(new_n567), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n630), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n622), .B1(new_n636), .B2(new_n540), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n565), .A2(new_n569), .ZN(new_n638));
  XOR2_X1   g0438(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n639));
  OR3_X1    g0439(.A1(new_n638), .A2(new_n540), .A3(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n637), .A2(new_n640), .B1(new_n624), .B2(new_n629), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n585), .A2(new_n604), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT88), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n585), .A2(new_n604), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT89), .B1(new_n510), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n508), .B1(new_n501), .B2(new_n502), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n646), .A2(new_n648), .A3(KEYINPUT89), .A4(new_n504), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n537), .A2(new_n540), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n636), .A2(new_n609), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n641), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n621), .B1(new_n462), .B2(new_n654), .ZN(G369));
  INV_X1    g0455(.A(new_n244), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .A3(G20), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT27), .B1(new_n656), .B2(G20), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n506), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n510), .B2(new_n514), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n510), .B2(new_n663), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n602), .A2(new_n603), .ZN(new_n668));
  INV_X1    g0468(.A(new_n608), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n668), .B(new_n588), .C1(new_n669), .C2(new_n606), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n604), .A2(new_n661), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n642), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n605), .A2(new_n661), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n662), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(new_n672), .ZN(new_n678));
  INV_X1    g0478(.A(new_n645), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n644), .B1(new_n585), .B2(new_n604), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n662), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(G399));
  NAND2_X1  g0484(.A1(new_n210), .A2(new_n276), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n557), .A2(G107), .A3(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n216), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n485), .A2(new_n487), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n288), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n505), .B1(new_n692), .B2(new_n511), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n537), .A2(new_n540), .ZN(new_n694));
  INV_X1    g0494(.A(new_n638), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n642), .A4(new_n670), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n676), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  AOI21_X1  g0498(.A(G179), .B1(new_n532), .B2(new_n534), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n699), .A2(new_n628), .A3(new_n580), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n485), .A3(new_n487), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n470), .A2(new_n533), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n524), .A2(new_n525), .B1(G33), .B2(G283), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n525), .B1(new_n268), .B2(G250), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n704), .B(new_n528), .C1(new_n262), .C2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n703), .B1(new_n706), .B2(new_n271), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n623), .A3(new_n571), .A4(new_n583), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n702), .B1(new_n708), .B2(new_n507), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n532), .A2(new_n534), .A3(new_n546), .A4(new_n550), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n583), .A2(new_n571), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n469), .A2(new_n470), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n482), .A2(new_n271), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT82), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n716), .B2(new_n478), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n712), .A2(KEYINPUT30), .A3(G179), .A4(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n701), .A2(new_n709), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT92), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT92), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n701), .A2(new_n721), .A3(new_n718), .A4(new_n709), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT31), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n697), .A2(new_n698), .B1(new_n723), .B2(new_n662), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n662), .A2(new_n698), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT91), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n690), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n651), .B1(new_n676), .B2(new_n605), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n630), .B(KEYINPUT93), .ZN(new_n731));
  INV_X1    g0531(.A(new_n635), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n568), .A3(new_n631), .ZN(new_n733));
  INV_X1    g0533(.A(new_n540), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(KEYINPUT26), .A3(new_n734), .A4(new_n630), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n639), .B1(new_n638), .B2(new_n540), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n731), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n661), .B1(new_n730), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT89), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n676), .B2(new_n681), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n649), .A3(new_n651), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n661), .B1(new_n742), .B2(new_n641), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n739), .B1(new_n743), .B2(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n729), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n689), .B1(new_n746), .B2(G1), .ZN(G364));
  NOR2_X1   g0547(.A1(new_n243), .A2(G20), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G45), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n685), .A2(G1), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n665), .A2(G330), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n667), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n665), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n250), .B1(G20), .B2(new_n296), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n341), .A2(new_n290), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT96), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n207), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n358), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT98), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n761), .A2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n207), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G97), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n207), .A2(new_n288), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n775), .A2(new_n290), .A3(G179), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n268), .B1(new_n777), .B2(new_n386), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT99), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n341), .A2(new_n290), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n762), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n330), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n341), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n762), .A2(new_n783), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n376), .B1(new_n785), .B2(new_n247), .ZN(new_n786));
  INV_X1    g0586(.A(new_n762), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(G179), .A3(new_n290), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n782), .B(new_n786), .C1(G107), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT95), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n774), .A2(new_n780), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(new_n774), .B2(new_n780), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n778), .A2(KEYINPUT99), .B1(G50), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n773), .A2(new_n779), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n769), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n781), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n777), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n788), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n803), .A2(new_n804), .B1(new_n785), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n784), .A2(new_n807), .ZN(new_n808));
  NOR4_X1   g0608(.A1(new_n802), .A2(new_n806), .A3(new_n268), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  INV_X1    g0610(.A(G326), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n771), .C1(new_n811), .C2(new_n793), .ZN(new_n812));
  INV_X1    g0612(.A(new_n766), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G329), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n759), .B1(new_n797), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n756), .A2(new_n759), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n210), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n372), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G355), .B1(new_n491), .B2(new_n818), .ZN(new_n820));
  INV_X1    g0620(.A(new_n216), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G45), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n238), .B2(G45), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n818), .A2(new_n268), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n820), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n817), .B1(new_n826), .B2(KEYINPUT94), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(KEYINPUT94), .B2(new_n826), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n815), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n753), .B1(new_n758), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n752), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NOR3_X1   g0632(.A1(new_n615), .A2(new_n616), .A3(new_n661), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n261), .A2(new_n661), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n292), .A2(new_n836), .B1(new_n615), .B2(new_n616), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n654), .B2(new_n661), .ZN(new_n839));
  INV_X1    g0639(.A(new_n837), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n833), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n653), .A2(new_n662), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n728), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n839), .A2(new_n728), .A3(new_n842), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n750), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(KEYINPUT100), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(KEYINPUT100), .B2(new_n845), .ZN(new_n847));
  INV_X1    g0647(.A(new_n785), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G150), .A2(new_n798), .B1(new_n848), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G143), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n784), .C1(new_n793), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n803), .A2(new_n330), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n268), .B1(new_n777), .B2(new_n202), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(new_n772), .C2(new_n354), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n813), .A2(G132), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n854), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n766), .A2(new_n805), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n777), .A2(new_n267), .B1(new_n785), .B2(new_n491), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n803), .A2(new_n386), .B1(new_n804), .B2(new_n781), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n372), .B1(new_n784), .B2(new_n810), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n773), .C1(new_n801), .C2(new_n793), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n860), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n759), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n759), .A2(new_n754), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n750), .B1(new_n247), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n868), .B(new_n870), .C1(new_n841), .C2(new_n755), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n847), .A2(new_n871), .ZN(G384));
  INV_X1    g0672(.A(new_n214), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n873), .B(G116), .C1(KEYINPUT35), .C2(new_n517), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(KEYINPUT35), .B2(new_n517), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT36), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n821), .B(G77), .C1(new_n330), .C2(new_n376), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n202), .A2(G68), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n206), .B(G13), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n833), .B1(new_n743), .B2(new_n841), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n380), .A2(new_n414), .ZN(new_n883));
  INV_X1    g0683(.A(new_n659), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n419), .B2(new_n426), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n659), .B(KEYINPUT102), .Z(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n415), .B2(new_n416), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n411), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT101), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n422), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT101), .B(new_n421), .C1(new_n415), .C2(new_n416), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n883), .B1(new_n421), .B2(new_n884), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n411), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n891), .A2(new_n895), .B1(KEYINPUT37), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n882), .B1(new_n886), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n382), .A2(new_n405), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT101), .B1(new_n901), .B2(new_n421), .ZN(new_n902));
  INV_X1    g0702(.A(new_n894), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n904), .B2(new_n890), .ZN(new_n905));
  INV_X1    g0705(.A(new_n885), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n413), .A2(new_n418), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n423), .A2(new_n425), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n899), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n342), .A2(new_n340), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n345), .A2(new_n346), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n336), .B1(new_n314), .B2(new_n319), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n336), .B(new_n661), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n336), .A2(new_n661), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n338), .B(new_n917), .C1(new_n347), .C2(new_n337), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n881), .A2(new_n911), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n888), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n908), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n411), .A2(new_n422), .A3(new_n889), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n904), .B2(new_n890), .ZN(new_n925));
  INV_X1    g0725(.A(new_n889), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n907), .B2(new_n908), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT103), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n899), .B(new_n910), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT39), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(new_n928), .ZN(new_n933));
  NOR2_X1   g0733(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n614), .A2(new_n662), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n922), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n461), .B(new_n739), .C1(KEYINPUT29), .C2(new_n743), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n621), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n940), .B(new_n942), .Z(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n720), .A2(new_n722), .A3(new_n725), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n838), .B1(new_n724), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n919), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n944), .B1(new_n948), .B2(new_n911), .ZN(new_n949));
  INV_X1    g0749(.A(new_n933), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n950), .A2(new_n946), .A3(KEYINPUT40), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n724), .A2(new_n945), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n461), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n690), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n943), .A2(new_n956), .B1(new_n206), .B2(new_n748), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n943), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n880), .B1(new_n957), .B2(new_n958), .ZN(G367));
  NAND2_X1  g0759(.A1(new_n234), .A2(new_n824), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n817), .B1(new_n818), .B2(new_n562), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n750), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n732), .A2(new_n662), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n630), .B2(new_n733), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n630), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n813), .A2(G137), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n772), .A2(G68), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n794), .A2(G143), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n777), .A2(new_n376), .B1(new_n785), .B2(new_n202), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n803), .A2(new_n247), .B1(new_n358), .B2(new_n781), .ZN(new_n970));
  INV_X1    g0770(.A(G150), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n268), .B1(new_n784), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n268), .B1(new_n798), .B2(G294), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n801), .B2(new_n784), .C1(new_n803), .C2(new_n556), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n776), .A2(G116), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT46), .Z(new_n978));
  AOI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(G311), .C2(new_n794), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n771), .A2(new_n267), .B1(new_n804), .B2(new_n785), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT105), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n979), .B(new_n981), .C1(new_n982), .C2(new_n766), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n980), .A2(KEYINPUT105), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n974), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT47), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n759), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n962), .B1(new_n965), .B2(new_n757), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n675), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n694), .B1(new_n523), .B2(new_n662), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n734), .A2(new_n661), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n993), .A2(new_n676), .A3(new_n662), .A4(new_n674), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n540), .B1(new_n991), .B2(new_n642), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n662), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n999), .A2(KEYINPUT43), .A3(new_n965), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT104), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n965), .B(KEYINPUT43), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  AND4_X1   g0803(.A1(new_n990), .A2(new_n1001), .A3(new_n993), .A4(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1001), .A2(new_n1003), .B1(new_n990), .B2(new_n993), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n749), .A2(G1), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n666), .A2(new_n672), .A3(new_n673), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n675), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n677), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1010), .A2(new_n678), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n683), .A2(new_n993), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT44), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n683), .A2(new_n993), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n990), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1013), .A2(new_n675), .A3(new_n1016), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1011), .A2(new_n1018), .A3(new_n746), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n746), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n685), .B(KEYINPUT41), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1007), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n989), .B1(new_n1006), .B2(new_n1024), .ZN(G387));
  XNOR2_X1  g0825(.A(new_n685), .B(KEYINPUT108), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1011), .A2(new_n746), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT109), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT109), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n1011), .B2(new_n746), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1029), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n674), .A2(new_n757), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n686), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n819), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(G107), .B2(new_n210), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n230), .A2(G45), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n259), .A2(new_n202), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT50), .Z(new_n1039));
  AOI211_X1 g0839(.A(G45), .B(new_n1034), .C1(G68), .C2(G77), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n825), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1036), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n753), .B1(new_n1042), .B2(new_n817), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n813), .A2(G150), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n772), .A2(new_n562), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n784), .A2(new_n202), .B1(new_n785), .B2(new_n330), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n268), .B1(new_n803), .B2(new_n556), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G77), .C2(new_n776), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n794), .A2(G159), .B1(new_n355), .B2(new_n798), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1044), .A2(new_n1045), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n268), .B1(new_n788), .B2(G116), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n784), .A2(new_n982), .B1(new_n785), .B2(new_n801), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT107), .Z(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n805), .B2(new_n781), .C1(new_n807), .C2(new_n793), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n772), .A2(G283), .B1(G294), .B2(new_n776), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT49), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1051), .B1(new_n811), .B2(new_n766), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1050), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1033), .B(new_n1043), .C1(new_n1063), .C2(new_n759), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1010), .A2(new_n678), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1007), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n1065), .A2(KEYINPUT106), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT106), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1032), .A2(new_n1069), .ZN(G393));
  OAI221_X1 g0870(.A(new_n816), .B1(new_n556), .B2(new_n210), .C1(new_n825), .C2(new_n241), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n753), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n848), .A2(new_n259), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n202), .B2(new_n781), .C1(new_n777), .C2(new_n330), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n372), .B(new_n1074), .C1(G87), .C2(new_n788), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n247), .B2(new_n771), .C1(new_n850), .C2(new_n766), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n793), .A2(new_n971), .B1(new_n358), .B2(new_n784), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  OAI22_X1  g0878(.A1(new_n793), .A2(new_n982), .B1(new_n805), .B2(new_n784), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT52), .Z(new_n1080));
  OAI21_X1  g0880(.A(new_n372), .B1(new_n803), .B2(new_n267), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n777), .A2(new_n804), .B1(new_n785), .B2(new_n810), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(G303), .C2(new_n798), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n491), .B2(new_n771), .C1(new_n807), .C2(new_n766), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1076), .A2(new_n1078), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1072), .B1(new_n1085), .B2(new_n759), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n757), .B2(new_n993), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1019), .A2(KEYINPUT110), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT110), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1013), .A2(new_n1016), .A3(new_n1089), .A4(new_n675), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1018), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1087), .B1(new_n1091), .B2(new_n1066), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1020), .A2(new_n1026), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n745), .B2(new_n1065), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(G390));
  INV_X1    g0896(.A(KEYINPUT114), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n937), .B1(new_n932), .B2(new_n928), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n730), .A2(new_n737), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n662), .A3(new_n837), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n919), .B1(new_n1100), .B2(new_n834), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n728), .A2(new_n841), .A3(new_n947), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n842), .A2(new_n834), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n938), .B1(new_n1105), .B2(new_n947), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1103), .B(new_n1104), .C1(new_n936), .C2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n930), .A2(KEYINPUT39), .B1(new_n933), .B2(new_n934), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n937), .B1(new_n881), .B2(new_n919), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1102), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n946), .A2(G330), .A3(new_n947), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1107), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n461), .A2(new_n953), .A3(G330), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n941), .A2(new_n621), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n833), .B1(new_n738), .B2(new_n837), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n720), .A2(new_n722), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n698), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1117), .A2(new_n661), .B1(new_n611), .B2(KEYINPUT31), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n727), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n841), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1115), .B1(new_n1120), .B2(new_n919), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n947), .B1(new_n946), .B2(G330), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n919), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n881), .B1(new_n1124), .B2(new_n1111), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1114), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT111), .B1(new_n1112), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1111), .B1(new_n1128), .B2(new_n1103), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT111), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n941), .A2(new_n621), .A3(new_n1113), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n945), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n841), .C1(new_n1118), .C2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n919), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n947), .B1(new_n728), .B2(new_n841), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1105), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n919), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n1104), .A3(new_n1115), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1132), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1130), .A2(new_n1131), .A3(new_n1140), .A4(new_n1107), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1127), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1027), .B1(new_n1112), .B2(new_n1126), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n869), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n753), .B1(new_n355), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n784), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G132), .A2(new_n1147), .B1(new_n798), .B2(G137), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1148), .B1(new_n785), .B2(new_n1149), .C1(new_n793), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n777), .A2(new_n971), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT53), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n268), .B1(new_n202), .B2(new_n803), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1151), .B(new_n1154), .C1(new_n1153), .C2(new_n1152), .ZN(new_n1155));
  INV_X1    g0955(.A(G125), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n766), .C1(new_n358), .C2(new_n771), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n781), .A2(new_n267), .B1(new_n785), .B2(new_n556), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n794), .B2(G283), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT112), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n268), .B(new_n855), .C1(G87), .C2(new_n776), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n810), .C2(new_n766), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n771), .A2(new_n247), .B1(new_n491), .B2(new_n784), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT113), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1157), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1146), .B1(new_n1165), .B2(new_n759), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n936), .B2(new_n755), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1112), .B2(new_n1066), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1097), .B1(new_n1144), .B2(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(KEYINPUT114), .B(new_n1168), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(G378));
  OAI22_X1  g0972(.A1(new_n781), .A2(new_n556), .B1(new_n785), .B2(new_n255), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n803), .A2(new_n376), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G107), .C2(new_n1147), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n372), .A2(new_n276), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n776), .B2(G77), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G116), .B2(new_n794), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(new_n967), .C1(new_n804), .C2(new_n766), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT58), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1176), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n784), .A2(new_n1150), .B1(new_n785), .B2(new_n851), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n777), .A2(new_n1149), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G132), .C2(new_n798), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n793), .B2(new_n1156), .C1(new_n971), .C2(new_n771), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n385), .B(new_n276), .C1(new_n803), .C2(new_n358), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n813), .B2(G124), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n759), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n750), .B1(new_n202), .B2(new_n869), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n460), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n445), .A2(new_n659), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT115), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n460), .A2(new_n1197), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1200), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1195), .B(new_n1196), .C1(new_n1204), .C2(new_n755), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n952), .B2(new_n690), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1204), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1208), .A2(new_n949), .A3(G330), .A4(new_n951), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n940), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n939), .A3(new_n1209), .A4(new_n922), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1206), .B1(new_n1214), .B2(new_n1007), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT116), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT57), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1132), .B1(new_n1127), .B2(new_n1141), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1216), .B(new_n1217), .C1(new_n1218), .C2(new_n1213), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1120), .A2(new_n919), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1102), .B(new_n1220), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1129), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1131), .B1(new_n1222), .B2(new_n1140), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1112), .A2(KEYINPUT111), .A3(new_n1126), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1114), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n1214), .A3(KEYINPUT57), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1219), .A2(new_n1226), .A3(new_n1026), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1214), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1216), .B1(new_n1228), .B2(new_n1217), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1215), .B1(new_n1227), .B2(new_n1229), .ZN(G375));
  XNOR2_X1  g1030(.A(new_n1007), .B(KEYINPUT118), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n919), .A2(new_n754), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n753), .B1(G68), .B2(new_n1145), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n777), .A2(new_n358), .B1(new_n785), .B2(new_n971), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n851), .A2(new_n784), .B1(new_n781), .B2(new_n1149), .ZN(new_n1236));
  OR4_X1    g1036(.A1(new_n372), .A2(new_n1235), .A3(new_n1174), .A4(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G132), .B2(new_n794), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n202), .B2(new_n771), .C1(new_n1150), .C2(new_n766), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n766), .A2(new_n801), .B1(new_n556), .B2(new_n777), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT119), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n794), .A2(G294), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n268), .B1(new_n788), .B2(G77), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n784), .A2(new_n804), .B1(new_n785), .B2(new_n267), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G116), .B2(new_n798), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1045), .A2(new_n1242), .A3(new_n1243), .A4(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1234), .B1(new_n1247), .B2(new_n759), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1233), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT120), .B1(new_n1232), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT120), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1252), .B(new_n1249), .C1(new_n1253), .C2(new_n1231), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1137), .A2(new_n1132), .A3(new_n1139), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT117), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n1132), .A4(new_n1139), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1258), .A2(new_n1023), .A3(new_n1126), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1255), .A2(new_n1260), .ZN(G381));
  AOI21_X1  g1061(.A(new_n1168), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n1215), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1032), .A2(new_n831), .A3(new_n1069), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(G384), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1095), .ZN(new_n1267));
  OR4_X1    g1067(.A1(G387), .A2(new_n1263), .A3(G381), .A4(new_n1267), .ZN(G407));
  OAI211_X1 g1068(.A(G407), .B(G213), .C1(G343), .C2(new_n1263), .ZN(G409));
  INV_X1    g1069(.A(KEYINPUT124), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(G387), .B2(new_n1095), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n831), .B1(new_n1032), .B2(new_n1069), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1265), .A2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1022), .B1(new_n1020), .B2(new_n746), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1007), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(G390), .A2(KEYINPUT124), .A3(new_n1276), .A4(new_n989), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G387), .A2(new_n1095), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1271), .A2(new_n1273), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(G390), .A2(new_n1276), .A3(new_n989), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1278), .A2(new_n1280), .A3(KEYINPUT125), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G387), .A2(new_n1282), .A3(new_n1095), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1265), .B2(new_n1272), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1279), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1215), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1225), .A2(new_n1023), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1213), .B1(new_n1287), .B2(new_n1231), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1262), .B1(new_n1288), .B2(new_n1206), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  INV_X1    g1091(.A(G213), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(G343), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1256), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1027), .B1(new_n1297), .B2(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1299), .A2(G384), .A3(new_n1255), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G384), .B1(new_n1299), .B2(new_n1255), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1290), .A2(new_n1291), .A3(new_n1294), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1255), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1266), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT122), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1299), .A2(G384), .A3(new_n1255), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT123), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1293), .A2(G2897), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1309), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT122), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1313), .A2(new_n1314), .A3(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1316), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1300), .A2(new_n1301), .A3(KEYINPUT122), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT123), .B1(new_n1319), .B2(new_n1311), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1309), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1317), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1293), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1303), .B(new_n1304), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1325));
  AOI211_X1 g1125(.A(new_n1293), .B(new_n1315), .C1(new_n1286), .C2(new_n1289), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(new_n1291), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1285), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1316), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1320), .A2(new_n1318), .A3(new_n1321), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1324), .A2(KEYINPUT121), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT121), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1334), .ZN(new_n1335));
  OR2_X1    g1135(.A1(new_n1326), .A2(KEYINPUT63), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1279), .B(new_n1304), .C1(new_n1281), .C2(new_n1284), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1337), .B1(new_n1326), .B2(KEYINPUT63), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1335), .A2(new_n1336), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1328), .A2(new_n1339), .ZN(G405));
  XNOR2_X1  g1140(.A(new_n1285), .B(new_n1302), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT126), .B1(G375), .B2(new_n1262), .ZN(new_n1342));
  AND3_X1   g1142(.A1(G375), .A2(KEYINPUT126), .A3(new_n1262), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1286), .ZN(new_n1344));
  OR2_X1    g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1341), .B1(new_n1342), .B2(new_n1345), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1285), .B(new_n1315), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1343), .A2(new_n1342), .A3(new_n1344), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1346), .A2(new_n1349), .ZN(G402));
endmodule


