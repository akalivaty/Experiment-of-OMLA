

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712;

  XNOR2_X1 U364 ( .A(n585), .B(n584), .ZN(n684) );
  INV_X1 U365 ( .A(n493), .ZN(n610) );
  XNOR2_X2 U366 ( .A(n390), .B(KEYINPUT19), .ZN(n544) );
  XNOR2_X1 U367 ( .A(n565), .B(n487), .ZN(n571) );
  NAND2_X1 U368 ( .A1(n576), .A2(n571), .ZN(n548) );
  NOR2_X2 U369 ( .A1(n632), .A2(n631), .ZN(n576) );
  XNOR2_X1 U370 ( .A(n383), .B(n382), .ZN(n526) );
  NOR2_X1 U371 ( .A1(n523), .A2(n504), .ZN(n501) );
  AND2_X1 U372 ( .A1(n565), .A2(n621), .ZN(n495) );
  OR2_X1 U373 ( .A1(n554), .A2(n634), .ZN(n631) );
  XNOR2_X1 U374 ( .A(n459), .B(n458), .ZN(n522) );
  XNOR2_X1 U375 ( .A(n361), .B(n360), .ZN(n634) );
  OR2_X1 U376 ( .A1(n663), .A2(G902), .ZN(n381) );
  NOR2_X1 U377 ( .A1(G902), .A2(n670), .ZN(n458) );
  XNOR2_X1 U378 ( .A(n358), .B(n453), .ZN(n464) );
  XNOR2_X2 U379 ( .A(n399), .B(KEYINPUT69), .ZN(n420) );
  XNOR2_X2 U380 ( .A(G101), .B(KEYINPUT68), .ZN(n399) );
  NAND2_X1 U381 ( .A1(n711), .A2(n712), .ZN(n363) );
  XOR2_X1 U382 ( .A(n429), .B(n693), .Z(n484) );
  BUF_X1 U383 ( .A(n452), .Z(n589) );
  INV_X1 U384 ( .A(KEYINPUT78), .ZN(n382) );
  NOR2_X1 U385 ( .A1(n626), .A2(KEYINPUT47), .ZN(n383) );
  XNOR2_X1 U386 ( .A(n478), .B(n477), .ZN(n635) );
  NAND2_X1 U387 ( .A1(n424), .A2(n423), .ZN(n438) );
  INV_X1 U388 ( .A(G131), .ZN(n421) );
  NOR2_X1 U389 ( .A1(G953), .A2(G237), .ZN(n480) );
  OR2_X1 U390 ( .A1(n613), .A2(n600), .ZN(n370) );
  NOR2_X1 U391 ( .A1(n709), .A2(n394), .ZN(n393) );
  NAND2_X1 U392 ( .A1(n388), .A2(n344), .ZN(n387) );
  XNOR2_X1 U393 ( .A(n363), .B(n350), .ZN(n388) );
  XNOR2_X1 U394 ( .A(n482), .B(n391), .ZN(n677) );
  XNOR2_X1 U395 ( .A(n417), .B(n411), .ZN(n391) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n453) );
  NAND2_X1 U397 ( .A1(n452), .A2(G234), .ZN(n358) );
  XOR2_X1 U398 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n449) );
  XNOR2_X1 U399 ( .A(G134), .B(G122), .ZN(n448) );
  XNOR2_X1 U400 ( .A(G116), .B(G107), .ZN(n446) );
  XNOR2_X1 U401 ( .A(n362), .B(KEYINPUT25), .ZN(n361) );
  NOR2_X1 U402 ( .A1(n672), .A2(G902), .ZN(n360) );
  AND2_X1 U403 ( .A1(n476), .A2(G217), .ZN(n362) );
  XNOR2_X1 U404 ( .A(KEYINPUT6), .B(KEYINPUT101), .ZN(n487) );
  XNOR2_X1 U405 ( .A(n558), .B(n557), .ZN(n559) );
  INV_X1 U406 ( .A(KEYINPUT66), .ZN(n557) );
  XNOR2_X1 U407 ( .A(n484), .B(n430), .ZN(n663) );
  XNOR2_X1 U408 ( .A(n514), .B(n384), .ZN(n626) );
  INV_X1 U409 ( .A(KEYINPUT99), .ZN(n384) );
  XNOR2_X1 U410 ( .A(G116), .B(G113), .ZN(n408) );
  INV_X1 U411 ( .A(KEYINPUT71), .ZN(n422) );
  INV_X1 U412 ( .A(KEYINPUT44), .ZN(n394) );
  XNOR2_X1 U413 ( .A(n367), .B(KEYINPUT86), .ZN(n400) );
  XNOR2_X1 U414 ( .A(n392), .B(n409), .ZN(n482) );
  XOR2_X1 U415 ( .A(KEYINPUT74), .B(G119), .Z(n409) );
  XNOR2_X1 U416 ( .A(n408), .B(n407), .ZN(n392) );
  INV_X1 U417 ( .A(KEYINPUT3), .ZN(n407) );
  XNOR2_X1 U418 ( .A(n428), .B(n427), .ZN(n693) );
  XOR2_X1 U419 ( .A(G134), .B(G137), .Z(n425) );
  XNOR2_X1 U420 ( .A(n359), .B(G953), .ZN(n452) );
  INV_X1 U421 ( .A(KEYINPUT64), .ZN(n359) );
  NAND2_X1 U422 ( .A1(G234), .A2(G237), .ZN(n470) );
  XNOR2_X1 U423 ( .A(KEYINPUT85), .B(KEYINPUT33), .ZN(n547) );
  XNOR2_X1 U424 ( .A(KEYINPUT20), .B(n469), .ZN(n476) );
  INV_X1 U425 ( .A(G469), .ZN(n380) );
  XNOR2_X1 U426 ( .A(G119), .B(G110), .ZN(n461) );
  XNOR2_X1 U427 ( .A(G128), .B(G137), .ZN(n460) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(G140), .Z(n432) );
  XNOR2_X1 U429 ( .A(G104), .B(G122), .ZN(n431) );
  INV_X1 U430 ( .A(KEYINPUT10), .ZN(n389) );
  XNOR2_X1 U431 ( .A(G113), .B(G143), .ZN(n437) );
  XOR2_X1 U432 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n434) );
  INV_X1 U433 ( .A(KEYINPUT45), .ZN(n584) );
  NOR2_X1 U434 ( .A1(n620), .A2(n386), .ZN(n385) );
  INV_X1 U435 ( .A(n619), .ZN(n386) );
  XNOR2_X1 U436 ( .A(G104), .B(G110), .ZN(n410) );
  XOR2_X1 U437 ( .A(G140), .B(KEYINPUT72), .Z(n467) );
  NOR2_X1 U438 ( .A1(n578), .A2(n497), .ZN(n499) );
  INV_X1 U439 ( .A(G475), .ZN(n444) );
  XNOR2_X1 U440 ( .A(n457), .B(n456), .ZN(n670) );
  XNOR2_X1 U441 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U442 ( .A(n379), .B(n588), .ZN(n378) );
  INV_X1 U443 ( .A(G953), .ZN(n698) );
  XNOR2_X1 U444 ( .A(n502), .B(n503), .ZN(n711) );
  AND2_X1 U445 ( .A1(n610), .A2(n539), .ZN(n502) );
  NOR2_X1 U446 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U447 ( .A(n570), .B(KEYINPUT102), .ZN(n708) );
  AND2_X1 U448 ( .A1(n371), .A2(n566), .ZN(n600) );
  NOR2_X1 U449 ( .A1(n595), .A2(n676), .ZN(n597) );
  NOR2_X1 U450 ( .A1(n667), .A2(n676), .ZN(n668) );
  AND2_X1 U451 ( .A1(n364), .A2(n590), .ZN(G54) );
  XNOR2_X1 U452 ( .A(n366), .B(n365), .ZN(n364) );
  XNOR2_X1 U453 ( .A(n663), .B(n355), .ZN(n365) );
  AND2_X1 U454 ( .A1(n537), .A2(n618), .ZN(n344) );
  XOR2_X1 U455 ( .A(n481), .B(KEYINPUT5), .Z(n345) );
  XOR2_X1 U456 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n346) );
  AND2_X1 U457 ( .A1(G210), .A2(n489), .ZN(n347) );
  AND2_X1 U458 ( .A1(n370), .A2(n519), .ZN(n348) );
  XOR2_X1 U459 ( .A(KEYINPUT67), .B(KEYINPUT1), .Z(n349) );
  XNOR2_X1 U460 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n350) );
  AND2_X1 U461 ( .A1(n395), .A2(G475), .ZN(n351) );
  AND2_X1 U462 ( .A1(n395), .A2(G472), .ZN(n352) );
  AND2_X1 U463 ( .A1(n395), .A2(G469), .ZN(n353) );
  AND2_X1 U464 ( .A1(n395), .A2(G210), .ZN(n354) );
  NOR2_X1 U465 ( .A1(n589), .A2(G952), .ZN(n676) );
  XNOR2_X1 U466 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n355) );
  XOR2_X1 U467 ( .A(n591), .B(KEYINPUT56), .Z(n356) );
  XNOR2_X1 U468 ( .A(n501), .B(n500), .ZN(n539) );
  NAND2_X1 U469 ( .A1(n357), .A2(n385), .ZN(n700) );
  XNOR2_X1 U470 ( .A(n387), .B(n538), .ZN(n357) );
  NAND2_X1 U471 ( .A1(n368), .A2(n353), .ZN(n366) );
  XNOR2_X1 U472 ( .A(n367), .B(n389), .ZN(n466) );
  XNOR2_X2 U473 ( .A(G146), .B(G125), .ZN(n367) );
  NAND2_X1 U474 ( .A1(n368), .A2(n351), .ZN(n665) );
  NAND2_X1 U475 ( .A1(n368), .A2(n352), .ZN(n594) );
  NAND2_X1 U476 ( .A1(n368), .A2(n354), .ZN(n379) );
  AND2_X1 U477 ( .A1(n368), .A2(n395), .ZN(n396) );
  XNOR2_X1 U478 ( .A(n368), .B(KEYINPUT82), .ZN(n659) );
  XNOR2_X2 U479 ( .A(n586), .B(n369), .ZN(n368) );
  INV_X1 U480 ( .A(KEYINPUT2), .ZN(n369) );
  XNOR2_X1 U481 ( .A(n580), .B(KEYINPUT92), .ZN(n371) );
  NAND2_X1 U482 ( .A1(n376), .A2(n372), .ZN(n375) );
  INV_X1 U483 ( .A(n709), .ZN(n372) );
  XNOR2_X2 U484 ( .A(n553), .B(KEYINPUT35), .ZN(n709) );
  AND2_X2 U485 ( .A1(n707), .A2(n708), .ZN(n376) );
  NAND2_X1 U486 ( .A1(n374), .A2(n373), .ZN(n583) );
  NAND2_X1 U487 ( .A1(n393), .A2(n376), .ZN(n373) );
  NAND2_X1 U488 ( .A1(n375), .A2(n394), .ZN(n374) );
  XNOR2_X1 U489 ( .A(n377), .B(n356), .ZN(G51) );
  NAND2_X1 U490 ( .A1(n378), .A2(n590), .ZN(n377) );
  XNOR2_X2 U491 ( .A(n508), .B(n349), .ZN(n632) );
  XNOR2_X2 U492 ( .A(n381), .B(n380), .ZN(n508) );
  XNOR2_X1 U493 ( .A(n400), .B(n420), .ZN(n401) );
  XNOR2_X1 U494 ( .A(n548), .B(n547), .ZN(n652) );
  XNOR2_X1 U495 ( .A(n402), .B(n401), .ZN(n406) );
  NAND2_X1 U496 ( .A1(n544), .A2(n545), .ZN(n546) );
  NAND2_X1 U497 ( .A1(n516), .A2(n621), .ZN(n390) );
  XNOR2_X2 U498 ( .A(n416), .B(n347), .ZN(n516) );
  XNOR2_X2 U499 ( .A(n563), .B(KEYINPUT32), .ZN(n707) );
  INV_X1 U500 ( .A(n587), .ZN(n395) );
  NAND2_X1 U501 ( .A1(n396), .A2(G478), .ZN(n669) );
  NAND2_X1 U502 ( .A1(n396), .A2(G217), .ZN(n673) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n513) );
  XNOR2_X1 U504 ( .A(n406), .B(n405), .ZN(n412) );
  XOR2_X1 U505 ( .A(n463), .B(n462), .Z(n397) );
  AND2_X1 U506 ( .A1(n498), .A2(n479), .ZN(n398) );
  INV_X1 U507 ( .A(KEYINPUT48), .ZN(n538) );
  XNOR2_X1 U508 ( .A(n482), .B(n345), .ZN(n483) );
  NOR2_X1 U509 ( .A1(n579), .A2(n652), .ZN(n550) );
  XNOR2_X1 U510 ( .A(n484), .B(n483), .ZN(n592) );
  XNOR2_X1 U511 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XOR2_X1 U512 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n414) );
  XOR2_X1 U513 ( .A(G143), .B(G128), .Z(n447) );
  XNOR2_X1 U514 ( .A(KEYINPUT4), .B(n447), .ZN(n427) );
  INV_X1 U515 ( .A(n427), .ZN(n402) );
  XOR2_X1 U516 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n404) );
  NAND2_X1 U517 ( .A1(G224), .A2(n589), .ZN(n403) );
  XNOR2_X1 U518 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U519 ( .A(G122), .B(KEYINPUT16), .Z(n411) );
  XNOR2_X1 U520 ( .A(n410), .B(G107), .ZN(n417) );
  XNOR2_X1 U521 ( .A(n412), .B(n677), .ZN(n415) );
  XNOR2_X1 U522 ( .A(n415), .B(KEYINPUT84), .ZN(n413) );
  XNOR2_X1 U523 ( .A(n414), .B(n413), .ZN(n588) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n587) );
  NAND2_X1 U525 ( .A1(n415), .A2(n587), .ZN(n416) );
  OR2_X1 U526 ( .A1(G237), .A2(G902), .ZN(n489) );
  XOR2_X1 U527 ( .A(n467), .B(n417), .Z(n419) );
  NAND2_X1 U528 ( .A1(G227), .A2(n589), .ZN(n418) );
  XNOR2_X1 U529 ( .A(n419), .B(n418), .ZN(n430) );
  XNOR2_X1 U530 ( .A(G146), .B(n420), .ZN(n429) );
  NAND2_X1 U531 ( .A1(KEYINPUT71), .A2(n421), .ZN(n424) );
  NAND2_X1 U532 ( .A1(n422), .A2(G131), .ZN(n423) );
  XNOR2_X1 U533 ( .A(n438), .B(KEYINPUT73), .ZN(n426) );
  XNOR2_X1 U534 ( .A(n426), .B(n425), .ZN(n428) );
  INV_X1 U535 ( .A(n632), .ZN(n567) );
  XNOR2_X1 U536 ( .A(KEYINPUT13), .B(KEYINPUT95), .ZN(n443) );
  XNOR2_X1 U537 ( .A(n432), .B(n431), .ZN(n436) );
  NAND2_X1 U538 ( .A1(G214), .A2(n480), .ZN(n433) );
  XNOR2_X1 U539 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U540 ( .A(n436), .B(n435), .ZN(n441) );
  XNOR2_X1 U541 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n466), .B(n439), .ZN(n440) );
  XNOR2_X1 U543 ( .A(n441), .B(n440), .ZN(n664) );
  NOR2_X1 U544 ( .A1(G902), .A2(n664), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U546 ( .A(KEYINPUT98), .B(G478), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n447), .B(n446), .ZN(n451) );
  XNOR2_X1 U548 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U549 ( .A(n451), .B(n450), .Z(n457) );
  NAND2_X1 U550 ( .A1(G217), .A2(n464), .ZN(n455) );
  XNOR2_X1 U551 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n454) );
  NAND2_X1 U552 ( .A1(n513), .A2(n522), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n460), .B(KEYINPUT24), .ZN(n463) );
  XNOR2_X1 U554 ( .A(n346), .B(n461), .ZN(n462) );
  NAND2_X1 U555 ( .A1(G221), .A2(n464), .ZN(n465) );
  XNOR2_X1 U556 ( .A(n397), .B(n465), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n467), .B(n466), .ZN(n692) );
  XNOR2_X1 U558 ( .A(n468), .B(n692), .ZN(n672) );
  NAND2_X1 U559 ( .A1(G234), .A2(n587), .ZN(n469) );
  XNOR2_X1 U560 ( .A(n470), .B(KEYINPUT14), .ZN(n472) );
  NAND2_X1 U561 ( .A1(G952), .A2(n472), .ZN(n471) );
  XOR2_X1 U562 ( .A(KEYINPUT87), .B(n471), .Z(n651) );
  NOR2_X1 U563 ( .A1(G953), .A2(n651), .ZN(n540) );
  INV_X1 U564 ( .A(n589), .ZN(n703) );
  AND2_X1 U565 ( .A1(G902), .A2(n472), .ZN(n541) );
  NAND2_X1 U566 ( .A1(n703), .A2(n541), .ZN(n473) );
  NOR2_X1 U567 ( .A1(G900), .A2(n473), .ZN(n474) );
  NOR2_X1 U568 ( .A1(n540), .A2(n474), .ZN(n475) );
  XNOR2_X1 U569 ( .A(KEYINPUT81), .B(n475), .ZN(n498) );
  XOR2_X1 U570 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n478) );
  NAND2_X1 U571 ( .A1(n476), .A2(G221), .ZN(n477) );
  INV_X1 U572 ( .A(n635), .ZN(n479) );
  AND2_X1 U573 ( .A1(n634), .A2(n398), .ZN(n506) );
  NAND2_X1 U574 ( .A1(n480), .A2(G210), .ZN(n481) );
  NOR2_X1 U575 ( .A1(n592), .A2(G902), .ZN(n486) );
  XNOR2_X1 U576 ( .A(G472), .B(KEYINPUT93), .ZN(n485) );
  XNOR2_X2 U577 ( .A(n486), .B(n485), .ZN(n565) );
  NAND2_X1 U578 ( .A1(n506), .A2(n571), .ZN(n488) );
  NOR2_X1 U579 ( .A1(n493), .A2(n488), .ZN(n490) );
  NAND2_X1 U580 ( .A1(G214), .A2(n489), .ZN(n621) );
  NAND2_X1 U581 ( .A1(n490), .A2(n621), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n567), .A2(n532), .ZN(n491) );
  XNOR2_X1 U583 ( .A(n491), .B(KEYINPUT43), .ZN(n492) );
  NOR2_X1 U584 ( .A1(n516), .A2(n492), .ZN(n620) );
  INV_X1 U585 ( .A(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U586 ( .A(n635), .B(KEYINPUT90), .ZN(n554) );
  NOR2_X1 U587 ( .A1(n631), .A2(n508), .ZN(n494) );
  XNOR2_X1 U588 ( .A(n494), .B(KEYINPUT91), .ZN(n578) );
  INV_X1 U589 ( .A(KEYINPUT30), .ZN(n496) );
  XNOR2_X1 U590 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U591 ( .A1(n499), .A2(n498), .ZN(n523) );
  INV_X1 U592 ( .A(n516), .ZN(n531) );
  XOR2_X1 U593 ( .A(KEYINPUT38), .B(n531), .Z(n504) );
  INV_X1 U594 ( .A(KEYINPUT39), .ZN(n500) );
  INV_X1 U595 ( .A(n504), .ZN(n622) );
  NAND2_X1 U596 ( .A1(n622), .A2(n621), .ZN(n625) );
  INV_X1 U597 ( .A(n513), .ZN(n521) );
  NAND2_X1 U598 ( .A1(n522), .A2(n521), .ZN(n624) );
  NOR2_X1 U599 ( .A1(n625), .A2(n624), .ZN(n505) );
  XNOR2_X1 U600 ( .A(KEYINPUT41), .B(n505), .ZN(n653) );
  AND2_X1 U601 ( .A1(n506), .A2(n565), .ZN(n507) );
  XNOR2_X1 U602 ( .A(KEYINPUT28), .B(n507), .ZN(n510) );
  INV_X1 U603 ( .A(n508), .ZN(n509) );
  NAND2_X1 U604 ( .A1(n510), .A2(n509), .ZN(n515) );
  NOR2_X1 U605 ( .A1(n653), .A2(n515), .ZN(n512) );
  XNOR2_X1 U606 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U607 ( .A(n512), .B(n511), .ZN(n712) );
  NOR2_X1 U608 ( .A1(n513), .A2(n522), .ZN(n612) );
  NOR2_X1 U609 ( .A1(n610), .A2(n612), .ZN(n514) );
  INV_X1 U610 ( .A(n626), .ZN(n519) );
  INV_X1 U611 ( .A(n515), .ZN(n517) );
  NAND2_X1 U612 ( .A1(n517), .A2(n544), .ZN(n605) );
  INV_X1 U613 ( .A(n605), .ZN(n518) );
  NAND2_X1 U614 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U615 ( .A1(n520), .A2(KEYINPUT47), .ZN(n525) );
  NOR2_X1 U616 ( .A1(n522), .A2(n521), .ZN(n551) );
  NOR2_X1 U617 ( .A1(n531), .A2(n523), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n551), .A2(n524), .ZN(n608) );
  NAND2_X1 U619 ( .A1(n525), .A2(n608), .ZN(n529) );
  NOR2_X1 U620 ( .A1(n605), .A2(n526), .ZN(n527) );
  XOR2_X1 U621 ( .A(KEYINPUT77), .B(n527), .Z(n528) );
  NOR2_X1 U622 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U623 ( .A(n530), .B(KEYINPUT76), .ZN(n537) );
  OR2_X1 U624 ( .A1(n532), .A2(n531), .ZN(n535) );
  XNOR2_X1 U625 ( .A(KEYINPUT104), .B(KEYINPUT36), .ZN(n533) );
  XNOR2_X1 U626 ( .A(n533), .B(KEYINPUT83), .ZN(n534) );
  XNOR2_X1 U627 ( .A(n535), .B(n534), .ZN(n536) );
  NAND2_X1 U628 ( .A1(n536), .A2(n567), .ZN(n618) );
  NAND2_X1 U629 ( .A1(n539), .A2(n612), .ZN(n619) );
  INV_X1 U630 ( .A(n540), .ZN(n543) );
  NOR2_X1 U631 ( .A1(G898), .A2(n698), .ZN(n679) );
  NAND2_X1 U632 ( .A1(n541), .A2(n679), .ZN(n542) );
  NAND2_X1 U633 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X2 U634 ( .A(n546), .B(KEYINPUT0), .ZN(n579) );
  XOR2_X1 U635 ( .A(KEYINPUT34), .B(KEYINPUT79), .Z(n549) );
  XNOR2_X1 U636 ( .A(n550), .B(n549), .ZN(n552) );
  NAND2_X1 U637 ( .A1(n552), .A2(n551), .ZN(n553) );
  INV_X1 U638 ( .A(n624), .ZN(n556) );
  NOR2_X1 U639 ( .A1(n579), .A2(n554), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n556), .A2(n555), .ZN(n560) );
  XOR2_X1 U641 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n558) );
  XNOR2_X2 U642 ( .A(n560), .B(n559), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n634), .A2(n573), .ZN(n564) );
  XNOR2_X1 U644 ( .A(KEYINPUT80), .B(n571), .ZN(n561) );
  NAND2_X1 U645 ( .A1(n567), .A2(n562), .ZN(n563) );
  INV_X1 U646 ( .A(n564), .ZN(n569) );
  INV_X1 U647 ( .A(n565), .ZN(n566) );
  NOR2_X1 U648 ( .A1(n567), .A2(n565), .ZN(n568) );
  NAND2_X1 U649 ( .A1(n569), .A2(n568), .ZN(n570) );
  INV_X1 U650 ( .A(n571), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U652 ( .A1(n634), .A2(n574), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n632), .A2(n575), .ZN(n598) );
  NAND2_X1 U654 ( .A1(n565), .A2(n576), .ZN(n642) );
  NOR2_X1 U655 ( .A1(n579), .A2(n642), .ZN(n577) );
  XOR2_X1 U656 ( .A(KEYINPUT31), .B(n577), .Z(n613) );
  NOR2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U658 ( .A(KEYINPUT100), .B(n348), .Z(n581) );
  AND2_X1 U659 ( .A1(n598), .A2(n581), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n585) );
  NOR2_X2 U661 ( .A1(n700), .A2(n684), .ZN(n586) );
  INV_X1 U662 ( .A(n676), .ZN(n590) );
  INV_X1 U663 ( .A(KEYINPUT115), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n594), .B(n593), .ZN(n595) );
  INV_X1 U665 ( .A(KEYINPUT63), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n597), .B(n596), .ZN(G57) );
  XNOR2_X1 U667 ( .A(G101), .B(n598), .ZN(G3) );
  NAND2_X1 U668 ( .A1(n600), .A2(n610), .ZN(n599) );
  XNOR2_X1 U669 ( .A(n599), .B(G104), .ZN(G6) );
  XOR2_X1 U670 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n602) );
  NAND2_X1 U671 ( .A1(n600), .A2(n612), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(n604) );
  XOR2_X1 U673 ( .A(G107), .B(KEYINPUT105), .Z(n603) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(G9) );
  XOR2_X1 U675 ( .A(G128), .B(KEYINPUT29), .Z(n607) );
  NAND2_X1 U676 ( .A1(n518), .A2(n612), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(G30) );
  XNOR2_X1 U678 ( .A(G143), .B(n608), .ZN(G45) );
  NAND2_X1 U679 ( .A1(n518), .A2(n610), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(G146), .ZN(G48) );
  NAND2_X1 U681 ( .A1(n613), .A2(n610), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(G113), .ZN(G15) );
  XOR2_X1 U683 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n615) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U686 ( .A(G116), .B(n616), .ZN(G18) );
  XOR2_X1 U687 ( .A(G125), .B(KEYINPUT37), .Z(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(G27) );
  XNOR2_X1 U689 ( .A(G134), .B(n619), .ZN(G36) );
  XOR2_X1 U690 ( .A(G140), .B(n620), .Z(G42) );
  XOR2_X1 U691 ( .A(KEYINPUT114), .B(KEYINPUT53), .Z(n662) );
  NOR2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n628) );
  NOR2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U695 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U696 ( .A1(n629), .A2(n652), .ZN(n630) );
  XNOR2_X1 U697 ( .A(n630), .B(KEYINPUT110), .ZN(n647) );
  NAND2_X1 U698 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U699 ( .A(n633), .B(KEYINPUT50), .ZN(n641) );
  XOR2_X1 U700 ( .A(KEYINPUT49), .B(KEYINPUT108), .Z(n637) );
  NAND2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U702 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U703 ( .A1(n638), .A2(n566), .ZN(n639) );
  XNOR2_X1 U704 ( .A(KEYINPUT109), .B(n639), .ZN(n640) );
  NAND2_X1 U705 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U706 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U707 ( .A(KEYINPUT51), .B(n644), .ZN(n645) );
  NOR2_X1 U708 ( .A1(n653), .A2(n645), .ZN(n646) );
  NOR2_X1 U709 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U710 ( .A(n648), .B(KEYINPUT52), .Z(n649) );
  XNOR2_X1 U711 ( .A(KEYINPUT111), .B(n649), .ZN(n650) );
  NOR2_X1 U712 ( .A1(n651), .A2(n650), .ZN(n656) );
  NOR2_X1 U713 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U714 ( .A(n654), .B(KEYINPUT112), .ZN(n655) );
  NOR2_X1 U715 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U716 ( .A(n657), .B(KEYINPUT113), .ZN(n658) );
  NOR2_X1 U717 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U718 ( .A1(n660), .A2(n698), .ZN(n661) );
  XNOR2_X1 U719 ( .A(n662), .B(n661), .ZN(G75) );
  XOR2_X1 U720 ( .A(n664), .B(KEYINPUT59), .Z(n666) );
  XNOR2_X1 U721 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U722 ( .A(n668), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U723 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U724 ( .A1(n676), .A2(n671), .ZN(G63) );
  XNOR2_X1 U725 ( .A(n672), .B(KEYINPUT116), .ZN(n674) );
  XNOR2_X1 U726 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U727 ( .A1(n676), .A2(n675), .ZN(G66) );
  XNOR2_X1 U728 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n691) );
  XNOR2_X1 U729 ( .A(G101), .B(n677), .ZN(n678) );
  XNOR2_X1 U730 ( .A(n678), .B(KEYINPUT119), .ZN(n680) );
  NOR2_X1 U731 ( .A1(n680), .A2(n679), .ZN(n689) );
  NAND2_X1 U732 ( .A1(G953), .A2(G224), .ZN(n681) );
  XNOR2_X1 U733 ( .A(KEYINPUT61), .B(n681), .ZN(n682) );
  NAND2_X1 U734 ( .A1(n682), .A2(G898), .ZN(n683) );
  XNOR2_X1 U735 ( .A(KEYINPUT117), .B(n683), .ZN(n687) );
  NOR2_X1 U736 ( .A1(G953), .A2(n684), .ZN(n685) );
  XNOR2_X1 U737 ( .A(n685), .B(KEYINPUT118), .ZN(n686) );
  NOR2_X1 U738 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U739 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U740 ( .A(n691), .B(n690), .ZN(G69) );
  XOR2_X1 U741 ( .A(n693), .B(n692), .Z(n699) );
  XNOR2_X1 U742 ( .A(G227), .B(n699), .ZN(n694) );
  XNOR2_X1 U743 ( .A(n694), .B(KEYINPUT123), .ZN(n695) );
  NAND2_X1 U744 ( .A1(G900), .A2(n695), .ZN(n696) );
  XOR2_X1 U745 ( .A(KEYINPUT124), .B(n696), .Z(n697) );
  NOR2_X1 U746 ( .A1(n698), .A2(n697), .ZN(n705) );
  XNOR2_X1 U747 ( .A(n699), .B(KEYINPUT122), .ZN(n701) );
  XNOR2_X1 U748 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U749 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U750 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U751 ( .A(KEYINPUT125), .B(n706), .ZN(G72) );
  XNOR2_X1 U752 ( .A(G119), .B(n707), .ZN(G21) );
  XNOR2_X1 U753 ( .A(G110), .B(n708), .ZN(G12) );
  XOR2_X1 U754 ( .A(n709), .B(G122), .Z(n710) );
  XNOR2_X1 U755 ( .A(KEYINPUT126), .B(n710), .ZN(G24) );
  XNOR2_X1 U756 ( .A(G131), .B(n711), .ZN(G33) );
  XNOR2_X1 U757 ( .A(G137), .B(n712), .ZN(G39) );
endmodule

