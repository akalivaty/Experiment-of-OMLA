//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G131), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G134), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT64), .A3(G137), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT11), .B1(new_n194), .B2(G134), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n192), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n196), .B2(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n195), .A2(new_n204), .A3(new_n197), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(new_n191), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G143), .B(G146), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT76), .A3(new_n223), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(G128), .B1(new_n225), .B2(new_n227), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n226), .A2(KEYINPUT1), .A3(G146), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n221), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n228), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT66), .B1(new_n234), .B2(new_n235), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n224), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n241), .B(new_n242), .C1(new_n231), .C2(G128), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n217), .A2(new_n220), .A3(KEYINPUT10), .ZN(new_n245));
  OAI22_X1  g059(.A1(new_n237), .A2(KEYINPUT10), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G101), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n226), .A2(G146), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT0), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(new_n222), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  OAI22_X1  g067(.A1(new_n250), .A2(new_n240), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n225), .B(new_n227), .C1(new_n251), .C2(new_n222), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n257));
  NAND3_X1  g071(.A1(new_n247), .A2(G101), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n249), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n209), .B1(new_n246), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n198), .A2(new_n201), .A3(new_n192), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n206), .A2(new_n191), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n262), .A2(KEYINPUT77), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT77), .B1(new_n262), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n241), .B1(new_n231), .B2(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n230), .B2(new_n232), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n269), .B2(new_n221), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n222), .B1(new_n250), .B2(new_n240), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n242), .B1(new_n271), .B2(new_n241), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n234), .A2(KEYINPUT66), .A3(new_n235), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n228), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n245), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n266), .A2(new_n259), .A3(new_n270), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n261), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(G110), .B(G140), .Z(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT74), .ZN(new_n280));
  INV_X1    g094(.A(G227), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G953), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n280), .B(new_n282), .Z(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n283), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n239), .A2(new_n243), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n228), .A3(new_n221), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT76), .B1(new_n231), .B2(new_n223), .ZN(new_n288));
  AND4_X1   g102(.A1(KEYINPUT76), .A2(new_n223), .A3(new_n225), .A4(new_n227), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n236), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n217), .A2(new_n220), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n208), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(KEYINPUT12), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT12), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n295), .B(new_n208), .C1(new_n287), .C2(new_n292), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n285), .B(new_n277), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n284), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n189), .B1(new_n298), .B2(new_n187), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n277), .B1(new_n294), .B2(new_n296), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n283), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n285), .A2(new_n277), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n261), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n246), .A2(new_n260), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n283), .B1(new_n305), .B2(new_n266), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(KEYINPUT78), .ZN(new_n307));
  OAI211_X1 g121(.A(G469), .B(new_n301), .C1(new_n304), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  OAI21_X1  g124(.A(G221), .B1(new_n310), .B2(G902), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g126(.A1(KEYINPUT91), .A2(G952), .ZN(new_n313));
  NAND2_X1  g127(.A1(KEYINPUT91), .A2(G952), .ZN(new_n314));
  AOI21_X1  g128(.A(G953), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(G234), .A2(G237), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n317), .A2(KEYINPUT92), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(KEYINPUT92), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT21), .B(G898), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n316), .A2(G902), .A3(G953), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT93), .Z(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT2), .B(G113), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G116), .B(G119), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n329), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n249), .A2(new_n333), .A3(new_n258), .ZN(new_n334));
  INV_X1    g148(.A(G113), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n336));
  INV_X1    g150(.A(G116), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G119), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT79), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT5), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n329), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  AND4_X1   g160(.A1(KEYINPUT80), .A2(new_n291), .A3(new_n346), .A4(new_n330), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n339), .A2(new_n345), .B1(new_n329), .B2(new_n328), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT80), .B1(new_n348), .B2(new_n291), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n334), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G122), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n334), .B(new_n351), .C1(new_n347), .C2(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT0), .B(G128), .Z(new_n356));
  OAI211_X1 g170(.A(new_n255), .B(G125), .C1(new_n356), .C2(new_n231), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT81), .ZN(new_n358));
  INV_X1    g172(.A(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n244), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT82), .B(G224), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(G953), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n361), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n350), .A2(new_n365), .A3(new_n352), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n355), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n363), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n360), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(KEYINPUT7), .ZN(new_n370));
  AOI211_X1 g184(.A(G125), .B(new_n238), .C1(new_n239), .C2(new_n243), .ZN(new_n371));
  INV_X1    g185(.A(new_n357), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n351), .B(KEYINPUT8), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n339), .B1(new_n340), .B2(new_n331), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n375), .A2(new_n330), .A3(new_n291), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n348), .A2(new_n291), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n354), .A2(new_n369), .A3(new_n373), .A4(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n379), .A2(new_n188), .ZN(new_n380));
  OAI21_X1  g194(.A(G210), .B1(G237), .B2(G902), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n367), .B2(new_n380), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n325), .B(new_n326), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n386));
  XNOR2_X1  g200(.A(G113), .B(G122), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(new_n210), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G214), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n390), .A2(G237), .A3(G953), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT83), .B1(new_n391), .B2(G143), .ZN(new_n392));
  NOR2_X1   g206(.A1(G237), .A2(G953), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G214), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n226), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n392), .A2(new_n396), .B1(G143), .B2(new_n391), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT84), .ZN(new_n399));
  INV_X1    g213(.A(G140), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n359), .B2(KEYINPUT72), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(G125), .A3(G140), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(G146), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(G125), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n359), .A2(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n224), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n397), .A2(new_n399), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n391), .A2(G143), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n391), .A2(KEYINPUT83), .A3(G143), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n395), .B1(new_n394), .B2(new_n226), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT18), .A3(G131), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n403), .ZN(new_n415));
  AOI21_X1  g229(.A(G140), .B1(new_n402), .B2(G125), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT16), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n405), .A2(KEYINPUT16), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(G146), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT19), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n401), .B2(new_n403), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT19), .B1(new_n405), .B2(new_n406), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n224), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n412), .A2(G131), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n397), .A2(new_n190), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n389), .B1(new_n414), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n408), .A2(new_n413), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT17), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n426), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT16), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n401), .B2(new_n403), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n224), .B1(new_n434), .B2(new_n418), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n420), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n412), .A2(KEYINPUT17), .A3(G131), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n388), .B(new_n430), .C1(new_n432), .C2(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n429), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g254(.A1(G475), .A2(G902), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n386), .B(KEYINPUT20), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n429), .B2(new_n439), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT85), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n444), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n337), .A2(G122), .ZN(new_n448));
  INV_X1    g262(.A(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n450), .A3(new_n213), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT89), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G128), .B(G143), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n196), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n448), .A2(KEYINPUT90), .A3(KEYINPUT14), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n457));
  INV_X1    g271(.A(new_n448), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT14), .B1(new_n449), .B2(G116), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n448), .A2(KEYINPUT14), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n453), .B(new_n455), .C1(new_n462), .C2(new_n213), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT13), .B1(new_n226), .B2(G128), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n222), .B2(G143), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n226), .A2(KEYINPUT13), .A3(G128), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT88), .B1(new_n467), .B2(G134), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n469), .B(new_n196), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n454), .A2(new_n196), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n213), .B1(new_n448), .B2(new_n450), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT87), .B1(new_n474), .B2(new_n451), .ZN(new_n475));
  INV_X1    g289(.A(new_n451), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n476), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n472), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n463), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n310), .A2(new_n481), .A3(G953), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  OAI221_X1 g298(.A(new_n472), .B1(new_n475), .B2(new_n478), .C1(new_n468), .C2(new_n470), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n485), .B2(new_n463), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n188), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n487), .A2(new_n489), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT86), .B(G475), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n430), .B1(new_n432), .B2(new_n438), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n388), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n495), .B2(G902), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n447), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n312), .A2(new_n385), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n420), .A2(new_n435), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n222), .A2(G119), .ZN(new_n502));
  INV_X1    g316(.A(G119), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT24), .B(G110), .Z(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n504), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G110), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n501), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n509), .B1(new_n506), .B2(new_n508), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n514), .A2(G110), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n420), .B(new_n407), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT22), .B(G137), .ZN(new_n520));
  INV_X1    g334(.A(G953), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(G221), .A3(G234), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n520), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n516), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n516), .B2(new_n519), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n500), .B(new_n188), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G234), .ZN(new_n528));
  OAI21_X1  g342(.A(G217), .B1(new_n528), .B2(G902), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT70), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n510), .A2(new_n515), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n519), .B1(new_n436), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n523), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n516), .A2(new_n519), .A3(new_n524), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n500), .B1(new_n536), .B2(new_n188), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n499), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n188), .B1(new_n525), .B2(new_n526), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT25), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(KEYINPUT73), .A3(new_n527), .A4(new_n530), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n529), .A2(new_n188), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n538), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT28), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n196), .A2(G137), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n194), .A2(G134), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n547), .A2(new_n548), .A3(G131), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n206), .B2(new_n190), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n286), .B2(new_n228), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n262), .A2(new_n263), .B1(new_n254), .B2(new_n255), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n333), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n256), .B1(new_n202), .B2(new_n207), .ZN(new_n554));
  INV_X1    g368(.A(new_n333), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n554), .B(new_n555), .C1(new_n244), .C2(new_n550), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n546), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n551), .A2(new_n552), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT28), .B1(new_n558), .B2(new_n555), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT68), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G101), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n393), .A2(G210), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n561), .B(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n557), .A2(new_n559), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(G902), .B1(new_n567), .B2(KEYINPUT29), .ZN(new_n568));
  INV_X1    g382(.A(new_n550), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n274), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n555), .B1(new_n570), .B2(new_n554), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n551), .A2(new_n333), .A3(new_n552), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT28), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n556), .A2(new_n546), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n565), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT30), .B1(new_n551), .B2(new_n552), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n554), .B(new_n577), .C1(new_n244), .C2(new_n550), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n555), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n566), .B1(new_n579), .B2(new_n572), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n577), .B1(new_n570), .B2(new_n554), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n551), .A2(KEYINPUT30), .A3(new_n552), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n333), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n556), .A2(new_n565), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(KEYINPUT31), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT31), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n579), .B2(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n573), .A2(new_n574), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n590), .A2(new_n592), .B1(new_n593), .B2(new_n566), .ZN(new_n594));
  NOR2_X1   g408(.A1(G472), .A2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n594), .A2(KEYINPUT32), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n566), .B1(new_n557), .B2(new_n559), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT31), .B1(new_n587), .B2(new_n589), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n579), .A2(new_n591), .A3(new_n588), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n598), .B1(new_n602), .B2(new_n595), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n584), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT69), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT32), .B1(new_n594), .B2(new_n596), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n602), .A2(new_n598), .A3(new_n595), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT69), .A3(new_n584), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n498), .A2(new_n545), .A3(new_n606), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n590), .A2(new_n592), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n596), .B1(new_n614), .B2(new_n599), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n594), .B2(G902), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n545), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n613), .B1(new_n618), .B2(new_n312), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n602), .B2(new_n188), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n538), .A2(new_n541), .A3(new_n544), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n621), .A2(new_n622), .A3(new_n615), .ZN(new_n623));
  INV_X1    g437(.A(new_n311), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n299), .B2(new_n308), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(KEYINPUT94), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n447), .A2(new_n496), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT33), .B1(new_n484), .B2(new_n486), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n480), .A2(new_n483), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n485), .A2(new_n482), .A3(new_n463), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(G902), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  MUX2_X1   g447(.A(new_n487), .B(new_n633), .S(G478), .Z(new_n634));
  NAND2_X1  g448(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n385), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n619), .A2(new_n626), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  NAND2_X1  g453(.A1(new_n367), .A2(new_n380), .ZN(new_n640));
  INV_X1    g454(.A(new_n381), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n382), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n326), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n447), .B(new_n496), .C1(new_n490), .C2(new_n491), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n325), .B(KEYINPUT95), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n619), .A3(new_n626), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR2_X1   g465(.A1(new_n524), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n533), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n543), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n538), .A2(new_n541), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n617), .A2(new_n616), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n498), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT96), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  AOI21_X1  g475(.A(new_n620), .B1(new_n568), .B2(new_n582), .ZN(new_n662));
  AOI211_X1 g476(.A(new_n605), .B(new_n662), .C1(new_n607), .C2(new_n608), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT69), .B1(new_n609), .B2(new_n584), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n655), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n312), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n323), .A2(G900), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT97), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n320), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n644), .A2(new_n645), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n665), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XNOR2_X1  g488(.A(new_n670), .B(KEYINPUT39), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n625), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT99), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n597), .A2(new_n603), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT98), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n587), .A2(new_n589), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(KEYINPUT98), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n620), .B1(new_n685), .B2(new_n188), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n326), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n492), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n690), .A2(new_n627), .A3(new_n666), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n643), .B(KEYINPUT38), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n678), .A2(new_n679), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT100), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NAND3_X1  g510(.A1(new_n627), .A2(new_n634), .A3(new_n670), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n644), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(KEYINPUT101), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n697), .B2(new_n644), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n665), .A2(new_n700), .A3(new_n667), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  AND3_X1   g518(.A1(new_n606), .A2(new_n545), .A3(new_n610), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n187), .A2(KEYINPUT102), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n293), .B(KEYINPUT12), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n708), .A2(new_n306), .B1(new_n278), .B2(new_n283), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n284), .A2(new_n297), .ZN(new_n711));
  INV_X1    g525(.A(new_n707), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n188), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n311), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n710), .A2(new_n713), .A3(KEYINPUT103), .A4(new_n311), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n705), .A2(new_n706), .A3(new_n636), .A4(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n606), .A3(new_n545), .A4(new_n610), .ZN(new_n720));
  INV_X1    g534(.A(new_n636), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT104), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  INV_X1    g539(.A(new_n720), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n648), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT105), .B(G116), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G18));
  AND3_X1   g543(.A1(new_n716), .A2(new_n655), .A3(new_n717), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n385), .A2(new_n497), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n606), .A3(new_n610), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NAND4_X1  g547(.A1(new_n623), .A2(new_n646), .A3(new_n716), .A4(new_n717), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n690), .A2(new_n627), .A3(new_n643), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT106), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n618), .A2(new_n647), .ZN(new_n737));
  INV_X1    g551(.A(new_n735), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n718), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NOR2_X1   g556(.A1(new_n697), .A2(new_n656), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n718), .A3(new_n699), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  XOR2_X1   g559(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n299), .A2(new_n747), .A3(new_n308), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n747), .B1(new_n299), .B2(new_n308), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n642), .A2(new_n311), .A3(new_n326), .A4(new_n382), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n545), .A3(new_n606), .A4(new_n610), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n746), .B1(new_n752), .B2(new_n697), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n622), .B1(new_n609), .B2(new_n584), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n751), .A2(KEYINPUT42), .A3(new_n698), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NOR2_X1   g571(.A1(new_n645), .A2(new_n671), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n665), .A2(new_n545), .A3(new_n751), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  NOR2_X1   g574(.A1(new_n643), .A2(new_n689), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n634), .A2(new_n496), .A3(new_n447), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT43), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n766), .B(new_n655), .C1(new_n615), .C2(new_n621), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n301), .B1(new_n304), .B2(new_n307), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n189), .B1(new_n771), .B2(G469), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .B1(new_n187), .B2(new_n298), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(KEYINPUT46), .B2(new_n772), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n311), .A3(new_n675), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n769), .B(new_n775), .C1(new_n768), .C2(new_n767), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n311), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT47), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n698), .A2(new_n622), .A3(new_n761), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n779), .A2(new_n665), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NOR2_X1   g596(.A1(G952), .A2(G953), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT118), .ZN(new_n784));
  INV_X1    g598(.A(new_n320), .ZN(new_n785));
  INV_X1    g599(.A(new_n718), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n762), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n766), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n754), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT48), .Z(new_n790));
  NAND3_X1  g604(.A1(new_n766), .A2(new_n785), .A3(new_n623), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n644), .A3(new_n786), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n787), .A2(new_n545), .A3(new_n785), .A4(new_n687), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n315), .B1(new_n793), .B2(new_n635), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n790), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n786), .A2(new_n326), .A3(new_n692), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT50), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT115), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n710), .A2(new_n713), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT110), .Z(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n779), .B1(new_n311), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n791), .A2(new_n762), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n798), .A2(KEYINPUT115), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n793), .A2(new_n627), .A3(new_n634), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n657), .B2(new_n788), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n799), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n803), .A2(new_n810), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n811), .A2(new_n804), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n798), .A2(KEYINPUT51), .A3(new_n808), .ZN(new_n814));
  OAI221_X1 g628(.A(new_n795), .B1(new_n809), .B2(KEYINPUT51), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT117), .Z(new_n816));
  NAND3_X1  g630(.A1(new_n703), .A2(new_n673), .A3(new_n744), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n687), .A2(new_n624), .A3(new_n655), .A4(new_n671), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n748), .A2(new_n749), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n818), .A2(new_n738), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  OR4_X1    g635(.A1(KEYINPUT113), .A2(new_n817), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n817), .B2(new_n820), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n673), .A2(new_n744), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n818), .A2(new_n738), .A3(new_n819), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n825), .A4(new_n703), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n826), .A3(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT111), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n606), .A2(new_n545), .A3(new_n610), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n831));
  INV_X1    g645(.A(new_n758), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n642), .A2(new_n326), .A3(new_n382), .A4(new_n670), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n497), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n667), .A2(new_n606), .A3(new_n610), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n743), .A2(new_n751), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n829), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n759), .A2(KEYINPUT111), .A3(new_n837), .A4(new_n836), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n756), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n646), .B(new_n326), .C1(new_n383), .C2(new_n384), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n635), .B2(new_n645), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n619), .A2(new_n626), .A3(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n611), .A2(new_n732), .A3(new_n844), .A4(new_n658), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n726), .A2(new_n648), .B1(new_n736), .B2(new_n740), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n723), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT112), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n839), .A2(new_n756), .A3(new_n840), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n723), .A2(new_n845), .A3(new_n846), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI211_X1 g666(.A(KEYINPUT53), .B(new_n828), .C1(new_n848), .C2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n823), .A2(new_n826), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n851), .B1(new_n849), .B2(new_n850), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n841), .A2(new_n847), .A3(KEYINPUT112), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n853), .B1(KEYINPUT53), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n854), .B1(new_n852), .B2(new_n848), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n864), .A2(KEYINPUT114), .A3(KEYINPUT53), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT53), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n863), .A2(new_n865), .B1(new_n828), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n860), .B1(KEYINPUT54), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n784), .B1(new_n816), .B2(new_n868), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n801), .B(KEYINPUT49), .Z(new_n870));
  NAND4_X1  g684(.A1(new_n687), .A2(new_n545), .A3(new_n311), .A4(new_n326), .ZN(new_n871));
  OR4_X1    g685(.A1(new_n692), .A2(new_n870), .A3(new_n763), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(G75));
  NAND2_X1  g687(.A1(new_n355), .A2(new_n366), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n364), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT55), .Z(new_n876));
  AOI21_X1  g690(.A(KEYINPUT119), .B1(new_n867), .B2(G902), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n828), .A2(new_n866), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT114), .B1(new_n864), .B2(KEYINPUT53), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n188), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  AOI211_X1 g698(.A(KEYINPUT56), .B(new_n876), .C1(new_n884), .C2(new_n641), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n881), .A2(new_n188), .A3(new_n381), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(new_n876), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n521), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(G51));
  XNOR2_X1  g704(.A(new_n867), .B(KEYINPUT54), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n189), .B(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n711), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n771), .A2(G469), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT120), .Z(new_n896));
  NAND2_X1  g710(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n889), .B1(new_n894), .B2(new_n897), .ZN(G54));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n899));
  INV_X1    g713(.A(new_n440), .ZN(new_n900));
  AND2_X1   g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n884), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n867), .A2(KEYINPUT119), .A3(G902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n882), .B1(new_n881), .B2(new_n188), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n889), .B1(new_n905), .B2(new_n440), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n903), .A2(new_n904), .A3(new_n900), .A4(new_n901), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT121), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n902), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n902), .A2(new_n906), .A3(new_n911), .A4(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(G60));
  AND2_X1   g727(.A1(new_n628), .A2(new_n632), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT59), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n891), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n868), .B2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n889), .ZN(G63));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(G217), .B2(G902), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n481), .A2(new_n188), .A3(KEYINPUT60), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n881), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n653), .ZN(new_n925));
  INV_X1    g739(.A(new_n889), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n925), .B(new_n926), .C1(new_n536), .C2(new_n924), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT61), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n927), .B(new_n929), .ZN(G66));
  OAI21_X1  g744(.A(G953), .B1(new_n321), .B2(new_n362), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT124), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n847), .B2(new_n521), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n874), .B1(G898), .B2(new_n521), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT125), .Z(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  NOR2_X1   g750(.A1(new_n585), .A2(new_n586), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n422), .A2(new_n423), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n937), .B(new_n938), .Z(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT126), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n695), .A2(new_n703), .A3(new_n824), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT62), .Z(new_n942));
  AND2_X1   g756(.A1(new_n635), .A2(new_n645), .ZN(new_n943));
  OR4_X1    g757(.A1(new_n830), .A2(new_n677), .A3(new_n762), .A4(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n781), .A2(new_n776), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n940), .B1(new_n946), .B2(new_n521), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n775), .A2(new_n738), .A3(new_n754), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT127), .Z(new_n949));
  NOR2_X1   g763(.A1(new_n817), .A2(new_n833), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n945), .A2(new_n756), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n951), .A2(G953), .ZN(new_n952));
  INV_X1    g766(.A(new_n939), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(G900), .B2(G953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n947), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(G900), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n281), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G72));
  NOR3_X1   g772(.A1(new_n579), .A2(new_n565), .A3(new_n572), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n951), .A2(new_n847), .ZN(new_n960));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT63), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n946), .A2(new_n847), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n565), .B1(new_n579), .B2(new_n572), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n963), .B(new_n926), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n962), .B1(new_n580), .B2(new_n683), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n859), .B2(new_n968), .ZN(G57));
endmodule


