//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204));
  NOR3_X1   g003(.A1(new_n204), .A2(G169gat), .A3(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(KEYINPUT65), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G183gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT66), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n204), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223));
  XNOR2_X1  g022(.A(G183gat), .B(G190gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n223), .B(new_n219), .C1(new_n224), .C2(new_n213), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n212), .A2(new_n221), .A3(new_n222), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT25), .ZN(new_n227));
  XOR2_X1   g026(.A(G113gat), .B(G120gat), .Z(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G127gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n231), .A2(KEYINPUT69), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(KEYINPUT69), .ZN(new_n233));
  OAI21_X1  g032(.A(G134gat), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G134gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n238));
  NAND2_X1  g037(.A1(G127gat), .A2(G134gat), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n236), .B2(new_n239), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n229), .B(new_n228), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n214), .B2(new_n216), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT26), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT27), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G183gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(G190gat), .B1(new_n249), .B2(KEYINPUT67), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n248), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT27), .B(G183gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(KEYINPUT28), .A3(new_n216), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n247), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n210), .A2(new_n261), .A3(new_n222), .A4(new_n206), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n219), .B1(new_n224), .B2(new_n213), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(KEYINPUT64), .ZN(new_n264));
  OR3_X1    g063(.A1(new_n218), .A2(KEYINPUT64), .A3(new_n220), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n227), .A2(new_n243), .A3(new_n260), .A4(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n255), .B1(KEYINPUT67), .B2(new_n257), .ZN(new_n270));
  INV_X1    g069(.A(new_n248), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n258), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n273), .A2(new_n247), .B1(new_n265), .B2(new_n264), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n274), .A2(KEYINPUT71), .A3(new_n243), .A4(new_n227), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n237), .A2(new_n242), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n266), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n218), .A2(new_n220), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(new_n223), .B1(new_n208), .B2(new_n211), .ZN(new_n279));
  INV_X1    g078(.A(new_n222), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n263), .B2(KEYINPUT66), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n261), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n276), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n269), .A2(new_n275), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  XNOR2_X1  g087(.A(G15gat), .B(G43gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G71gat), .B(G99gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n288), .B1(new_n292), .B2(KEYINPUT72), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(KEYINPUT72), .B2(new_n292), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT73), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n284), .B2(new_n286), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n294), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n291), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n287), .A2(new_n288), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n296), .A2(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n269), .A2(new_n285), .A3(new_n275), .A4(new_n283), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n305), .B(KEYINPUT34), .Z(new_n306));
  NOR3_X1   g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(new_n308), .A3(new_n292), .ZN(new_n309));
  AND4_X1   g108(.A1(new_n299), .A2(new_n287), .A3(KEYINPUT32), .A4(new_n294), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n299), .B1(new_n298), .B2(new_n294), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n306), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT77), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n309), .B(new_n306), .C1(new_n310), .C2(new_n311), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT76), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n202), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n312), .A2(KEYINPUT74), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n309), .B(new_n321), .C1(new_n310), .C2(new_n311), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n322), .A3(new_n313), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n202), .B1(new_n303), .B2(new_n306), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n319), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n319), .A3(new_n324), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n318), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT81), .B1(new_n329), .B2(G141gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(G148gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n330), .B(new_n333), .C1(new_n332), .C2(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335));
  INV_X1    g134(.A(G155gat), .ZN(new_n336));
  INV_X1    g135(.A(G162gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n336), .B2(new_n337), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n329), .A2(G141gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n332), .A2(G148gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G155gat), .B(G162gat), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351));
  AND2_X1   g150(.A1(G211gat), .A2(G218gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(KEYINPUT22), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(G211gat), .A2(G218gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n353), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n346), .A2(KEYINPUT84), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n345), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n347), .B1(new_n356), .B2(new_n349), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n358), .B(new_n359), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n357), .B2(KEYINPUT29), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n340), .A2(new_n345), .A3(KEYINPUT82), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT82), .B1(new_n340), .B2(new_n345), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n367), .A2(new_n371), .B1(new_n350), .B2(new_n357), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n365), .B1(new_n359), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G22gat), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n365), .B(new_n375), .C1(new_n359), .C2(new_n372), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378));
  INV_X1    g177(.A(G50gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT86), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n382), .B(KEYINPUT86), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n374), .A2(new_n376), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G226gat), .ZN(new_n388));
  INV_X1    g187(.A(G233gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n277), .A2(new_n282), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(KEYINPUT29), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(new_n274), .B2(new_n227), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n357), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n392), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n277), .B2(new_n282), .ZN(new_n396));
  INV_X1    g195(.A(new_n390), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n274), .A2(new_n397), .A3(new_n227), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n398), .A3(new_n356), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  NAND4_X1  g201(.A1(new_n394), .A2(KEYINPUT30), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n402), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n396), .A2(new_n398), .A3(new_n356), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n356), .B1(new_n396), .B2(new_n398), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n405), .A2(new_n406), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n410), .A2(KEYINPUT78), .A3(KEYINPUT30), .A4(new_n402), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT79), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n243), .A2(new_n360), .A3(new_n414), .A4(new_n362), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n276), .A2(new_n346), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n346), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n368), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n276), .B(new_n348), .C1(new_n420), .C2(new_n366), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n417), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n369), .A2(new_n370), .A3(new_n366), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n276), .B1(new_n346), .B2(new_n347), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n243), .A2(new_n360), .A3(KEYINPUT4), .A4(new_n362), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(KEYINPUT4), .B2(new_n416), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n416), .B1(new_n371), .B2(new_n276), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT5), .B1(new_n431), .B2(new_n423), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n424), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT0), .ZN(new_n435));
  XNOR2_X1  g234(.A(G57gat), .B(G85gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n435), .B(new_n436), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n424), .B(new_n437), .C1(new_n430), .C2(new_n432), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(KEYINPUT6), .A3(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n394), .A2(new_n399), .A3(new_n402), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n394), .A2(KEYINPUT80), .A3(new_n399), .A4(new_n402), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n387), .B1(new_n413), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n447), .A2(new_n449), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n399), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT90), .A4(new_n356), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n394), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT37), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n404), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n410), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n453), .A2(new_n463), .A3(new_n442), .A4(new_n443), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT37), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT37), .B1(new_n405), .B2(new_n406), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n404), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n467), .B2(KEYINPUT91), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n469), .A3(new_n404), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n459), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n387), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n431), .A2(new_n423), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT39), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n423), .B1(new_n417), .B2(new_n421), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n438), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(KEYINPUT40), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n439), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT40), .B1(new_n477), .B2(new_n479), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n412), .A2(new_n485), .A3(new_n450), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n412), .B2(new_n450), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n484), .B(KEYINPUT89), .C1(new_n486), .C2(new_n487), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n452), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n323), .A2(new_n387), .A3(new_n316), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n413), .A2(new_n451), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT35), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT76), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n316), .B(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n384), .A2(new_n386), .ZN(new_n497));
  INV_X1    g296(.A(new_n444), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT35), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n304), .B1(new_n303), .B2(new_n306), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n312), .A2(KEYINPUT77), .A3(new_n313), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n496), .A2(new_n499), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n328), .A2(new_n491), .B1(new_n494), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(G1gat), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n506), .B1(new_n509), .B2(KEYINPUT93), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(G1gat), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI221_X1 g311(.A(new_n509), .B1(KEYINPUT93), .B2(new_n506), .C1(G1gat), .C2(new_n507), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G29gat), .ZN(new_n515));
  INV_X1    g314(.A(G36gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT15), .A4(new_n520), .ZN(new_n524));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n514), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n527), .B(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(new_n514), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT18), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n527), .B(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n533), .B(new_n528), .C1(new_n536), .C2(new_n514), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n514), .B(new_n527), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n533), .B(KEYINPUT13), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n534), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n539), .A3(new_n542), .A4(new_n549), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n543), .A2(KEYINPUT94), .A3(new_n550), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n505), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n336), .ZN(new_n559));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G57gat), .B(G64gat), .Z(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OR3_X1    g366(.A1(KEYINPUT95), .A2(G71gat), .A3(G78gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n567), .A2(new_n564), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G71gat), .ZN(new_n571));
  INV_X1    g370(.A(G78gat), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n571), .B(new_n572), .C1(KEYINPUT96), .C2(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n564), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n566), .A2(KEYINPUT96), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n563), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G127gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n577), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n514), .B1(KEYINPUT21), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n582), .A2(new_n585), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n562), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n586), .A3(new_n561), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595));
  XOR2_X1   g394(.A(G99gat), .B(G106gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT97), .B(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n598), .A2(new_n599), .B1(KEYINPUT8), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT7), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n597), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n577), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n603), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n596), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n601), .A2(KEYINPUT98), .A3(new_n597), .A4(new_n603), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n596), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT99), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n604), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n613), .A2(new_n615), .B1(new_n608), .B2(new_n609), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n595), .B(new_n611), .C1(new_n616), .C2(new_n583), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n605), .A2(new_n610), .A3(KEYINPUT101), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT10), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n583), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n594), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(new_n610), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n604), .B(KEYINPUT99), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n577), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT101), .B1(new_n605), .B2(new_n610), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n594), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n630), .ZN(new_n638));
  INV_X1    g437(.A(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(G232gat), .A2(G233gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT41), .ZN(new_n643));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n530), .B1(new_n624), .B2(new_n625), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(KEYINPUT100), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n648), .A2(KEYINPUT100), .B1(KEYINPUT41), .B2(new_n642), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n616), .B2(new_n527), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n647), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n650), .B1(new_n647), .B2(new_n653), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n646), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n645), .A3(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n593), .A2(new_n641), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n557), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n498), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n663), .A2(new_n503), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G8gat), .B1(new_n663), .B2(new_n503), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(KEYINPUT104), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n669), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n670), .A2(new_n671), .B1(new_n668), .B2(new_n675), .ZN(G1325gat));
  NOR2_X1   g475(.A1(new_n315), .A2(new_n317), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n663), .A2(G15gat), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n663), .B2(new_n328), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n663), .A2(new_n387), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  OAI21_X1  g483(.A(KEYINPUT44), .B1(new_n505), .B2(new_n660), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n494), .A2(new_n504), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT36), .B1(new_n496), .B2(new_n502), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n323), .A2(new_n319), .A3(new_n324), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(new_n325), .ZN(new_n689));
  INV_X1    g488(.A(new_n452), .ZN(new_n690));
  AND4_X1   g489(.A1(new_n443), .A2(new_n453), .A3(new_n463), .A4(new_n442), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n468), .A2(new_n470), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT38), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n497), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n483), .A2(new_n482), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n480), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n412), .A2(new_n450), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n412), .A2(new_n485), .A3(new_n450), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n694), .B1(new_n700), .B2(KEYINPUT89), .ZN(new_n701));
  INV_X1    g500(.A(new_n490), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n690), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n686), .B1(new_n689), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n661), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n641), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n593), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n556), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n498), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n515), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n712), .B2(new_n711), .ZN(new_n714));
  NOR4_X1   g513(.A1(new_n505), .A2(new_n556), .A3(new_n660), .A4(new_n709), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n515), .A3(new_n498), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT106), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(new_n719), .ZN(G1328gat));
  INV_X1    g519(.A(new_n503), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n715), .A2(new_n516), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT46), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n710), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n724), .B2(new_n503), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1329gat));
  AND2_X1   g525(.A1(new_n715), .A2(new_n677), .ZN(new_n727));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n328), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n727), .A2(G43gat), .B1(new_n724), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT47), .ZN(G1330gat));
  AND2_X1   g531(.A1(new_n715), .A2(new_n497), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n387), .A2(new_n379), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n733), .A2(G50gat), .B1(new_n724), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g536(.A1(new_n592), .A2(new_n556), .A3(new_n660), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n704), .A2(new_n641), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n498), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n721), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  AOI21_X1  g544(.A(new_n571), .B1(new_n739), .B2(new_n689), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n678), .A2(G71gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n739), .A2(new_n497), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(G78gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1335gat));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n704), .A2(new_n661), .ZN(new_n754));
  INV_X1    g553(.A(new_n556), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n592), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n661), .A4(new_n756), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(new_n498), .A3(new_n598), .A4(new_n641), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n757), .A2(new_n708), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n707), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n444), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n764), .B2(new_n598), .ZN(G1336gat));
  NAND3_X1  g564(.A1(new_n758), .A2(KEYINPUT110), .A3(new_n759), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n767), .B(new_n753), .C1(new_n754), .C2(new_n757), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n503), .A2(new_n708), .A3(G92gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G92gat), .B1(new_n763), .B2(new_n503), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n760), .A2(new_n769), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(G1337gat));
  XOR2_X1   g576(.A(KEYINPUT112), .B(G99gat), .Z(new_n778));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n677), .A3(new_n641), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n328), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n778), .ZN(G1338gat));
  INV_X1    g580(.A(new_n762), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n387), .B(new_n782), .C1(new_n685), .C2(new_n706), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT113), .B(G106gat), .Z(new_n784));
  OAI21_X1  g583(.A(KEYINPUT114), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n707), .A2(new_n497), .A3(new_n762), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787));
  INV_X1    g586(.A(new_n784), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n387), .A2(G106gat), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n641), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n766), .A2(new_n768), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n785), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT53), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT53), .B1(new_n786), .B2(new_n788), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n760), .A2(new_n641), .A3(new_n790), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(G1339gat));
  OAI211_X1 g597(.A(new_n629), .B(new_n620), .C1(new_n628), .C2(KEYINPUT10), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n622), .A2(new_n799), .A3(KEYINPUT54), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n801), .B(new_n594), .C1(new_n619), .C2(new_n621), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n639), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n637), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n802), .A2(new_n639), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT55), .B1(new_n805), .B2(new_n800), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n532), .A2(new_n533), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n540), .A2(new_n541), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n548), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n657), .A2(new_n659), .A3(new_n553), .A4(new_n809), .ZN(new_n810));
  NOR4_X1   g609(.A1(new_n804), .A2(new_n806), .A3(KEYINPUT116), .A4(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n803), .A2(new_n637), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n800), .A2(new_n639), .A3(new_n802), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n810), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n812), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n553), .A2(new_n809), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n641), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n637), .A3(new_n554), .A4(new_n555), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n806), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n660), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n592), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n738), .A2(KEYINPUT115), .A3(new_n708), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT115), .B1(new_n738), .B2(new_n708), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n828), .A2(new_n444), .A3(new_n492), .A4(new_n721), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n755), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n503), .A2(new_n498), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n824), .A2(new_n827), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT117), .A3(new_n387), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n828), .B2(new_n497), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n678), .B(new_n831), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n755), .A2(G113gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n830), .B1(new_n836), .B2(new_n837), .ZN(G1340gat));
  AOI21_X1  g637(.A(G120gat), .B1(new_n829), .B2(new_n641), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n641), .A2(G120gat), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n836), .B2(new_n840), .ZN(G1341gat));
  NAND2_X1  g640(.A1(new_n836), .A2(new_n592), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n232), .A2(new_n233), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n593), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(G1342gat));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n235), .A3(new_n661), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT56), .Z(new_n849));
  AND2_X1   g648(.A1(new_n836), .A2(new_n661), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n235), .ZN(G1343gat));
  NOR3_X1   g650(.A1(new_n689), .A2(new_n387), .A3(new_n721), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n832), .A2(new_n498), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n332), .B1(new_n853), .B2(new_n556), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n622), .A2(new_n799), .A3(KEYINPUT54), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n802), .A2(new_n639), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n814), .A2(KEYINPUT119), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n820), .B1(new_n863), .B2(new_n821), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n660), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n818), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n827), .B1(new_n866), .B2(new_n593), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT57), .B1(new_n867), .B2(new_n387), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n689), .A2(new_n831), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n497), .B1(new_n824), .B2(new_n827), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n868), .B(new_n869), .C1(KEYINPUT57), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n755), .A2(G141gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n854), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g673(.A(new_n853), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n329), .A3(new_n641), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n871), .A2(new_n708), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .A3(new_n329), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n738), .A2(KEYINPUT120), .A3(new_n708), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n738), .B2(new_n708), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n804), .A2(new_n806), .A3(new_n810), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n864), .B2(new_n660), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n592), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n387), .A2(KEYINPUT57), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n870), .A2(KEYINPUT57), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n641), .A3(new_n869), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n879), .B1(new_n888), .B2(G148gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n876), .B1(new_n878), .B2(new_n889), .ZN(G1345gat));
  OAI21_X1  g689(.A(G155gat), .B1(new_n871), .B2(new_n593), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n336), .A3(new_n592), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n871), .B2(new_n660), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n337), .A3(new_n661), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n721), .A2(new_n444), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n828), .A2(new_n492), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n755), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n678), .B(new_n897), .C1(new_n833), .C2(new_n835), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n755), .A2(G169gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(G1348gat));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903));
  INV_X1    g702(.A(new_n898), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G176gat), .A3(new_n708), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n900), .A2(new_n641), .ZN(new_n907));
  INV_X1    g706(.A(G176gat), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n903), .B(new_n906), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n900), .B2(new_n641), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT121), .B1(new_n910), .B2(new_n905), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1349gat));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n904), .A2(new_n252), .A3(new_n593), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n900), .A2(new_n592), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n913), .B(new_n915), .C1(new_n916), .C2(new_n214), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n214), .B1(new_n900), .B2(new_n592), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT60), .B1(new_n918), .B2(new_n914), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1350gat));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n661), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G190gat), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n898), .A2(new_n216), .A3(new_n661), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT122), .Z(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(G1351gat));
  INV_X1    g727(.A(new_n870), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n689), .A2(new_n897), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n755), .ZN(new_n933));
  OR3_X1    g732(.A1(new_n689), .A2(KEYINPUT123), .A3(new_n897), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n689), .B2(new_n897), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n887), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n755), .A2(G197gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  NOR3_X1   g739(.A1(new_n931), .A2(G204gat), .A3(new_n708), .ZN(new_n941));
  XNOR2_X1  g740(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(G204gat), .B1(new_n937), .B2(new_n708), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1353gat));
  INV_X1    g744(.A(G211gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n932), .A2(new_n946), .A3(new_n592), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n887), .A2(new_n592), .A3(new_n936), .ZN(new_n948));
  AND2_X1   g747(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n949));
  OAI21_X1  g748(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n949), .B1(new_n948), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n956), .B(new_n947), .C1(new_n952), .C2(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1354gat));
  AND3_X1   g757(.A1(new_n938), .A2(G218gat), .A3(new_n661), .ZN(new_n959));
  AOI21_X1  g758(.A(G218gat), .B1(new_n932), .B2(new_n661), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1355gat));
endmodule


