//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n459), .A2(G137), .A3(new_n458), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT66), .ZN(G160));
  NAND2_X1  g046(.A1(new_n459), .A2(new_n458), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n458), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n474), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n475), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n485), .B(new_n489), .C1(new_n475), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n458), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n478), .B2(G126), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(G75), .A2(G543), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n503), .A2(G651), .B1(new_n508), .B2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT67), .B1(new_n506), .B2(new_n501), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n507), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n509), .B1(new_n510), .B2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n508), .A2(G51), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT68), .B(KEYINPUT7), .Z(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n519), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT69), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT69), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n524), .B1(new_n530), .B2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n501), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G651), .B1(new_n508), .B2(G52), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n511), .A2(G90), .A3(new_n518), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n501), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(new_n508), .B2(G43), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n511), .A2(G81), .A3(new_n518), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT70), .Z(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND3_X1  g126(.A1(new_n511), .A2(G91), .A3(new_n518), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT72), .B(G65), .Z(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(new_n501), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n508), .A2(new_n558), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n516), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n559), .B2(new_n562), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n557), .B1(new_n565), .B2(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n530), .A2(new_n531), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(new_n523), .ZN(G286));
  INV_X1    g144(.A(G651), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n570), .B1(new_n501), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(G49), .B2(new_n508), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n511), .A2(G87), .A3(new_n518), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n511), .A2(G86), .A3(new_n518), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n508), .A2(G48), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n513), .B2(new_n514), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n581), .B2(KEYINPUT73), .ZN(new_n582));
  OAI211_X1 g157(.A(KEYINPUT73), .B(G61), .C1(new_n499), .C2(new_n500), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n578), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n508), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  XOR2_X1   g163(.A(KEYINPUT74), .B(G85), .Z(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n570), .B2(new_n588), .C1(new_n519), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n511), .A2(G92), .A3(new_n518), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n501), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n508), .B2(G54), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n603), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G168), .B2(new_n603), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n543), .A2(new_n544), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n603), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n599), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n473), .A2(G135), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G111), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G2105), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n478), .B2(G123), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n459), .A2(new_n466), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n622), .A2(G2096), .B1(G2100), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(G2100), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n627), .B(new_n628), .C1(G2096), .C2(new_n622), .ZN(G156));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT77), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n647), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n654), .A2(new_n649), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n655), .B1(new_n648), .B2(new_n649), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n654), .B2(new_n649), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n652), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2096), .B(G2100), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT79), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  OR2_X1    g245(.A1(new_n663), .A2(new_n665), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n668), .A3(new_n666), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n670), .B(new_n672), .C1(new_n668), .C2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n676), .ZN(new_n680));
  INV_X1    g255(.A(new_n678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G23), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n573), .A2(new_n574), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT83), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT33), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT84), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(G6), .A2(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G305), .B2(new_n684), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT32), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT82), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n684), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n684), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G1971), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n695), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(G1971), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n696), .A2(new_n699), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n691), .A2(KEYINPUT34), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(KEYINPUT34), .B1(new_n691), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n478), .A2(G119), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT80), .Z(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(G107), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G2105), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n473), .B2(G131), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n706), .B1(new_n714), .B2(new_n705), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XOR2_X1   g291(.A(new_n715), .B(new_n716), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n684), .A2(G24), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT81), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G290), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1986), .Z(new_n721));
  NOR2_X1   g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n703), .A2(new_n704), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT36), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(KEYINPUT36), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(G160), .A2(G29), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n728), .B2(KEYINPUT24), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT24), .B2(new_n728), .ZN(new_n730));
  AOI21_X1  g305(.A(G2084), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n705), .A2(G33), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n459), .A2(G127), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n458), .B1(new_n735), .B2(KEYINPUT89), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(KEYINPUT89), .B2(new_n735), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT25), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n473), .A2(KEYINPUT88), .A3(G139), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n741));
  INV_X1    g316(.A(G139), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n472), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n732), .B1(new_n745), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n731), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n727), .A2(G2084), .A3(new_n730), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n545), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G16), .B2(G19), .ZN(new_n754));
  INV_X1    g329(.A(G1341), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NOR2_X1   g332(.A1(G5), .A2(G16), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT91), .Z(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G301), .B2(new_n684), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n756), .A2(new_n757), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n705), .A2(G32), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n459), .A2(G2105), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n466), .A2(G105), .ZN(new_n771));
  INV_X1    g346(.A(G141), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n472), .B2(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n765), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT92), .B(G2078), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n705), .A2(G27), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n705), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G11), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(G11), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(G28), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n705), .B1(new_n786), .B2(G28), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n784), .B(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n621), .B2(G29), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n705), .A2(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n705), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT29), .B(G2090), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n775), .A2(new_n776), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n790), .B(new_n794), .C1(new_n792), .C2(new_n793), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n752), .A2(new_n764), .A3(new_n782), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n684), .A2(G20), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT23), .ZN(new_n798));
  INV_X1    g373(.A(G299), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n684), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1956), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n684), .A2(G21), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G168), .B2(new_n684), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT90), .B(G1966), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n600), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G4), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT85), .B(G1348), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n705), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT28), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n478), .A2(G128), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n458), .A2(G116), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n813), .B1(new_n814), .B2(new_n815), .C1(new_n816), .C2(new_n472), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT86), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT87), .B(G2067), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n809), .A2(new_n810), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n796), .A2(new_n801), .A3(new_n805), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT93), .B1(new_n726), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n826), .B(new_n823), .C1(new_n724), .C2(new_n725), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n726), .A2(new_n824), .ZN(G150));
  NAND2_X1  g404(.A1(new_n600), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  INV_X1    g407(.A(G80), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n501), .A2(new_n832), .B1(new_n833), .B2(new_n507), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI221_X1 g411(.A(KEYINPUT94), .B1(new_n833), .B2(new_n507), .C1(new_n501), .C2(new_n832), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(G651), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n508), .A2(G55), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n511), .A2(G93), .A3(new_n518), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n609), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n840), .A2(new_n839), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n545), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n831), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT95), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n841), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  XNOR2_X1  g429(.A(KEYINPUT100), .B(G37), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n818), .ZN(new_n857));
  INV_X1    g432(.A(G126), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n768), .A2(new_n858), .B1(new_n492), .B2(new_n493), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  INV_X1    g435(.A(new_n490), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n489), .B1(new_n459), .B2(new_n485), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n488), .A2(KEYINPUT97), .A3(new_n490), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n488), .A2(KEYINPUT97), .A3(new_n490), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT97), .B1(new_n488), .B2(new_n490), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n495), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n818), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n866), .A2(new_n774), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n774), .B1(new_n866), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n745), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n818), .B(new_n869), .ZN(new_n874));
  INV_X1    g449(.A(new_n774), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n745), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n866), .A2(new_n774), .A3(new_n870), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n713), .B(new_n624), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n473), .A2(G142), .B1(G130), .B2(new_n478), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G118), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n883), .A2(KEYINPUT98), .B1(new_n884), .B2(G2105), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(KEYINPUT98), .B2(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n881), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT99), .B1(new_n880), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n891));
  AOI211_X1 g466(.A(new_n891), .B(new_n888), .C1(new_n873), .C2(new_n879), .ZN(new_n892));
  OAI22_X1  g467(.A1(new_n890), .A2(new_n892), .B1(new_n880), .B2(new_n889), .ZN(new_n893));
  XNOR2_X1  g468(.A(G160), .B(new_n482), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n622), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n856), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n889), .B1(new_n880), .B2(KEYINPUT101), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(KEYINPUT101), .B2(new_n880), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n871), .A2(new_n872), .A3(new_n745), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n889), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n891), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n880), .A2(KEYINPUT99), .A3(new_n889), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n905), .A3(new_n895), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT40), .B1(new_n897), .B2(new_n906), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(G395));
  NOR2_X1   g484(.A1(new_n841), .A2(G868), .ZN(new_n910));
  XNOR2_X1  g485(.A(G305), .B(G290), .ZN(new_n911));
  XNOR2_X1  g486(.A(G303), .B(G288), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n914));
  XOR2_X1   g489(.A(new_n913), .B(new_n914), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n611), .B(new_n845), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n599), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n559), .A2(new_n562), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT71), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n564), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n594), .A2(new_n920), .A3(new_n557), .A4(new_n598), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT41), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n921), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n594), .A2(new_n598), .B1(new_n920), .B2(new_n557), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n915), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n930), .B(new_n931), .Z(new_n932));
  AOI21_X1  g507(.A(new_n910), .B1(new_n932), .B2(G868), .ZN(G295));
  AOI21_X1  g508(.A(new_n910), .B1(new_n932), .B2(G868), .ZN(G331));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n842), .A2(new_n844), .A3(G301), .ZN(new_n936));
  AOI21_X1  g511(.A(G301), .B1(new_n842), .B2(new_n844), .ZN(new_n937));
  OAI21_X1  g512(.A(G286), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n845), .A2(G171), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n842), .A2(new_n844), .A3(G301), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(G168), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n925), .B2(new_n926), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n938), .A2(new_n941), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT104), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n923), .A2(new_n922), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n941), .A4(new_n938), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n938), .A2(new_n941), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n927), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n946), .A2(new_n949), .A3(new_n913), .A4(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n945), .A2(KEYINPUT104), .B1(new_n950), .B2(new_n927), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(KEYINPUT105), .A3(new_n913), .A4(new_n949), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n951), .A2(KEYINPUT106), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n913), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n951), .A2(KEYINPUT106), .A3(new_n945), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n856), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n957), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n913), .B1(new_n955), .B2(new_n949), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(G37), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n958), .B1(new_n957), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n935), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n957), .A2(new_n965), .A3(new_n958), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n958), .B1(new_n957), .B2(new_n962), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT44), .B(new_n968), .C1(new_n969), .C2(KEYINPUT107), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n969), .A2(KEYINPUT107), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G397));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT108), .B(G1384), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n869), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G40), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n462), .A2(new_n468), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n973), .B1(new_n978), .B2(G1996), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  INV_X1    g555(.A(new_n974), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n865), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n463), .A2(new_n469), .A3(G40), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT109), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n774), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT110), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n818), .B(G2067), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n875), .A2(new_n985), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n713), .B(new_n716), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT111), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n988), .B(new_n991), .C1(new_n978), .C2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(G290), .B(G1986), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n984), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT112), .B1(new_n865), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(new_n998), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n869), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1384), .B1(new_n491), .B2(new_n495), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n977), .B1(new_n1004), .B2(KEYINPUT45), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT113), .ZN(new_n1008));
  INV_X1    g583(.A(G1971), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1010), .A3(new_n1006), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT50), .B1(new_n869), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n977), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(G2090), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n997), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT55), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT114), .B(G8), .Z(new_n1024));
  NOR2_X1   g599(.A1(new_n865), .A2(G1384), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n977), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n686), .A2(G1976), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n869), .A2(new_n1013), .A3(new_n977), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1024), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n1028), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1031), .A2(new_n1035), .B1(new_n1036), .B2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n578), .A2(KEYINPUT116), .A3(new_n1038), .A4(new_n585), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n585), .A2(new_n1038), .A3(new_n576), .A4(new_n577), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1039), .A2(new_n1042), .B1(G1981), .B2(G305), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT49), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1049), .A3(new_n1026), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1037), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1023), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1026), .B1(new_n1048), .B2(KEYINPUT49), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1044), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n686), .A2(new_n1029), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1043), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1052), .B1(new_n1026), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n1059));
  INV_X1    g634(.A(G2078), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1010), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1061));
  AOI211_X1 g636(.A(KEYINPUT113), .B(new_n1005), .C1(new_n999), .C2(new_n1002), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n983), .B1(KEYINPUT45), .B2(new_n1004), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1025), .B2(KEYINPUT45), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1060), .A2(KEYINPUT53), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n761), .B2(new_n1017), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1059), .B1(new_n1072), .B2(G301), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1064), .B1(new_n1075), .B2(new_n1060), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n865), .B2(G1384), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n983), .B1(new_n1078), .B2(new_n1015), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT123), .B1(new_n1079), .B2(G1961), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1017), .A2(new_n1081), .A3(new_n761), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1069), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n983), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n982), .B2(new_n977), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1003), .B(new_n1084), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1074), .B1(new_n1076), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1066), .A2(KEYINPUT125), .A3(new_n1088), .A4(new_n1083), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(G171), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1073), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n983), .B1(new_n1077), .B2(new_n1004), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1025), .B2(new_n1077), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT120), .B(G1956), .Z(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT56), .B(G2072), .Z(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1003), .A2(new_n1006), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n559), .B2(new_n562), .ZN(new_n1102));
  AOI22_X1  g677(.A1(G299), .A2(KEYINPUT57), .B1(new_n557), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1079), .A2(G1348), .B1(G2067), .B2(new_n1032), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1105), .A2(new_n600), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1094), .B(new_n1104), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1107), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1104), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(new_n1107), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1117));
  OAI221_X1 g692(.A(KEYINPUT60), .B1(G2067), .B2(new_n1032), .C1(new_n1079), .C2(G1348), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n600), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1112), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1007), .A2(G1996), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1025), .B2(new_n977), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n545), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1118), .A2(new_n600), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT59), .B(new_n545), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1108), .B(new_n1110), .C1(new_n1120), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1093), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT117), .B1(new_n1135), .B2(new_n1055), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1037), .A2(new_n1050), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1096), .A2(G2090), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n1009), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1021), .B1(new_n1142), .B2(new_n1024), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1139), .A2(new_n1023), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G168), .A2(new_n1024), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(KEYINPUT51), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT45), .B1(new_n869), .B2(new_n1013), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1004), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n977), .B1(new_n1149), .B2(new_n980), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n804), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1068), .A2(KEYINPUT118), .A3(new_n804), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n983), .A2(G2084), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT119), .B(new_n1156), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1147), .B1(new_n1162), .B2(new_n1033), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(G8), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1145), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(G168), .B(new_n1024), .C1(new_n1155), .C2(new_n1161), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1163), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1076), .A2(new_n1089), .A3(G171), .ZN(new_n1171));
  AOI21_X1  g746(.A(G301), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1059), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1144), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1058), .B1(new_n1131), .B2(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(G286), .B(new_n1024), .C1(new_n1155), .C2(new_n1161), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1139), .A2(new_n1143), .A3(new_n1023), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1051), .A2(new_n1178), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1180), .A2(new_n1023), .A3(new_n1176), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1162), .A2(new_n1033), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1146), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n997), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT51), .B1(new_n1186), .B2(new_n1145), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1185), .B1(new_n1187), .B2(new_n1168), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AND4_X1   g765(.A1(new_n1139), .A2(new_n1143), .A3(new_n1023), .A4(new_n1172), .ZN(new_n1191));
  OAI211_X1 g766(.A(KEYINPUT62), .B(new_n1185), .C1(new_n1187), .C2(new_n1168), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1183), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n996), .B1(new_n1175), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n979), .A2(new_n986), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT46), .Z(new_n1197));
  INV_X1    g772(.A(KEYINPUT47), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n984), .B1(new_n989), .B2(new_n774), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1198), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  OAI22_X1  g779(.A1(new_n1201), .A2(new_n1202), .B1(new_n994), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n714), .A2(new_n716), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT126), .Z(new_n1207));
  NAND3_X1  g782(.A1(new_n988), .A2(new_n991), .A3(new_n1207), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n818), .A2(G2067), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n978), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT127), .B1(new_n1205), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1210), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n994), .A2(new_n1204), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1202), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n1200), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1211), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1195), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g794(.A(new_n456), .ZN(new_n1221));
  OR3_X1    g795(.A1(G401), .A2(new_n1221), .A3(G227), .ZN(new_n1222));
  AOI21_X1  g796(.A(new_n1222), .B1(new_n679), .B2(new_n682), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n880), .A2(new_n889), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1224), .B1(new_n903), .B2(new_n904), .ZN(new_n1225));
  OAI21_X1  g799(.A(new_n855), .B1(new_n1225), .B2(new_n895), .ZN(new_n1226));
  AND3_X1   g800(.A1(new_n899), .A2(new_n905), .A3(new_n895), .ZN(new_n1227));
  OAI21_X1  g801(.A(new_n1223), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g802(.A1(new_n963), .A2(new_n966), .ZN(new_n1229));
  NOR2_X1   g803(.A1(new_n1228), .A2(new_n1229), .ZN(G308));
  OAI221_X1 g804(.A(new_n1223), .B1(new_n1226), .B2(new_n1227), .C1(new_n963), .C2(new_n966), .ZN(G225));
endmodule


