

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U325 ( .A(n323), .B(n322), .ZN(n327) );
  XNOR2_X1 U326 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n412) );
  XNOR2_X1 U328 ( .A(n413), .B(n412), .ZN(n434) );
  XNOR2_X1 U329 ( .A(KEYINPUT109), .B(KEYINPUT48), .ZN(n397) );
  XNOR2_X1 U330 ( .A(n398), .B(n397), .ZN(n529) );
  NOR2_X1 U331 ( .A1(n451), .A2(n521), .ZN(n571) );
  XOR2_X1 U332 ( .A(n329), .B(n328), .Z(n558) );
  XNOR2_X1 U333 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(G211GAT), .B(KEYINPUT84), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n293), .B(KEYINPUT21), .ZN(n294) );
  XOR2_X1 U337 ( .A(n294), .B(KEYINPUT85), .Z(n296) );
  XNOR2_X1 U338 ( .A(G197GAT), .B(G218GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n399) );
  XNOR2_X1 U340 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n297), .B(KEYINPUT2), .ZN(n426) );
  XOR2_X1 U342 ( .A(G50GAT), .B(G162GAT), .Z(n317) );
  XOR2_X1 U343 ( .A(n426), .B(n317), .Z(n299) );
  NAND2_X1 U344 ( .A1(G228GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n399), .B(n300), .ZN(n312) );
  XOR2_X1 U347 ( .A(KEYINPUT87), .B(KEYINPUT82), .Z(n302) );
  XNOR2_X1 U348 ( .A(KEYINPUT24), .B(KEYINPUT83), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U350 ( .A(n303), .B(G204GAT), .Z(n305) );
  XOR2_X1 U351 ( .A(G22GAT), .B(G155GAT), .Z(n372) );
  XNOR2_X1 U352 ( .A(n372), .B(KEYINPUT86), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U354 ( .A(n306), .B(KEYINPUT23), .Z(n310) );
  XOR2_X1 U355 ( .A(G78GAT), .B(G148GAT), .Z(n308) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n356) );
  XNOR2_X1 U358 ( .A(n356), .B(KEYINPUT22), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n463) );
  XOR2_X1 U361 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n314) );
  XNOR2_X1 U362 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n329) );
  XOR2_X1 U364 ( .A(G29GAT), .B(G43GAT), .Z(n316) );
  XNOR2_X1 U365 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n336) );
  XOR2_X1 U367 ( .A(n317), .B(n336), .Z(n323) );
  XOR2_X1 U368 ( .A(KEYINPUT66), .B(G92GAT), .Z(n319) );
  XNOR2_X1 U369 ( .A(G134GAT), .B(G106GAT), .ZN(n318) );
  XOR2_X1 U370 ( .A(n319), .B(n318), .Z(n321) );
  NAND2_X1 U371 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n324), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U374 ( .A(G36GAT), .B(G190GAT), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n325), .B(KEYINPUT75), .ZN(n403) );
  XNOR2_X1 U376 ( .A(n355), .B(n403), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U378 ( .A(G141GAT), .B(G22GAT), .Z(n331) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(G197GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U381 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n333) );
  XNOR2_X1 U382 ( .A(G113GAT), .B(G8GAT), .ZN(n332) );
  XNOR2_X1 U383 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n343) );
  XOR2_X1 U385 ( .A(n336), .B(KEYINPUT29), .Z(n338) );
  NAND2_X1 U386 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G1GAT), .Z(n379) );
  XOR2_X1 U389 ( .A(n339), .B(n379), .Z(n341) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(G50GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n563) );
  XOR2_X1 U393 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n345) );
  XNOR2_X1 U394 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n360) );
  XNOR2_X1 U396 ( .A(G64GAT), .B(G92GAT), .ZN(n347) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(G204GAT), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n349) );
  INV_X1 U399 ( .A(n349), .ZN(n408) );
  NAND2_X1 U400 ( .A1(n408), .A2(KEYINPUT31), .ZN(n351) );
  INV_X1 U401 ( .A(KEYINPUT31), .ZN(n348) );
  NAND2_X1 U402 ( .A1(n349), .A2(n348), .ZN(n350) );
  NAND2_X1 U403 ( .A1(n351), .A2(n350), .ZN(n353) );
  AND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U406 ( .A(n355), .B(n354), .Z(n358) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U408 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U409 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U410 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n362) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G57GAT), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U413 ( .A(KEYINPUT13), .B(n363), .ZN(n371) );
  XNOR2_X1 U414 ( .A(n364), .B(n371), .ZN(n388) );
  XNOR2_X1 U415 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n388), .B(n365), .ZN(n501) );
  NAND2_X1 U417 ( .A1(n563), .A2(n501), .ZN(n367) );
  INV_X1 U418 ( .A(KEYINPUT46), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n384) );
  XOR2_X1 U420 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n369) );
  XNOR2_X1 U421 ( .A(G127GAT), .B(KEYINPUT12), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U423 ( .A(n371), .B(n370), .Z(n383) );
  XOR2_X1 U424 ( .A(G8GAT), .B(G183GAT), .Z(n400) );
  XOR2_X1 U425 ( .A(n400), .B(n372), .Z(n374) );
  XNOR2_X1 U426 ( .A(G211GAT), .B(G78GAT), .ZN(n373) );
  XNOR2_X1 U427 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U428 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n376) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U431 ( .A(n378), .B(n377), .Z(n381) );
  XNOR2_X1 U432 ( .A(n379), .B(G64GAT), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U434 ( .A(n383), .B(n382), .ZN(n555) );
  XNOR2_X1 U435 ( .A(n555), .B(KEYINPUT106), .ZN(n572) );
  NOR2_X1 U436 ( .A1(n384), .A2(n572), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n385), .B(KEYINPUT107), .ZN(n386) );
  NOR2_X1 U438 ( .A1(n558), .A2(n386), .ZN(n387) );
  XNOR2_X1 U439 ( .A(KEYINPUT47), .B(n387), .ZN(n396) );
  INV_X1 U440 ( .A(n388), .ZN(n392) );
  INV_X1 U441 ( .A(KEYINPUT36), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n389), .B(n558), .ZN(n482) );
  INV_X1 U443 ( .A(n555), .ZN(n585) );
  NOR2_X1 U444 ( .A1(n482), .A2(n585), .ZN(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT45), .B(n390), .Z(n391) );
  NOR2_X1 U446 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n393), .B(KEYINPUT108), .ZN(n394) );
  INV_X1 U448 ( .A(n563), .ZN(n577) );
  NAND2_X1 U449 ( .A1(n394), .A2(n577), .ZN(n395) );
  NAND2_X1 U450 ( .A1(n396), .A2(n395), .ZN(n398) );
  XOR2_X1 U451 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U453 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U454 ( .A(n404), .B(n403), .Z(n410) );
  XOR2_X1 U455 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n406) );
  XNOR2_X1 U456 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n405) );
  XNOR2_X1 U457 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U458 ( .A(G169GAT), .B(n407), .Z(n437) );
  XNOR2_X1 U459 ( .A(n437), .B(n408), .ZN(n409) );
  XNOR2_X1 U460 ( .A(n410), .B(n409), .ZN(n505) );
  XNOR2_X1 U461 ( .A(n505), .B(KEYINPUT119), .ZN(n411) );
  NOR2_X1 U462 ( .A1(n529), .A2(n411), .ZN(n413) );
  XOR2_X1 U463 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n415) );
  XNOR2_X1 U464 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n414) );
  XNOR2_X1 U465 ( .A(n415), .B(n414), .ZN(n433) );
  XOR2_X1 U466 ( .A(G85GAT), .B(G162GAT), .Z(n417) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(G148GAT), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U469 ( .A(KEYINPUT5), .B(G57GAT), .Z(n419) );
  XNOR2_X1 U470 ( .A(G1GAT), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U472 ( .A(n421), .B(n420), .Z(n431) );
  XNOR2_X1 U473 ( .A(G127GAT), .B(G134GAT), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n422), .B(KEYINPUT0), .ZN(n423) );
  XOR2_X1 U475 ( .A(n423), .B(KEYINPUT78), .Z(n425) );
  XNOR2_X1 U476 ( .A(G113GAT), .B(G120GAT), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n436) );
  XOR2_X1 U478 ( .A(n426), .B(KEYINPUT1), .Z(n428) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n436), .B(n429), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n433), .B(n432), .ZN(n516) );
  NAND2_X1 U484 ( .A1(n434), .A2(n516), .ZN(n575) );
  NOR2_X1 U485 ( .A1(n463), .A2(n575), .ZN(n435) );
  XNOR2_X1 U486 ( .A(n435), .B(KEYINPUT55), .ZN(n451) );
  XNOR2_X1 U487 ( .A(n437), .B(n436), .ZN(n450) );
  XOR2_X1 U488 ( .A(G99GAT), .B(G190GAT), .Z(n439) );
  XNOR2_X1 U489 ( .A(G15GAT), .B(G43GAT), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U492 ( .A(G183GAT), .B(G176GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n448) );
  XOR2_X1 U495 ( .A(KEYINPUT65), .B(KEYINPUT80), .Z(n445) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U498 ( .A(KEYINPUT79), .B(n446), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n521) );
  NAND2_X1 U501 ( .A1(n571), .A2(n558), .ZN(n455) );
  XOR2_X1 U502 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n453) );
  INV_X1 U503 ( .A(G190GAT), .ZN(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT34), .B(KEYINPUT92), .Z(n473) );
  NAND2_X1 U505 ( .A1(n388), .A2(n563), .ZN(n456) );
  XNOR2_X1 U506 ( .A(n456), .B(KEYINPUT74), .ZN(n487) );
  INV_X1 U507 ( .A(n521), .ZN(n531) );
  XNOR2_X1 U508 ( .A(n463), .B(KEYINPUT28), .ZN(n508) );
  NOR2_X1 U509 ( .A1(n516), .A2(n508), .ZN(n458) );
  XOR2_X1 U510 ( .A(n505), .B(KEYINPUT27), .Z(n461) );
  INV_X1 U511 ( .A(n461), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n458), .A2(n457), .ZN(n530) );
  XNOR2_X1 U513 ( .A(KEYINPUT90), .B(n530), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n531), .A2(n459), .ZN(n468) );
  INV_X1 U515 ( .A(n516), .ZN(n546) );
  NAND2_X1 U516 ( .A1(n463), .A2(n521), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT26), .ZN(n574) );
  NOR2_X1 U518 ( .A1(n574), .A2(n461), .ZN(n545) );
  INV_X1 U519 ( .A(n505), .ZN(n519) );
  NOR2_X1 U520 ( .A1(n521), .A2(n519), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NOR2_X1 U523 ( .A1(n545), .A2(n465), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n546), .A2(n466), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n483) );
  NOR2_X1 U526 ( .A1(n558), .A2(n585), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  NOR2_X1 U528 ( .A1(n483), .A2(n470), .ZN(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT91), .B(n471), .ZN(n502) );
  NOR2_X1 U530 ( .A1(n487), .A2(n502), .ZN(n479) );
  NAND2_X1 U531 ( .A1(n479), .A2(n546), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n474), .Z(G1324GAT) );
  NAND2_X1 U534 ( .A1(n479), .A2(n505), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT93), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U537 ( .A1(n479), .A2(n531), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NAND2_X1 U540 ( .A1(n508), .A2(n479), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT94), .ZN(n481) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  NOR2_X1 U543 ( .A1(n555), .A2(n483), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT95), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n482), .A2(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n486), .ZN(n514) );
  NOR2_X1 U547 ( .A1(n487), .A2(n514), .ZN(n489) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(KEYINPUT96), .Z(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n498) );
  NOR2_X1 U550 ( .A1(n516), .A2(n498), .ZN(n491) );
  XNOR2_X1 U551 ( .A(KEYINPUT97), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NOR2_X1 U554 ( .A1(n519), .A2(n498), .ZN(n493) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(n493), .Z(n494) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  NOR2_X1 U557 ( .A1(n521), .A2(n498), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT99), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  INV_X1 U561 ( .A(n508), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n525), .A2(n498), .ZN(n499) );
  XOR2_X1 U563 ( .A(KEYINPUT100), .B(n499), .Z(n500) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  NAND2_X1 U566 ( .A1(n577), .A2(n501), .ZN(n513) );
  NOR2_X1 U567 ( .A1(n513), .A2(n502), .ZN(n509) );
  NAND2_X1 U568 ( .A1(n546), .A2(n509), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n509), .A2(n505), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n531), .A2(n509), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n512), .Z(G1335GAT) );
  NOR2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U579 ( .A(KEYINPUT102), .B(n515), .Z(n524) );
  NOR2_X1 U580 ( .A1(n524), .A2(n516), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT103), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n524), .A2(n519), .ZN(n520) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n524), .ZN(n522) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(n522), .Z(n523) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  XNOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT105), .ZN(n527) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n529), .A2(n530), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n534) );
  NOR2_X1 U594 ( .A1(n577), .A2(n534), .ZN(n533) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  INV_X1 U596 ( .A(n534), .ZN(n542) );
  AND2_X1 U597 ( .A1(n501), .A2(n542), .ZN(n539) );
  XOR2_X1 U598 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n536) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT110), .B(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n572), .A2(n542), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U607 ( .A1(n542), .A2(n558), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT113), .Z(n549) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U611 ( .A1(n529), .A2(n547), .ZN(n559) );
  NAND2_X1 U612 ( .A1(n559), .A2(n563), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n551) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(n552), .Z(n554) );
  NAND2_X1 U618 ( .A1(n559), .A2(n501), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n559), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n561) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  XOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U628 ( .A1(n571), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT122), .B(n568), .Z(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n501), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U639 ( .A(n576), .B(KEYINPUT125), .ZN(n587) );
  NOR2_X1 U640 ( .A1(n577), .A2(n587), .ZN(n582) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n579) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT126), .B(n580), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n388), .A2(n587), .ZN(n584) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n482), .A2(n587), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

