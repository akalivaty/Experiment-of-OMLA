//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1322, new_n1323, new_n1324, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1380, new_n1381, new_n1382;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n213), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n216), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G200), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT76), .B(KEYINPUT13), .Z(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G226), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT75), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n255), .A2(KEYINPUT75), .A3(G226), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G97), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n255), .A2(G232), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n254), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n252), .B2(new_n253), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n271), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n254), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n273), .B1(G238), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n251), .B1(new_n266), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n264), .B1(new_n259), .B2(new_n260), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n250), .C1(new_n280), .C2(new_n254), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n249), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G13), .A3(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G68), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT12), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G68), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n210), .A2(G33), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n209), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n284), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n295), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT71), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n210), .B2(G1), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n283), .A2(KEYINPUT71), .A3(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(G68), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n287), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT11), .B1(new_n293), .B2(new_n295), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT78), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n304), .A2(KEYINPUT78), .A3(new_n305), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n282), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n281), .A2(G190), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT13), .B1(new_n266), .B2(new_n278), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT77), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AND4_X1   g0114(.A1(KEYINPUT77), .A2(new_n313), .A3(new_n281), .A4(G190), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n295), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT15), .B(G87), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT74), .ZN(new_n319));
  INV_X1    g0119(.A(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT8), .B(G58), .Z(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n317), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n298), .A2(G77), .A3(new_n302), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G77), .B2(new_n284), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G244), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n272), .B1(new_n275), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(G107), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n331), .B1(new_n332), .B2(new_n255), .C1(new_n263), .C2(G1698), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G169), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n328), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(G190), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n328), .B(new_n341), .C1(new_n249), .C2(new_n335), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G223), .A2(G1698), .ZN(new_n344));
  INV_X1    g0144(.A(G222), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n255), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n291), .B2(new_n255), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT68), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n254), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n349), .B2(new_n348), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n273), .B1(G226), .B2(new_n276), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n323), .A2(new_n321), .B1(G150), .B2(new_n288), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n203), .A2(G20), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n317), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT69), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n358), .A2(new_n359), .B1(new_n202), .B2(new_n297), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n356), .A2(new_n357), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT69), .B1(new_n361), .B2(new_n317), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n302), .A2(G50), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT72), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT70), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n297), .B2(new_n295), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n209), .A4(new_n294), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n360), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n351), .A2(new_n338), .A3(new_n352), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n355), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT73), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n355), .A2(new_n374), .A3(new_n370), .A4(new_n371), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n343), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n353), .A2(G200), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n351), .A2(G190), .A3(new_n352), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n360), .A2(new_n362), .A3(new_n369), .A4(KEYINPUT9), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT9), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n370), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n383), .A2(new_n381), .A3(new_n377), .A4(new_n378), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT10), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n354), .B1(new_n279), .B2(new_n281), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT14), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n313), .A2(G179), .A3(new_n281), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n310), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AND4_X1   g0193(.A1(new_n316), .A2(new_n376), .A3(new_n387), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G33), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n398), .A2(KEYINPUT79), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n255), .B2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(G20), .B1(new_n396), .B2(new_n397), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT79), .B1(new_n403), .B2(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G58), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n289), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n407), .A2(new_n201), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(G20), .B1(G159), .B2(new_n288), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n409), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT81), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT81), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n396), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n397), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n400), .A2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n395), .A2(G33), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n210), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT80), .B1(new_n420), .B2(new_n400), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n403), .A2(new_n422), .A3(KEYINPUT7), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n418), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n411), .B1(new_n424), .B2(G68), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n295), .B(new_n410), .C1(new_n425), .C2(KEYINPUT16), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n283), .A2(KEYINPUT71), .A3(G20), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT71), .B1(new_n283), .B2(G20), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT8), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G58), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n406), .A2(KEYINPUT8), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n427), .A2(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT82), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT82), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n323), .A2(new_n302), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n368), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n323), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n297), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT83), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n441), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n256), .A2(G226), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n255), .B(new_n444), .C1(G223), .C2(G1698), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G87), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n254), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G232), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n272), .B1(new_n275), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G190), .ZN(new_n451));
  OAI21_X1  g0251(.A(G200), .B1(new_n447), .B2(new_n449), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n426), .A2(new_n443), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n424), .A2(G68), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT16), .B1(new_n458), .B2(new_n409), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n410), .A2(new_n295), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n443), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n426), .A2(KEYINPUT84), .A3(new_n443), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n450), .A2(G179), .ZN(new_n465));
  OAI21_X1  g0265(.A(G169), .B1(new_n447), .B2(new_n449), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n457), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n469), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n463), .A2(new_n464), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n455), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n394), .B1(new_n473), .B2(KEYINPUT86), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT86), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n455), .C1(new_n470), .C2(new_n472), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT95), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT94), .A2(KEYINPUT23), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G20), .A3(new_n332), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n210), .A2(G107), .B1(KEYINPUT94), .B2(KEYINPUT23), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT94), .A2(KEYINPUT23), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT88), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT88), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G116), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n292), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n478), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n486), .A2(G116), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n484), .A2(KEYINPUT88), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n321), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n482), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n210), .A2(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n479), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT95), .A4(new_n481), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n255), .A2(new_n210), .A3(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT22), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT22), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n255), .A2(new_n500), .A3(new_n210), .A4(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT24), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n497), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n317), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n332), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT25), .B1(new_n297), .B2(new_n332), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n283), .A2(G33), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n284), .A2(new_n511), .A3(new_n209), .A4(new_n294), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n509), .A2(new_n510), .B1(new_n332), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT96), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n506), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n505), .B1(new_n497), .B2(new_n502), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n295), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT96), .ZN(new_n518));
  INV_X1    g0318(.A(new_n513), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n270), .A2(G1), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  NOR2_X1   g0322(.A1(KEYINPUT5), .A2(G41), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(G264), .A3(new_n254), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n219), .A2(new_n256), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n221), .A2(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n396), .A2(new_n527), .A3(new_n397), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G294), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n254), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n524), .A2(new_n334), .A3(new_n267), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n526), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G179), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n354), .B2(new_n533), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n514), .A2(new_n520), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(G190), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n526), .A2(new_n531), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n283), .A2(G45), .ZN(new_n539));
  OR2_X1    g0339(.A1(KEYINPUT5), .A2(G41), .ZN(new_n540));
  NAND2_X1  g0340(.A1(KEYINPUT5), .A2(G41), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n268), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G200), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n517), .A2(new_n519), .A3(new_n537), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n334), .B1(new_n521), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(G270), .B1(new_n268), .B2(new_n542), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n396), .A2(new_n397), .A3(G257), .A4(new_n256), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n396), .A2(new_n397), .A3(G264), .A4(G1698), .ZN(new_n551));
  INV_X1    g0351(.A(G303), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n255), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n334), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G13), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(G1), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n557), .A2(new_n485), .A3(new_n487), .A4(G20), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n512), .B2(new_n484), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(G20), .B1(G33), .B2(G283), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n320), .A2(G97), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(new_n294), .B2(new_n209), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n485), .A2(new_n487), .A3(G20), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT20), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT92), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n555), .A2(new_n567), .A3(new_n568), .A4(G169), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n354), .B1(new_n549), .B2(new_n554), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n572), .B2(new_n567), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT93), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n555), .A2(new_n567), .A3(G169), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT92), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT93), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(new_n570), .A4(new_n569), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n567), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n549), .A2(new_n554), .A3(G179), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n567), .B1(new_n555), .B2(G200), .ZN(new_n585));
  INV_X1    g0385(.A(G190), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(new_n555), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n297), .A2(new_n220), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n512), .B2(new_n220), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n288), .A2(G77), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT6), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n593), .A2(new_n220), .A3(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(G97), .B(G107), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n596), .B2(new_n210), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n424), .B2(G107), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n591), .B1(new_n598), .B2(new_n317), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n524), .A2(G257), .A3(new_n254), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n543), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n396), .A2(new_n397), .A3(G244), .A4(new_n256), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n255), .A2(KEYINPUT4), .A3(G244), .A4(new_n256), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G283), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n255), .A2(G250), .A3(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n604), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n608), .B2(new_n334), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(G169), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n334), .ZN(new_n613));
  INV_X1    g0413(.A(new_n601), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n612), .B1(new_n615), .B2(G179), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n609), .A2(KEYINPUT87), .A3(new_n338), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n599), .A2(new_n611), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n609), .A2(G190), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n609), .A2(new_n249), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n595), .A2(new_n593), .ZN(new_n622));
  INV_X1    g0422(.A(new_n594), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(G20), .B1(G77), .B2(new_n288), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n422), .B1(new_n403), .B2(KEYINPUT7), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT80), .B(new_n400), .C1(new_n255), .C2(G20), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n416), .B2(new_n417), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n628), .B2(new_n332), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n590), .B1(new_n629), .B2(new_n295), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n485), .A2(new_n487), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G33), .ZN(new_n633));
  OR2_X1    g0433(.A1(G238), .A2(G1698), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n329), .A2(G1698), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n396), .A2(new_n634), .A3(new_n397), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n334), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n219), .B1(new_n283), .B2(G45), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n268), .A2(new_n521), .B1(new_n254), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(G169), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  NOR2_X1   g0442(.A1(G238), .A2(G1698), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n329), .B2(G1698), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n644), .A2(new_n255), .B1(new_n632), .B2(G33), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n640), .B1(new_n645), .B2(new_n254), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n646), .B2(G179), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n254), .B1(new_n633), .B2(new_n636), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n268), .A2(new_n521), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n254), .A2(new_n639), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(KEYINPUT89), .A3(new_n338), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n641), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n396), .A2(new_n397), .A3(new_n210), .A4(G68), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT91), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT19), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n655), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n255), .A2(KEYINPUT91), .A3(new_n210), .A4(G68), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n210), .B1(new_n262), .B2(new_n657), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n218), .A2(new_n220), .A3(new_n332), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n659), .B(new_n660), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n295), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT74), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n318), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n318), .A2(new_n668), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n284), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n512), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n319), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n512), .A2(new_n218), .ZN(new_n676));
  AOI211_X1 g0476(.A(new_n676), .B(new_n671), .C1(new_n666), .C2(new_n295), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n586), .B(new_n640), .C1(new_n645), .C2(new_n254), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n652), .B2(G200), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n654), .A2(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n618), .A2(new_n631), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n588), .A2(new_n681), .ZN(new_n682));
  AND4_X1   g0482(.A1(new_n477), .A2(new_n536), .A3(new_n546), .A4(new_n682), .ZN(G372));
  NAND2_X1  g0483(.A1(new_n373), .A2(new_n375), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n461), .A2(new_n467), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT18), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n316), .A2(new_n339), .A3(new_n337), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n393), .ZN(new_n688));
  INV_X1    g0488(.A(new_n455), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n387), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n468), .A2(new_n469), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n472), .A3(new_n456), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n689), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n475), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n473), .A2(KEYINPUT86), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n394), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n646), .A2(G179), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n641), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n677), .A2(new_n679), .B1(new_n675), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n546), .A2(new_n618), .A3(new_n631), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n583), .B1(new_n574), .B2(new_n578), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n517), .A2(new_n519), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n535), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n703), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n676), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n679), .A2(new_n672), .A3(new_n667), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n641), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT89), .B1(new_n652), .B2(new_n338), .ZN(new_n711));
  NOR4_X1   g0511(.A1(new_n648), .A2(new_n651), .A3(new_n642), .A4(G179), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI221_X4 g0513(.A(new_n671), .B1(new_n673), .B2(new_n319), .C1(new_n666), .C2(new_n295), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT26), .B1(new_n618), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n675), .A2(new_n701), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT26), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n630), .A2(new_n610), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n609), .A2(KEYINPUT87), .A3(new_n338), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT87), .B1(new_n609), .B2(new_n338), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n702), .A2(new_n718), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n716), .A2(new_n717), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT97), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT97), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n716), .A2(new_n723), .A3(new_n726), .A4(new_n717), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n707), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n693), .B1(new_n699), .B2(new_n728), .ZN(G369));
  INV_X1    g0529(.A(new_n704), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n557), .A2(new_n210), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT27), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT27), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G213), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G343), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n580), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n730), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n588), .B2(new_n738), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n514), .A2(new_n520), .A3(new_n736), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n536), .A2(new_n743), .A3(new_n546), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n536), .B2(new_n737), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n536), .A2(new_n546), .A3(new_n737), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n730), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(new_n706), .B2(new_n736), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n747), .A2(new_n750), .ZN(G399));
  NOR2_X1   g0551(.A1(new_n663), .A2(G116), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n214), .A2(new_n269), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(G1), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n207), .B2(new_n753), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT29), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n704), .A2(new_n536), .ZN(new_n758));
  AND4_X1   g0558(.A1(new_n546), .A2(new_n618), .A3(new_n631), .A4(new_n702), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n717), .A2(new_n709), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT26), .B1(new_n618), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n680), .A2(new_n718), .A3(new_n719), .A4(new_n722), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n762), .A2(new_n717), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n757), .B1(new_n765), .B2(new_n737), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n725), .A2(new_n727), .ZN(new_n767));
  INV_X1    g0567(.A(new_n707), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n736), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n766), .B1(new_n769), .B2(new_n757), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT98), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n613), .A2(new_n538), .A3(new_n652), .A4(new_n614), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n772), .B2(new_n582), .ZN(new_n773));
  INV_X1    g0573(.A(new_n582), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G250), .A2(G1698), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n221), .B2(G1698), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(new_n255), .B1(G33), .B2(G294), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n525), .B1(new_n777), .B2(new_n254), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n646), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n774), .A2(KEYINPUT98), .A3(new_n779), .A4(new_n609), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT99), .B(KEYINPUT30), .Z(new_n781));
  NAND3_X1  g0581(.A1(new_n773), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n772), .A2(new_n582), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT30), .ZN(new_n784));
  AND3_X1   g0584(.A1(new_n555), .A2(new_n338), .A3(new_n646), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT100), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n615), .B2(new_n544), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n609), .A2(new_n533), .A3(KEYINPUT100), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n782), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n736), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT31), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n615), .A2(new_n786), .A3(new_n544), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT100), .B1(new_n609), .B2(new_n533), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(new_n785), .B1(new_n783), .B2(KEYINPUT30), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n737), .B1(new_n797), .B2(new_n782), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT31), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n719), .A2(new_n722), .B1(new_n621), .B2(new_n630), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n704), .A2(new_n587), .A3(new_n680), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n536), .A2(new_n546), .A3(new_n737), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n793), .B(new_n799), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G330), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n770), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n756), .B1(new_n805), .B2(G1), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT101), .ZN(G364));
  NOR2_X1   g0607(.A1(new_n556), .A2(G20), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n283), .B1(new_n808), .B2(G45), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n753), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n742), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(G330), .B2(new_n740), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n255), .A2(new_n214), .ZN(new_n815));
  INV_X1    g0615(.A(G355), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n816), .B1(G116), .B2(new_n214), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n247), .A2(G45), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n398), .A2(new_n214), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n270), .B2(new_n208), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n817), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G13), .A2(G33), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n209), .B1(G20), .B2(new_n354), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n812), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n210), .A2(new_n338), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G200), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n586), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(G190), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n202), .A2(new_n832), .B1(new_n834), .B2(new_n289), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n338), .A2(new_n249), .A3(G190), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G20), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n220), .ZN(new_n839));
  NOR2_X1   g0639(.A1(G190), .A2(G200), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n829), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n255), .B1(new_n841), .B2(new_n291), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n835), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n829), .A2(G190), .A3(new_n249), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT102), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(G58), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n210), .A2(G179), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(G190), .A3(G200), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT103), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(G87), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT32), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(new_n840), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n858), .B2(G159), .ZN(new_n859));
  INV_X1    g0659(.A(G159), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n857), .A2(KEYINPUT32), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n848), .A2(new_n586), .A3(G200), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n332), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n859), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n843), .A2(new_n847), .A3(new_n855), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n853), .A2(new_n552), .ZN(new_n866));
  INV_X1    g0666(.A(G322), .ZN(new_n867));
  INV_X1    g0667(.A(G311), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n844), .A2(new_n867), .B1(new_n841), .B2(new_n868), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n255), .B(new_n869), .C1(G329), .C2(new_n858), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n831), .A2(G326), .B1(G294), .B2(new_n837), .ZN(new_n871));
  XNOR2_X1  g0671(.A(KEYINPUT33), .B(G317), .ZN(new_n872));
  INV_X1    g0672(.A(new_n862), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n833), .A2(new_n872), .B1(new_n873), .B2(G283), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n865), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n828), .B1(new_n876), .B2(new_n825), .ZN(new_n877));
  INV_X1    g0677(.A(new_n824), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n740), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n814), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(G396));
  OAI21_X1  g0681(.A(new_n736), .B1(new_n325), .B2(new_n327), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n342), .A2(new_n882), .B1(new_n337), .B2(new_n339), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n337), .A2(new_n339), .A3(new_n737), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT105), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n342), .A2(new_n882), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n340), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n769), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT106), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT106), .B1(new_n886), .B2(new_n890), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n769), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n812), .B1(new_n896), .B2(new_n804), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n804), .B2(new_n896), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n825), .A2(new_n822), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n812), .B1(G77), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(G283), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n834), .A2(new_n901), .B1(new_n218), .B2(new_n862), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n839), .B(new_n902), .C1(G303), .C2(new_n831), .ZN(new_n903));
  INV_X1    g0703(.A(new_n632), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n904), .A2(new_n841), .B1(new_n868), .B2(new_n857), .ZN(new_n905));
  INV_X1    g0705(.A(new_n844), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n255), .B(new_n905), .C1(G294), .C2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n903), .B(new_n907), .C1(new_n332), .C2(new_n853), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT104), .ZN(new_n909));
  INV_X1    g0709(.A(new_n841), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n831), .A2(G137), .B1(new_n910), .B2(G159), .ZN(new_n911));
  INV_X1    g0711(.A(G150), .ZN(new_n912));
  INV_X1    g0712(.A(G143), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n911), .B1(new_n912), .B2(new_n834), .C1(new_n845), .C2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT34), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n862), .A2(new_n289), .ZN(new_n918));
  INV_X1    g0718(.A(G132), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n255), .B1(new_n857), .B2(new_n919), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n918), .B(new_n920), .C1(G58), .C2(new_n837), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n917), .B(new_n921), .C1(new_n202), .C2(new_n853), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n909), .B1(new_n916), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n900), .B1(new_n923), .B2(new_n825), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n891), .B2(new_n823), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n898), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(G384));
  OR2_X1    g0727(.A1(new_n624), .A2(KEYINPUT35), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n624), .A2(KEYINPUT35), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n928), .A2(G116), .A3(new_n211), .A4(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  OR3_X1    g0732(.A1(new_n207), .A2(new_n291), .A3(new_n407), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n202), .A2(G68), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n283), .B(G13), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n426), .A2(KEYINPUT84), .A3(new_n443), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT84), .B1(new_n426), .B2(new_n443), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n734), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n685), .A2(new_n453), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT37), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT108), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n734), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n463), .A2(new_n464), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT37), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n468), .A2(new_n945), .A3(new_n946), .A4(new_n453), .ZN(new_n947));
  AND4_X1   g0747(.A1(new_n426), .A2(new_n443), .A3(new_n451), .A4(new_n452), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n426), .A2(new_n443), .B1(new_n466), .B2(new_n465), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n946), .B1(new_n950), .B2(new_n945), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT108), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n943), .A2(new_n947), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n939), .B1(new_n686), .B2(new_n455), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT16), .B1(new_n405), .B2(new_n409), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n438), .B(new_n436), .C1(new_n460), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n944), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n695), .B2(new_n689), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT38), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n467), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n961), .A3(new_n453), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT37), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n947), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n959), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n955), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n310), .A2(new_n736), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n393), .A2(new_n316), .A3(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n310), .B(new_n736), .C1(new_n390), .C2(new_n392), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n891), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n682), .A2(new_n748), .B1(KEYINPUT31), .B2(new_n798), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT110), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n791), .B2(new_n792), .ZN(new_n974));
  AOI211_X1 g0774(.A(KEYINPUT110), .B(KEYINPUT31), .C1(new_n790), .C2(new_n736), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n972), .A2(new_n976), .A3(KEYINPUT111), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT111), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT110), .B1(new_n798), .B2(KEYINPUT31), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n791), .A2(new_n973), .A3(new_n792), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n971), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT40), .B1(new_n966), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n960), .B1(new_n959), .B2(new_n964), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n947), .A2(new_n963), .ZN(new_n988));
  OAI211_X1 g0788(.A(KEYINPUT38), .B(new_n988), .C1(new_n473), .C2(new_n958), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT40), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(new_n991), .A3(new_n984), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n977), .A2(new_n983), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(new_n477), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G330), .ZN(new_n997));
  INV_X1    g0797(.A(new_n995), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n993), .A2(new_n699), .A3(new_n998), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n970), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n892), .B2(new_n884), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n1002), .A2(new_n990), .B1(new_n686), .B2(new_n734), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT39), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n955), .B2(new_n965), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n393), .A2(new_n736), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n987), .A2(KEYINPUT39), .A3(new_n989), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT109), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n770), .B2(new_n699), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n717), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n680), .A2(new_n719), .A3(new_n722), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(new_n1014), .B2(KEYINPUT26), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n726), .B1(new_n1015), .B2(new_n723), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n727), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n768), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n757), .A3(new_n737), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n765), .A2(new_n737), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT29), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n477), .A3(KEYINPUT109), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n692), .B1(new_n1012), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1010), .B(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1000), .A2(new_n1025), .B1(new_n283), .B2(new_n808), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1000), .A2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n936), .B1(new_n1026), .B2(new_n1027), .ZN(G367));
  OAI21_X1  g0828(.A(new_n800), .B1(new_n630), .B2(new_n737), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n618), .B2(new_n737), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n749), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT42), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1031), .A2(new_n536), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n736), .B1(new_n1035), .B2(new_n618), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT43), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n677), .A2(new_n737), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1013), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n761), .B2(new_n1038), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1034), .A2(new_n1036), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1037), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n746), .A2(new_n1031), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT113), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1044), .A2(KEYINPUT113), .A3(new_n1045), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n753), .B(KEYINPUT41), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1031), .A2(new_n750), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n1052));
  XNOR2_X1  g0852(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1031), .A2(new_n750), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT44), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n1053), .A2(new_n1055), .A3(new_n747), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n747), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n704), .A2(new_n736), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n749), .B1(new_n745), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(new_n741), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n805), .A2(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1050), .B1(new_n1064), .B2(new_n805), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1048), .B(new_n1049), .C1(new_n810), .C2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n239), .A2(new_n819), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n319), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n826), .B1(new_n1068), .B2(new_n214), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n812), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n844), .A2(new_n912), .B1(new_n841), .B2(new_n202), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n398), .B(new_n1071), .C1(G137), .C2(new_n858), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n854), .A2(G58), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n838), .A2(new_n289), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G143), .B2(new_n831), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n833), .A2(G159), .B1(new_n873), .B2(G77), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G317), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n398), .B1(new_n857), .B2(new_n1078), .C1(new_n841), .C2(new_n901), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n846), .B2(G303), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n854), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n873), .A2(G97), .B1(new_n837), .B2(G107), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G294), .A2(new_n833), .B1(new_n831), .B2(G311), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT46), .B1(new_n854), .B2(new_n632), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT47), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1070), .B1(new_n1087), .B2(new_n825), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1040), .B2(new_n878), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(G387));
  AOI21_X1  g0890(.A(new_n753), .B1(new_n805), .B2(new_n1062), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n805), .B2(new_n1062), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n745), .A2(new_n878), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n815), .A2(new_n752), .B1(G107), .B2(new_n214), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n235), .A2(G45), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n323), .A2(new_n202), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT50), .Z(new_n1097));
  INV_X1    g0897(.A(new_n752), .ZN(new_n1098));
  AOI211_X1 g0898(.A(G45), .B(new_n1098), .C1(G68), .C2(G77), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n819), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1094), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n812), .B1(new_n1101), .B2(new_n827), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n832), .A2(new_n860), .B1(new_n220), .B2(new_n862), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n323), .B2(new_n833), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n854), .A2(G77), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n319), .A2(new_n837), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n844), .A2(new_n202), .B1(new_n857), .B2(new_n912), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n398), .B(new_n1107), .C1(G68), .C2(new_n910), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n255), .B1(new_n858), .B2(G326), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n833), .A2(G311), .B1(new_n910), .B2(G303), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n867), .B2(new_n832), .C1(new_n845), .C2(new_n1078), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT48), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n854), .A2(G294), .B1(G283), .B2(new_n837), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT49), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1110), .B1(new_n904), .B2(new_n862), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1109), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1102), .B1(new_n1121), .B2(new_n825), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1062), .A2(new_n810), .B1(new_n1093), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1092), .A2(new_n1123), .ZN(G393));
  NAND2_X1  g0924(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1064), .A2(new_n811), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1058), .A2(new_n809), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1031), .A2(new_n824), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n244), .A2(new_n214), .A3(new_n398), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n826), .B1(new_n220), .B2(new_n214), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n812), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n832), .A2(new_n1078), .B1(new_n868), .B2(new_n844), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT52), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n863), .B1(new_n632), .B2(new_n837), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n552), .B2(new_n834), .ZN(new_n1135));
  INV_X1    g0935(.A(G294), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n398), .B1(new_n857), .B2(new_n867), .C1(new_n841), .C2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1133), .B(new_n1138), .C1(new_n901), .C2(new_n853), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n833), .A2(G50), .B1(new_n910), .B2(new_n323), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT115), .Z(new_n1141));
  OAI221_X1 g0941(.A(new_n255), .B1(new_n857), .B2(new_n913), .C1(new_n218), .C2(new_n862), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G77), .B2(new_n837), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(new_n289), .C2(new_n853), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G150), .A2(new_n831), .B1(new_n906), .B2(G159), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT51), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1139), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1131), .B1(new_n1147), .B2(new_n825), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1127), .B1(new_n1128), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1126), .A2(new_n1149), .ZN(G390));
  AOI21_X1  g0950(.A(new_n736), .B1(new_n760), .B2(new_n764), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n885), .B1(new_n1151), .B2(new_n891), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n970), .A2(new_n803), .A3(G330), .A4(new_n891), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(G330), .B1(new_n893), .B2(new_n894), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n977), .B2(new_n983), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1154), .B1(new_n1156), .B2(new_n970), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n803), .A2(G330), .A3(new_n891), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n984), .A2(G330), .B1(new_n1001), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n891), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n728), .A2(new_n736), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(new_n885), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n376), .A2(new_n387), .A3(new_n393), .A4(new_n316), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n696), .B2(new_n475), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n995), .A2(G330), .A3(new_n698), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT116), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n477), .A2(new_n995), .A3(KEYINPUT116), .A4(G330), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1163), .A2(new_n1170), .A3(new_n1024), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT117), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1163), .A2(new_n1170), .A3(new_n1024), .A4(KEYINPUT117), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT119), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n985), .A2(new_n997), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n970), .B1(new_n1161), .B2(new_n885), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1005), .A2(new_n1008), .B1(new_n1006), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1006), .B1(new_n1152), .B2(new_n1001), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n966), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1177), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1006), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n947), .B1(new_n951), .B2(KEYINPUT108), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n941), .A2(new_n942), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n954), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n960), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT39), .B1(new_n1187), .B2(new_n989), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n987), .A2(KEYINPUT39), .A3(new_n989), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n966), .A2(new_n1180), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1153), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1182), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT119), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1173), .A2(new_n1194), .A3(new_n1174), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1176), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1193), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1175), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(KEYINPUT118), .A3(new_n811), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT118), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n1201), .B2(new_n753), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1196), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1197), .A2(new_n810), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n822), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n812), .B1(new_n323), .B2(new_n899), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n854), .A2(G150), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT53), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n398), .B1(new_n858), .B2(G125), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT54), .B(G143), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1209), .B1(new_n919), .B2(new_n844), .C1(new_n841), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G137), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n834), .A2(new_n1212), .B1(new_n860), .B2(new_n838), .ZN(new_n1213));
  INV_X1    g1013(.A(G128), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n832), .A2(new_n1214), .B1(new_n202), .B2(new_n862), .ZN(new_n1215));
  OR3_X1    g1015(.A1(new_n1211), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1208), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n841), .A2(new_n220), .B1(new_n857), .B2(new_n1136), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n255), .B(new_n1219), .C1(G116), .C2(new_n906), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n918), .B1(G77), .B2(new_n837), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G107), .A2(new_n833), .B1(new_n831), .B2(G283), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1220), .A2(new_n855), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1217), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1206), .B1(new_n1225), .B2(new_n825), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT121), .Z(new_n1227));
  NAND2_X1  g1027(.A1(new_n1205), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1204), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1203), .A2(new_n1230), .ZN(G378));
  OAI21_X1  g1031(.A(new_n812), .B1(G50), .B2(new_n899), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n255), .A2(G41), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n901), .B2(new_n857), .C1(new_n332), .C2(new_n844), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n319), .B2(new_n910), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1074), .B1(G97), .B2(new_n833), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n831), .A2(G116), .B1(new_n873), .B2(G58), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1235), .A2(new_n1105), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT58), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1233), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT122), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n844), .A2(new_n1214), .B1(new_n841), .B2(new_n1212), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G132), .B2(new_n833), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n831), .A2(G125), .B1(G150), .B2(new_n837), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n853), .C2(new_n1210), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT123), .Z(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n873), .A2(G159), .ZN(new_n1254));
  AOI211_X1 g1054(.A(G33), .B(G41), .C1(new_n858), .C2(G124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1246), .B1(new_n1243), .B2(new_n1242), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1232), .B1(new_n1258), .B2(new_n825), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n387), .A2(new_n372), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n370), .A2(new_n944), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1260), .B(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1262), .B(new_n1263), .Z(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1259), .B1(new_n1265), .B2(new_n823), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT124), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1003), .A2(new_n1009), .A3(new_n1265), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1265), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1268), .A2(new_n1269), .B1(new_n993), .B2(new_n997), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1010), .A2(new_n1264), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n997), .B1(new_n986), .B2(new_n992), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1003), .A2(new_n1009), .A3(new_n1265), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1267), .B1(new_n1275), .B2(new_n810), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1170), .A2(new_n1024), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1198), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT57), .B1(new_n1279), .B2(new_n1275), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(KEYINPUT57), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1277), .B1(new_n1175), .B2(new_n1197), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n811), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1276), .B1(new_n1280), .B2(new_n1283), .ZN(G375));
  AND3_X1   g1084(.A1(new_n1173), .A2(new_n1194), .A3(new_n1174), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1194), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1050), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1163), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1277), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1163), .A2(new_n810), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n812), .B1(G68), .B2(new_n899), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n255), .B1(new_n857), .B2(new_n1214), .C1(new_n841), .C2(new_n912), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n846), .B2(G137), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n834), .A2(new_n1210), .B1(new_n406), .B2(new_n862), .ZN(new_n1296));
  OAI22_X1  g1096(.A1(new_n832), .A2(new_n919), .B1(new_n202), .B2(new_n838), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1295), .B(new_n1298), .C1(new_n860), .C2(new_n853), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n853), .A2(new_n220), .B1(new_n552), .B2(new_n857), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(KEYINPUT125), .Z(new_n1301));
  OAI21_X1  g1101(.A(new_n398), .B1(new_n844), .B2(new_n901), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(G107), .B2(new_n910), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n833), .A2(new_n632), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n831), .A2(G294), .B1(new_n873), .B2(G77), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1303), .A2(new_n1106), .A3(new_n1304), .A4(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1299), .B1(new_n1301), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1293), .B1(new_n1307), .B2(new_n825), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n970), .B2(new_n823), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1292), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1291), .A2(new_n1311), .ZN(G381));
  NAND3_X1  g1112(.A1(new_n1092), .A2(new_n880), .A3(new_n1123), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1126), .A2(new_n1149), .A3(new_n926), .A4(new_n1314), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(G387), .A2(G381), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n753), .B1(new_n1175), .B2(new_n1197), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1287), .A2(new_n1193), .B1(new_n1317), .B2(KEYINPUT118), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1229), .B1(new_n1318), .B2(new_n1202), .ZN(new_n1319));
  INV_X1    g1119(.A(G375), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1316), .A2(new_n1319), .A3(new_n1320), .ZN(G407));
  NAND2_X1  g1121(.A1(new_n735), .A2(G213), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1320), .A2(new_n1319), .A3(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(G407), .A2(G213), .A3(new_n1324), .ZN(G409));
  INV_X1    g1125(.A(new_n1275), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1282), .A2(new_n1326), .A3(new_n1050), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1266), .B1(new_n1326), .B2(new_n809), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1203), .B(new_n1230), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1319), .B2(G375), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT60), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n811), .B1(new_n1290), .B2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1173), .A2(KEYINPUT60), .A3(new_n1174), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1332), .B1(new_n1333), .B2(new_n1290), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(G384), .A3(new_n1311), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n926), .B1(new_n1334), .B2(new_n1310), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1330), .A2(new_n1322), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT62), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1330), .A2(new_n1322), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1323), .A2(G2897), .ZN(new_n1343));
  XOR2_X1   g1143(.A(new_n1343), .B(KEYINPUT126), .Z(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1338), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1336), .A2(new_n1337), .A3(new_n1344), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1342), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT61), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT62), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1330), .A2(new_n1351), .A3(new_n1322), .A4(new_n1339), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1341), .A2(new_n1349), .A3(new_n1350), .A4(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n880), .B1(new_n1092), .B2(new_n1123), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(G390), .A2(new_n1313), .A3(new_n1355), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1126), .B(new_n1149), .C1(new_n1314), .C2(new_n1354), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(G387), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1356), .A2(new_n1066), .A3(new_n1089), .A4(new_n1357), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1353), .A2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT127), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1342), .A2(new_n1363), .A3(new_n1348), .ZN(new_n1364));
  OAI211_X1 g1164(.A(KEYINPUT57), .B(new_n1275), .C1(new_n1201), .C2(new_n1277), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1282), .A2(new_n1326), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n811), .B(new_n1365), .C1(new_n1366), .C2(KEYINPUT57), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(G378), .A2(new_n1367), .A3(new_n1276), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1323), .B1(new_n1368), .B2(new_n1329), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1370));
  OAI21_X1  g1170(.A(KEYINPUT127), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1364), .A2(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT63), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1340), .A2(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1359), .A2(new_n1350), .A3(new_n1360), .ZN(new_n1375));
  AOI211_X1 g1175(.A(new_n1323), .B(new_n1338), .C1(new_n1368), .C2(new_n1329), .ZN(new_n1376));
  AOI21_X1  g1176(.A(new_n1375), .B1(new_n1376), .B2(KEYINPUT63), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1372), .A2(new_n1374), .A3(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1362), .A2(new_n1378), .ZN(G405));
  NAND2_X1  g1179(.A1(new_n1319), .A2(G375), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1380), .A2(new_n1368), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1381), .B(new_n1339), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(new_n1382), .B(new_n1361), .ZN(G402));
endmodule


