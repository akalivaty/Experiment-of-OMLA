//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT95), .ZN(new_n205));
  MUX2_X1   g004(.A(G1gat), .B(new_n203), .S(new_n205), .Z(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(G8gat), .Z(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G43gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT93), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n209), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT94), .B(G50gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G43gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT92), .B(G29gat), .Z(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT14), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n212), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n225), .B1(new_n212), .B2(new_n224), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(KEYINPUT17), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n206), .B(G8gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT96), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n229), .B(new_n226), .Z(new_n236));
  XOR2_X1   g035(.A(new_n233), .B(KEYINPUT13), .Z(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n231), .A2(new_n234), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n235), .A2(KEYINPUT97), .A3(new_n239), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G169gat), .B(G197gat), .Z(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(KEYINPUT12), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n245), .A2(new_n255), .A3(new_n239), .A4(new_n235), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT98), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n235), .A2(new_n239), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT98), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n255), .A4(new_n245), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G85gat), .A2(G92gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT7), .ZN(new_n265));
  INV_X1    g064(.A(G99gat), .ZN(new_n266));
  INV_X1    g065(.A(G106gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT8), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n265), .B(new_n268), .C1(G85gat), .C2(G92gat), .ZN(new_n269));
  XOR2_X1   g068(.A(G99gat), .B(G106gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n228), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n226), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT41), .ZN(new_n275));
  NAND2_X1  g074(.A1(G232gat), .A2(G233gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n272), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n275), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n283), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G78gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT9), .ZN(new_n289));
  XNOR2_X1  g088(.A(G57gat), .B(G64gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n287), .B(KEYINPUT99), .ZN(new_n292));
  INV_X1    g091(.A(new_n290), .ZN(new_n293));
  AND2_X1   g092(.A1(G71gat), .A2(G78gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n292), .B(new_n293), .C1(KEYINPUT9), .C2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n273), .A2(KEYINPUT10), .A3(new_n291), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n291), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n297), .B(new_n271), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n296), .B1(new_n299), .B2(KEYINPUT10), .ZN(new_n300));
  AND2_X1   g099(.A1(G230gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(new_n298), .B2(new_n302), .ZN(new_n304));
  XNOR2_X1  g103(.A(G120gat), .B(G148gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G176gat), .B(G204gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n304), .B(new_n307), .Z(new_n308));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n229), .B1(new_n309), .B2(new_n297), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT101), .ZN(new_n311));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(new_n312), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G155gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n315), .B(KEYINPUT20), .Z(new_n316));
  OR3_X1    g115(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n313), .B2(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n309), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT100), .B(KEYINPUT19), .Z(new_n320));
  XNOR2_X1  g119(.A(G183gat), .B(G211gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n319), .B(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n286), .B(new_n308), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  INV_X1    g126(.A(G85gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT0), .B(G57gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  XOR2_X1   g133(.A(G127gat), .B(G134gat), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT71), .B(G120gat), .ZN(new_n337));
  INV_X1    g136(.A(G113gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n338), .A2(G120gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n334), .B(new_n336), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(KEYINPUT1), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G141gat), .B(G148gat), .Z(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  INV_X1    g145(.A(G162gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(KEYINPUT2), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G141gat), .B(G148gat), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n349), .B(new_n348), .C1(new_n353), .C2(KEYINPUT2), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OR3_X1    g154(.A1(new_n344), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT4), .B1(new_n344), .B2(new_n355), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n343), .A2(new_n341), .B1(new_n355), .B2(KEYINPUT3), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n356), .A2(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n344), .B(new_n355), .ZN(new_n364));
  INV_X1    g163(.A(new_n362), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n333), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT5), .B1(new_n361), .B2(new_n362), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n332), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n364), .A2(new_n365), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n361), .B2(new_n362), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n370), .B(new_n331), .C1(new_n372), .C2(new_n333), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n367), .A2(new_n368), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT6), .A3(new_n331), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G211gat), .ZN(new_n379));
  INV_X1    g178(.A(G218gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G211gat), .A2(G218gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT22), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(G197gat), .A2(G204gat), .ZN(new_n388));
  AND2_X1   g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n381), .A2(KEYINPUT77), .A3(new_n382), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n385), .A2(KEYINPUT78), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n394));
  INV_X1    g193(.A(G197gat), .ZN(new_n395));
  INV_X1    g194(.A(G204gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G197gat), .A2(G204gat), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n397), .A2(new_n398), .B1(new_n386), .B2(new_n382), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n394), .B1(new_n399), .B2(new_n383), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n392), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G183gat), .ZN(new_n411));
  INV_X1    g210(.A(G190gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(G169gat), .A2(G176gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT23), .ZN(new_n416));
  NAND2_X1  g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(G169gat), .B2(G176gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT65), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT25), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT65), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n416), .A2(new_n417), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n414), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT70), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n411), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n429), .A3(KEYINPUT27), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n412), .A2(KEYINPUT69), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OR3_X1    g233(.A1(new_n411), .A2(KEYINPUT70), .A3(KEYINPUT27), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT27), .B(G183gat), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n431), .B2(new_n433), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n436), .A2(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n415), .A2(KEYINPUT26), .ZN(new_n441));
  NAND2_X1  g240(.A1(G183gat), .A2(G190gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n417), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n441), .B(new_n442), .C1(new_n444), .C2(new_n415), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n425), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n405), .B(KEYINPUT66), .ZN(new_n447));
  NAND2_X1  g246(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n434), .A2(new_n429), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n406), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n420), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n422), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n404), .B1(new_n446), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G226gat), .A2(G233gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n429), .A2(new_n448), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT69), .B(G190gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n453), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n405), .B(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n455), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT25), .ZN(new_n466));
  INV_X1    g265(.A(new_n445), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n411), .A2(KEYINPUT70), .A3(KEYINPUT27), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT28), .B1(new_n469), .B2(new_n430), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n439), .A2(new_n438), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n466), .A2(new_n473), .A3(new_n425), .ZN(new_n474));
  INV_X1    g273(.A(new_n458), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n403), .B1(new_n459), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n474), .B2(new_n404), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(KEYINPUT79), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n402), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481));
  INV_X1    g280(.A(new_n446), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n458), .B1(new_n482), .B2(new_n466), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n459), .A2(KEYINPUT80), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n401), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(KEYINPUT81), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n484), .A2(new_n488), .A3(new_n401), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G8gat), .B(G36gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(G64gat), .B(G92gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n487), .A2(new_n489), .A3(new_n493), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT30), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n498), .A3(new_n494), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n378), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n400), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n503), .B2(new_n392), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n355), .B1(new_n504), .B2(KEYINPUT3), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n359), .A2(new_n404), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n359), .A2(KEYINPUT83), .A3(new_n404), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n402), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G228gat), .ZN(new_n511));
  INV_X1    g310(.A(G233gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n505), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n390), .A2(new_n382), .A3(new_n381), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n399), .A2(new_n383), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT29), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n355), .B1(new_n517), .B2(KEYINPUT3), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n359), .A2(new_n404), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(new_n401), .ZN(new_n520));
  INV_X1    g319(.A(new_n513), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT82), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT82), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n514), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(G22gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n514), .B(new_n527), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G78gat), .B(G106gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G50gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n521), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n522), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n539), .A2(KEYINPUT84), .A3(new_n527), .A4(new_n514), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n535), .A2(new_n526), .A3(new_n540), .A4(new_n532), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n533), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n500), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n344), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n446), .B2(new_n456), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n466), .A2(new_n344), .A3(new_n473), .A4(new_n425), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G227gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(new_n512), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT34), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT74), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n548), .A2(new_n552), .A3(new_n549), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n559));
  XNOR2_X1  g358(.A(G15gat), .B(G43gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(G71gat), .B(G99gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT33), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n559), .B1(KEYINPUT72), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n563), .A2(new_n564), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n556), .B(new_n557), .C1(new_n566), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n569), .B(new_n563), .C1(new_n558), .C2(new_n564), .ZN(new_n573));
  AOI211_X1 g372(.A(KEYINPUT72), .B(new_n563), .C1(new_n558), .C2(new_n564), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n559), .A2(new_n573), .B1(new_n574), .B2(new_n568), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n557), .B1(new_n575), .B2(new_n556), .ZN(new_n576));
  OAI22_X1  g375(.A1(new_n572), .A2(new_n576), .B1(new_n556), .B2(new_n575), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(KEYINPUT76), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT76), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n575), .A2(new_n556), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n556), .B1(new_n566), .B2(new_n570), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT74), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n582), .B1(new_n584), .B2(new_n571), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n581), .B1(new_n585), .B2(new_n578), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT73), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n556), .B1(new_n575), .B2(new_n587), .ZN(new_n588));
  OAI221_X1 g387(.A(KEYINPUT73), .B1(new_n573), .B2(new_n559), .C1(new_n574), .C2(new_n568), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n584), .A2(new_n571), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n580), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n361), .A2(new_n362), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n593), .B(KEYINPUT39), .C1(new_n365), .C2(new_n364), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(new_n332), .C1(KEYINPUT39), .C2(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT87), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT40), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT40), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(KEYINPUT87), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n373), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n496), .A2(KEYINPUT30), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n493), .B1(new_n487), .B2(new_n489), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n499), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n499), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT79), .B1(new_n478), .B2(new_n483), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n459), .A2(new_n403), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n401), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n484), .A2(new_n402), .A3(new_n485), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT37), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n489), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n488), .B1(new_n611), .B2(new_n402), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(new_n486), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n493), .B(new_n614), .C1(new_n617), .C2(KEYINPUT37), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n617), .B2(KEYINPUT37), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT37), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n494), .B1(new_n490), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n375), .A2(new_n377), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n603), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n545), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n608), .A2(new_n627), .A3(KEYINPUT88), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT88), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n597), .A2(new_n373), .A3(new_n599), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n499), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT86), .B1(new_n497), .B2(new_n499), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n529), .A2(new_n532), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n540), .A2(new_n532), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n635), .A2(KEYINPUT85), .A3(new_n526), .A4(new_n535), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n541), .A2(new_n542), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT37), .B1(new_n487), .B2(new_n489), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n612), .A2(KEYINPUT37), .A3(new_n613), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n639), .A2(new_n640), .A3(new_n494), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n493), .B1(new_n617), .B2(KEYINPUT37), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT38), .B1(new_n490), .B2(new_n621), .ZN(new_n643));
  OAI22_X1  g442(.A1(new_n641), .A2(KEYINPUT38), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n638), .B1(new_n644), .B2(new_n625), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n629), .B1(new_n633), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n546), .B(new_n592), .C1(new_n628), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n606), .A2(new_n624), .A3(new_n607), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT89), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT35), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n638), .A2(new_n577), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n606), .A2(KEYINPUT89), .A3(new_n624), .A4(new_n607), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT90), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n587), .B1(new_n566), .B2(new_n570), .ZN(new_n656));
  INV_X1    g455(.A(new_n556), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n589), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n572), .B2(new_n576), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n638), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n655), .B(new_n651), .C1(new_n660), .C2(new_n500), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n497), .A2(new_n499), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n662), .A2(new_n624), .A3(new_n545), .A4(new_n590), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT90), .B1(new_n663), .B2(KEYINPUT35), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n654), .A2(new_n665), .ZN(new_n666));
  AOI211_X1 g465(.A(new_n263), .B(new_n326), .C1(new_n647), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n378), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(G1gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1324gat));
  NOR2_X1   g469(.A1(new_n631), .A2(new_n632), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT16), .B(G8gat), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT103), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n673), .A2(G8gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(KEYINPUT103), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n678), .A2(new_n679), .A3(new_n680), .A4(new_n681), .ZN(G1325gat));
  AOI21_X1  g481(.A(G15gat), .B1(new_n667), .B2(new_n585), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n592), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n580), .A2(new_n586), .A3(new_n591), .A4(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n667), .A2(G15gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n667), .A2(new_n638), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NAND2_X1  g492(.A1(new_n647), .A2(new_n666), .ZN(new_n694));
  INV_X1    g493(.A(new_n286), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n324), .A2(new_n325), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n308), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n698), .A2(new_n263), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n378), .A3(new_n219), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n546), .B(new_n687), .C1(new_n628), .C2(new_n646), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n286), .B1(new_n707), .B2(new_n666), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n701), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n624), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n705), .B1(new_n219), .B2(new_n713), .ZN(G1328gat));
  OAI21_X1  g513(.A(G36gat), .B1(new_n712), .B2(new_n671), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n702), .A2(new_n220), .A3(new_n672), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n716), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(KEYINPUT46), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT106), .B1(new_n716), .B2(KEYINPUT46), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n715), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(G1329gat));
  AOI21_X1  g519(.A(new_n709), .B1(new_n694), .B2(new_n695), .ZN(new_n721));
  AOI211_X1 g520(.A(KEYINPUT44), .B(new_n286), .C1(new_n707), .C2(new_n666), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n688), .B(new_n700), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G43gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n702), .A2(new_n211), .A3(new_n585), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n724), .B(new_n725), .C1(KEYINPUT107), .C2(KEYINPUT47), .ZN(new_n726));
  NAND2_X1  g525(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1330gat));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n216), .B1(new_n711), .B2(new_n638), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n702), .A2(new_n216), .A3(new_n638), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n729), .B(new_n733), .C1(new_n730), .C2(new_n731), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1331gat));
  NAND2_X1  g536(.A1(new_n698), .A2(new_n286), .ZN(new_n738));
  AOI211_X1 g537(.A(new_n738), .B(new_n308), .C1(new_n707), .C2(new_n666), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n263), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n378), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g541(.A(new_n671), .B(KEYINPUT110), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT49), .B(G64gat), .Z(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(G1333gat));
  NAND3_X1  g546(.A1(new_n740), .A2(G71gat), .A3(new_n688), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n740), .A2(new_n585), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(G71gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n740), .A2(new_n638), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n698), .A2(new_n262), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n308), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n721), .B2(new_n722), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n624), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n708), .A2(new_n759), .A3(new_n754), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n708), .B2(new_n754), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n699), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n624), .A2(G85gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n758), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT111), .ZN(G1336gat));
  OAI211_X1 g566(.A(new_n743), .B(new_n756), .C1(new_n721), .C2(new_n722), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n761), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n708), .A2(new_n759), .A3(new_n754), .ZN(new_n771));
  INV_X1    g570(.A(new_n743), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n770), .A2(new_n699), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n769), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT114), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n769), .A2(new_n774), .A3(new_n778), .A4(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n672), .B(new_n756), .C1(new_n721), .C2(new_n722), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n708), .A2(new_n754), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n760), .B2(new_n761), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n787), .A3(new_n759), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n772), .A2(G92gat), .A3(new_n308), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n784), .A2(new_n785), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n780), .A2(new_n794), .ZN(G1337gat));
  OAI21_X1  g594(.A(G99gat), .B1(new_n757), .B2(new_n687), .ZN(new_n796));
  INV_X1    g595(.A(new_n762), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n308), .A2(G99gat), .A3(new_n577), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT115), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(G1338gat));
  NAND2_X1  g599(.A1(new_n789), .A2(new_n790), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n308), .A2(G106gat), .A3(new_n545), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT116), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n757), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n267), .B1(new_n805), .B2(new_n638), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n797), .B2(new_n803), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(new_n806), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n236), .A2(new_n812), .A3(new_n238), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n236), .B2(new_n238), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n813), .B(new_n814), .C1(new_n234), .C2(new_n231), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n257), .A2(new_n260), .B1(new_n252), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n286), .A3(new_n699), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n304), .A2(new_n307), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n300), .A2(new_n302), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT54), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n303), .B1(KEYINPUT117), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n819), .A2(KEYINPUT117), .A3(KEYINPUT54), .A4(new_n303), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n307), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT55), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n823), .A2(new_n827), .A3(new_n307), .A4(new_n824), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n818), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n816), .B2(new_n286), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n262), .A2(new_n695), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n817), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n326), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n832), .A2(new_n697), .B1(new_n833), .B2(new_n263), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n834), .A2(new_n624), .A3(new_n638), .A4(new_n659), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n772), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n338), .A3(new_n262), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n697), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n263), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n652), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n743), .A2(new_n624), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n263), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n837), .A2(new_n846), .ZN(G1340gat));
  INV_X1    g646(.A(new_n337), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n836), .A2(new_n848), .A3(new_n699), .ZN(new_n849));
  OAI21_X1  g648(.A(G120gat), .B1(new_n845), .B2(new_n308), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n836), .B2(new_n698), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n698), .A2(G127gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n844), .B2(new_n853), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n672), .A2(new_n286), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n835), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT56), .Z(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n845), .B2(new_n286), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1343gat));
  NOR4_X1   g659(.A1(new_n834), .A2(new_n624), .A3(new_n545), .A4(new_n688), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n772), .ZN(new_n862));
  INV_X1    g661(.A(G141gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n262), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n840), .A2(new_n865), .A3(new_n638), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n834), .B2(new_n545), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n843), .A2(new_n688), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n263), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g670(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n871), .B(new_n872), .ZN(G1344gat));
  INV_X1    g672(.A(G148gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n874), .A3(new_n699), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n866), .A2(new_n867), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n638), .A2(new_n878), .A3(new_n865), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n834), .A2(new_n878), .A3(new_n865), .A4(new_n638), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n699), .A3(new_n868), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n876), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n876), .B(G148gat), .C1(new_n869), .C2(new_n308), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n875), .B1(new_n883), .B2(new_n885), .ZN(G1345gat));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n346), .A3(new_n697), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n698), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n346), .B2(new_n888), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n869), .B2(new_n286), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n861), .A2(new_n347), .A3(new_n856), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT121), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n671), .A2(new_n378), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n840), .A2(new_n652), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n263), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT124), .Z(new_n897));
  NAND3_X1  g696(.A1(new_n840), .A2(KEYINPUT122), .A3(new_n624), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n834), .B2(new_n378), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n898), .A2(new_n900), .A3(new_n660), .A4(new_n743), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n263), .A2(G169gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n897), .A2(new_n905), .ZN(G1348gat));
  INV_X1    g705(.A(G176gat), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n895), .A2(new_n907), .A3(new_n308), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n902), .A2(new_n699), .A3(new_n903), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n907), .ZN(G1349gat));
  OR3_X1    g709(.A1(new_n895), .A2(KEYINPUT125), .A3(new_n697), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT125), .B1(new_n895), .B2(new_n697), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n460), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n698), .A2(new_n438), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n901), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n913), .B(new_n916), .C1(new_n901), .C2(new_n914), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1350gat));
  NAND4_X1  g719(.A1(new_n902), .A2(new_n434), .A3(new_n695), .A4(new_n903), .ZN(new_n921));
  OAI21_X1  g720(.A(G190gat), .B1(new_n895), .B2(new_n286), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n898), .A2(new_n900), .ZN(new_n925));
  NOR4_X1   g724(.A1(new_n925), .A2(new_n545), .A3(new_n688), .A4(new_n772), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n395), .A3(new_n262), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n687), .A2(new_n894), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n880), .A2(new_n881), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n262), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n395), .ZN(G1352gat));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n396), .A3(new_n699), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n880), .A2(new_n699), .A3(new_n881), .A4(new_n928), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G204gat), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n926), .A2(new_n936), .A3(new_n396), .A4(new_n699), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(G1353gat));
  NAND4_X1  g737(.A1(new_n880), .A2(new_n698), .A3(new_n881), .A4(new_n928), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(G211gat), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n379), .A3(new_n698), .ZN(new_n946));
  INV_X1    g745(.A(new_n944), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n939), .A2(G211gat), .A3(new_n947), .A4(new_n942), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(G1354gat));
  AOI21_X1  g748(.A(G218gat), .B1(new_n926), .B2(new_n695), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n286), .A2(new_n380), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n929), .B2(new_n951), .ZN(G1355gat));
endmodule


