//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:34:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1232, new_n1233;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  INV_X1    g0007(.A(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G68), .A2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G244), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n215), .C1(G77), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n203), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(G58), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT64), .Z(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n206), .B(new_n227), .C1(new_n230), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n219), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n210), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(KEYINPUT66), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n209), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT67), .B(G45), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n254), .B(G274), .C1(new_n255), .C2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT68), .B(G226), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(new_n263), .B(KEYINPUT69), .Z(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  INV_X1    g0069(.A(G223), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n267), .B(new_n269), .C1(new_n270), .C2(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(new_n259), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n271), .B(new_n272), .C1(G77), .C2(new_n267), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G190), .ZN(new_n275));
  OR3_X1    g0075(.A1(new_n274), .A2(KEYINPUT72), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n232), .B2(G50), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n229), .A2(G33), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n228), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT70), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n229), .A2(G1), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n283), .A2(new_n286), .B1(new_n223), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n286), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n288), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n291), .B1(new_n223), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT9), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT72), .B1(new_n274), .B2(new_n275), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n274), .A2(G200), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n276), .A2(new_n295), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(new_n274), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n302), .B(new_n294), .C1(G169), .C2(new_n300), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n261), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G238), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  OAI211_X1 g0108(.A(G232), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT73), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n267), .A2(new_n311), .A3(G232), .A4(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT74), .ZN(new_n315));
  AOI21_X1  g0115(.A(G1698), .B1(new_n265), .B2(new_n266), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G226), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n313), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n256), .B(new_n306), .C1(new_n318), .C2(new_n259), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT75), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n310), .A2(new_n312), .B1(G226), .B2(new_n316), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n315), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n272), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(new_n256), .A4(new_n306), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n320), .A2(KEYINPUT13), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(G190), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT76), .ZN(new_n330));
  INV_X1    g0130(.A(G68), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT77), .B1(new_n290), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g0132(.A(new_n332), .B(KEYINPUT12), .Z(new_n333));
  NOR2_X1   g0133(.A1(new_n285), .A2(new_n287), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(G68), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n279), .A2(G50), .B1(G20), .B2(new_n331), .ZN(new_n336));
  INV_X1    g0136(.A(G77), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n281), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n286), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT11), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n319), .B(KEYINPUT13), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT76), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n326), .A2(new_n328), .A3(new_n344), .A4(G190), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n330), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G238), .A2(G1698), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n267), .B(new_n347), .C1(new_n219), .C2(G1698), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n272), .C1(G107), .C2(new_n267), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n305), .A2(new_n216), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n256), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n275), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G200), .B2(new_n351), .ZN(new_n353));
  INV_X1    g0153(.A(new_n282), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT15), .B(G87), .Z(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n281), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n285), .B1(G77), .B2(new_n334), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n290), .A2(new_n337), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n351), .A2(G179), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT71), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n362), .B1(new_n367), .B2(new_n351), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n363), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n326), .A2(G179), .A3(new_n328), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT78), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT78), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n326), .A2(new_n328), .A3(new_n374), .A4(G179), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n376));
  OAI21_X1  g0176(.A(G169), .B1(new_n376), .B2(new_n327), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n342), .A2(KEYINPUT14), .A3(G169), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n373), .A2(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n341), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n346), .B(new_n371), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT85), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT84), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT83), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n270), .A2(new_n268), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n224), .A2(G1698), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(new_n307), .C2(new_n308), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n389), .A2(KEYINPUT82), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT82), .B1(new_n389), .B2(new_n390), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n391), .A2(new_n392), .A3(new_n259), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n256), .B1(new_n261), .B2(new_n219), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n386), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n389), .A2(new_n390), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT82), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n389), .A2(KEYINPUT82), .A3(new_n390), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n272), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n394), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT83), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G200), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n400), .A2(new_n401), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G190), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(G58), .B(G68), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(G20), .B1(G159), .B2(new_n279), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n266), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n307), .A2(new_n308), .A3(G20), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT79), .B1(new_n414), .B2(KEYINPUT7), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT79), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n267), .C2(G20), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(KEYINPUT16), .B(new_n411), .C1(new_n419), .C2(new_n331), .ZN(new_n420));
  INV_X1    g0220(.A(new_n411), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT80), .B1(new_n414), .B2(KEYINPUT7), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT80), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n417), .C1(new_n267), .C2(G20), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n412), .A2(KEYINPUT81), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n307), .A2(new_n308), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT7), .A4(new_n229), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n422), .A2(new_n424), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n421), .B1(new_n429), .B2(G68), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n420), .B(new_n285), .C1(new_n430), .C2(KEYINPUT16), .ZN(new_n431));
  INV_X1    g0231(.A(new_n290), .ZN(new_n432));
  MUX2_X1   g0232(.A(new_n432), .B(new_n293), .S(new_n354), .Z(new_n433));
  AND2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n385), .B1(new_n409), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n433), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT84), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n384), .B(KEYINPUT17), .C1(new_n435), .C2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G169), .B1(new_n395), .B2(new_n402), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n406), .A2(G179), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n437), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n436), .A2(new_n437), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n385), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT84), .B1(new_n436), .B2(new_n437), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n446), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n439), .B(new_n445), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n304), .A2(new_n383), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n267), .A2(new_n229), .A3(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT22), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT22), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n267), .A2(new_n457), .A3(new_n229), .A4(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT24), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n207), .A2(G20), .ZN(new_n461));
  OAI22_X1  g0261(.A1(KEYINPUT23), .A2(new_n461), .B1(new_n281), .B2(new_n209), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(KEYINPUT23), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT92), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT92), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(new_n465), .A3(KEYINPUT23), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n459), .A2(new_n460), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n459), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n285), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n254), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n292), .A2(new_n432), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G107), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n290), .A2(new_n207), .ZN(new_n475));
  XOR2_X1   g0275(.A(new_n475), .B(KEYINPUT25), .Z(new_n476));
  NAND3_X1  g0276(.A1(new_n470), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n221), .A2(G1698), .ZN(new_n478));
  OAI221_X1 g0278(.A(new_n478), .B1(G250), .B2(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n479));
  INV_X1    g0279(.A(G294), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n257), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT88), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(G41), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n258), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n488), .A2(new_n259), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n481), .A2(new_n272), .B1(new_n489), .B2(G264), .ZN(new_n490));
  INV_X1    g0290(.A(G274), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G169), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n492), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n301), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n477), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT93), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n495), .A2(new_n404), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n494), .A2(new_n275), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n477), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G244), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G1698), .ZN(new_n505));
  OAI221_X1 g0305(.A(new_n505), .B1(G238), .B2(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G116), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n272), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n486), .A2(new_n491), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(new_n259), .C1(G250), .C2(new_n486), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n275), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(G200), .B2(new_n512), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n229), .B1(new_n315), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n213), .A2(new_n220), .A3(new_n207), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n267), .A2(new_n229), .A3(G68), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n515), .B1(new_n281), .B2(new_n220), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(new_n285), .B1(new_n290), .B2(new_n357), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n473), .A2(G87), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n514), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n512), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n301), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n512), .A2(new_n367), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n521), .A2(new_n285), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n357), .A2(new_n290), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n472), .A2(new_n357), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n526), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n488), .A2(new_n259), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n492), .B1(new_n221), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT89), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n426), .A2(new_n504), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(KEYINPUT4), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n267), .A2(G250), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n268), .B1(new_n541), .B2(KEYINPUT4), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n272), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT89), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n492), .B(new_n544), .C1(new_n221), .C2(new_n534), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n367), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(G179), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n285), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n429), .A2(KEYINPUT87), .A3(G107), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT87), .B1(new_n429), .B2(G107), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n220), .A2(new_n207), .A3(KEYINPUT6), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT86), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT6), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G97), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n554), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n207), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n560), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(G107), .A3(new_n558), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n550), .B1(new_n553), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n432), .A2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n472), .B2(new_n220), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n547), .B(new_n549), .C1(new_n566), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n429), .A2(G107), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n429), .A2(KEYINPUT87), .A3(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n565), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n569), .B1(new_n575), .B2(new_n285), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n546), .A2(G200), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n536), .A2(new_n543), .A3(new_n545), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT90), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n533), .A2(new_n570), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n538), .B(new_n229), .C1(G33), .C2(new_n220), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT91), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n284), .A2(new_n228), .B1(G20), .B2(new_n209), .ZN(new_n586));
  AOI21_X1  g0386(.A(G20), .B1(new_n257), .B2(G97), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(KEYINPUT91), .A3(new_n538), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n290), .A2(new_n209), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n432), .A2(G116), .A3(new_n550), .A4(new_n471), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n489), .A2(G270), .ZN(new_n595));
  INV_X1    g0395(.A(G303), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n259), .B1(new_n426), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n267), .B1(new_n208), .B2(new_n268), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n221), .A2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n492), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n594), .A2(G169), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT21), .ZN(new_n603));
  INV_X1    g0403(.A(new_n594), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n595), .A2(new_n600), .A3(G179), .A4(new_n492), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n601), .A2(G200), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n604), .B(new_n607), .C1(new_n275), .C2(new_n601), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n603), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n533), .A2(new_n570), .A3(new_n580), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(KEYINPUT90), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n454), .A2(new_n503), .A3(new_n582), .A4(new_n611), .ZN(G372));
  INV_X1    g0412(.A(new_n303), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n381), .A2(new_n382), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT95), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n366), .B2(new_n369), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT95), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n346), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n439), .B1(new_n450), .B2(new_n452), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n445), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n613), .B1(new_n621), .B2(new_n299), .ZN(new_n622));
  INV_X1    g0422(.A(new_n547), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n576), .A2(new_n623), .A3(new_n548), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n533), .A3(KEYINPUT26), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT26), .B1(new_n624), .B2(new_n533), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n532), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n502), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT94), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n497), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n603), .A2(new_n606), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(new_n610), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n454), .B1(new_n628), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n622), .A2(new_n635), .ZN(G369));
  NOR2_X1   g0436(.A1(new_n289), .A2(G20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n228), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT96), .ZN(new_n640));
  INV_X1    g0440(.A(G213), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n638), .B2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(KEYINPUT96), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n604), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n632), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n609), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n497), .B(KEYINPUT93), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n629), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n477), .A2(new_n646), .ZN(new_n655));
  OAI22_X1  g0455(.A1(new_n654), .A2(new_n655), .B1(new_n497), .B2(new_n647), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n646), .B1(new_n603), .B2(new_n606), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n503), .A2(new_n659), .B1(new_n631), .B2(new_n647), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n204), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n517), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n233), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(new_n532), .ZN(new_n669));
  INV_X1    g0469(.A(new_n627), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n625), .ZN(new_n671));
  INV_X1    g0471(.A(new_n610), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n672), .B(new_n629), .C1(new_n632), .C2(new_n631), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n646), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT29), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n672), .B(new_n629), .C1(new_n499), .C2(new_n632), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n646), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT29), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n601), .A2(new_n301), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n546), .A2(new_n680), .A3(new_n494), .A4(new_n512), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n481), .A2(new_n272), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n489), .A2(G264), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n509), .A4(new_n511), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT97), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n605), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n525), .A2(KEYINPUT97), .A3(new_n490), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n578), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT98), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT30), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT30), .B1(new_n688), .B2(new_n689), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n681), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT100), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT100), .B(new_n681), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n694), .A2(new_n646), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n611), .A2(new_n503), .A3(new_n582), .A4(new_n647), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(KEYINPUT31), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT99), .Z(new_n700));
  OAI21_X1  g0500(.A(G330), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n679), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n668), .B1(new_n703), .B2(G1), .ZN(G364));
  NOR2_X1   g0504(.A1(G13), .A2(G33), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G20), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n650), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n662), .A2(new_n267), .ZN(new_n710));
  OAI221_X1 g0510(.A(new_n710), .B1(new_n234), .B2(new_n255), .C1(new_n252), .C2(new_n485), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n662), .A2(new_n426), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(G355), .B(KEYINPUT101), .ZN(new_n714));
  OAI221_X1 g0514(.A(new_n711), .B1(G116), .B2(new_n204), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n228), .B1(G20), .B2(new_n367), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n637), .A2(G45), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n664), .A2(G1), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n229), .A2(new_n301), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(G190), .A3(G200), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT103), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n229), .A2(new_n301), .A3(G190), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n404), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT102), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n728), .A2(G50), .B1(G77), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n404), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G20), .A3(G190), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n213), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n426), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT105), .Z(new_n739));
  NAND3_X1  g0539(.A1(new_n722), .A2(G190), .A3(new_n404), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G58), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n229), .A2(G190), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT104), .B(KEYINPUT32), .Z(new_n748));
  XNOR2_X1  g0548(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n734), .A2(new_n739), .A3(new_n742), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n229), .B1(new_n744), .B2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n220), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n729), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n735), .A2(new_n743), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n331), .B1(new_n754), .B2(new_n207), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n750), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n736), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n733), .A2(G311), .B1(G303), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n745), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G329), .ZN(new_n760));
  INV_X1    g0560(.A(G317), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n753), .B1(KEYINPUT33), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(KEYINPUT33), .B2(new_n761), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n758), .A2(new_n426), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G326), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n727), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n740), .A2(new_n769), .B1(new_n751), .B2(new_n480), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n764), .A2(new_n766), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n716), .B1(new_n756), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n709), .A2(new_n718), .A3(new_n721), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n650), .A2(G330), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(new_n651), .A3(new_n720), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(G396));
  OAI211_X1 g0576(.A(new_n371), .B(new_n647), .C1(new_n634), .C2(new_n628), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n616), .A2(new_n361), .A3(new_n617), .A4(new_n646), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n370), .B1(new_n362), .B2(new_n647), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n777), .B1(new_n674), .B2(new_n781), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n701), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n701), .A2(new_n782), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(new_n720), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n716), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n728), .A2(G137), .B1(G143), .B2(new_n741), .ZN(new_n787));
  INV_X1    g0587(.A(new_n733), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n787), .B1(new_n278), .B2(new_n753), .C1(new_n746), .C2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT34), .Z(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G50), .B2(new_n757), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n426), .B1(new_n759), .B2(G132), .ZN(new_n792));
  INV_X1    g0592(.A(new_n751), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G58), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n754), .A2(new_n331), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n791), .A2(new_n792), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n754), .A2(new_n213), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n788), .A2(new_n209), .B1(new_n727), .B2(new_n596), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G294), .C2(new_n741), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n267), .B(new_n752), .C1(new_n804), .C2(G283), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n207), .B2(new_n736), .C1(new_n807), .C2(new_n745), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n786), .B1(new_n797), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n781), .A2(new_n706), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n809), .A2(new_n720), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n716), .A2(new_n705), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(G77), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n785), .A2(new_n814), .ZN(G384));
  INV_X1    g0615(.A(new_n644), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n419), .A2(new_n331), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n421), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n286), .B1(new_n818), .B2(KEYINPUT16), .ZN(new_n819));
  INV_X1    g0619(.A(new_n420), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n433), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n453), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n644), .B1(new_n440), .B2(new_n441), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT37), .B1(new_n823), .B2(new_n437), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n435), .B2(new_n438), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n448), .A2(new_n449), .B1(new_n823), .B2(new_n821), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT40), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n822), .A2(KEYINPUT38), .A3(new_n828), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n341), .A2(new_n646), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n346), .B(new_n835), .C1(new_n381), .C2(new_n382), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n381), .A2(new_n835), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n780), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n694), .A2(new_n646), .A3(new_n695), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT31), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n698), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT109), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT40), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n834), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n825), .A2(KEYINPUT107), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n823), .A2(new_n437), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT37), .B1(new_n848), .B2(new_n447), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT107), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n824), .C1(new_n435), .C2(new_n438), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT108), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n453), .A2(new_n437), .A3(new_n816), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT108), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n847), .A2(new_n855), .A3(new_n849), .A4(new_n851), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n830), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n833), .A2(new_n858), .B1(new_n842), .B2(new_n844), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n846), .B1(new_n859), .B2(new_n832), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n454), .B1(new_n698), .B2(new_n841), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(G330), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n822), .A2(KEYINPUT38), .A3(new_n828), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n822), .B2(new_n828), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n366), .A2(new_n369), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n647), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n777), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n836), .A2(new_n837), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n866), .A2(new_n871), .B1(new_n445), .B2(new_n816), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT39), .B1(new_n858), .B2(new_n833), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n864), .A2(new_n865), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n614), .A2(new_n647), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n872), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n675), .A2(new_n678), .A3(new_n454), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n622), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n879), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n863), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n254), .B2(new_n637), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n209), .B1(new_n564), .B2(KEYINPUT35), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n230), .C1(KEYINPUT35), .C2(new_n564), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT36), .ZN(new_n887));
  OAI21_X1  g0687(.A(G77), .B1(new_n218), .B2(new_n331), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n233), .A2(new_n888), .B1(G50), .B2(new_n331), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(G1), .A3(new_n289), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(new_n887), .A3(new_n890), .ZN(G367));
  NAND2_X1  g0691(.A1(new_n728), .A2(G311), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n736), .A2(new_n209), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n267), .B1(new_n893), .B2(KEYINPUT46), .ZN(new_n894));
  INV_X1    g0694(.A(new_n754), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(G97), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n733), .A2(G283), .B1(G107), .B2(new_n793), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n892), .A2(new_n894), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n803), .A2(new_n480), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n893), .A2(KEYINPUT46), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n740), .A2(new_n596), .B1(new_n745), .B2(new_n761), .ZN(new_n901));
  NOR4_X1   g0701(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n267), .B1(new_n331), .B2(new_n751), .C1(new_n788), .C2(new_n223), .ZN(new_n903));
  AOI22_X1  g0703(.A1(G143), .A2(new_n728), .B1(new_n804), .B2(G159), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n904), .B1(new_n337), .B2(new_n754), .C1(new_n278), .C2(new_n740), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n903), .B(new_n905), .C1(G137), .C2(new_n759), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n757), .A2(G58), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT47), .Z(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n716), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n522), .A2(new_n523), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n646), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n532), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n533), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n707), .ZN(new_n915));
  INV_X1    g0715(.A(new_n710), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n717), .B1(new_n204), .B2(new_n357), .C1(new_n243), .C2(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n910), .A2(new_n721), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n570), .B(new_n580), .C1(new_n576), .C2(new_n647), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n570), .B2(new_n647), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n657), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT43), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT110), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n921), .B(new_n924), .Z(new_n925));
  NOR2_X1   g0725(.A1(new_n914), .A2(new_n922), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n656), .A2(new_n659), .A3(new_n920), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT42), .Z(new_n928));
  OAI21_X1  g0728(.A(new_n570), .B1(new_n919), .B2(new_n653), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n647), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n925), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n719), .A2(G1), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n660), .A2(new_n920), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT45), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n660), .A2(new_n920), .A3(KEYINPUT44), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT44), .B1(new_n660), .B2(new_n920), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n503), .A2(new_n659), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n656), .B2(new_n659), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n657), .B1(new_n651), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n703), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n663), .B(KEYINPUT41), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n918), .B1(new_n932), .B2(new_n946), .ZN(G387));
  NAND2_X1  g0747(.A1(new_n703), .A2(new_n942), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n664), .B1(new_n702), .B2(new_n943), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n942), .A2(new_n933), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n426), .B1(new_n745), .B2(new_n765), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n733), .A2(G303), .B1(G317), .B2(new_n741), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n807), .B2(new_n803), .C1(new_n769), .C2(new_n727), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT48), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n767), .B2(new_n751), .C1(new_n480), .C2(new_n736), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT49), .Z(new_n957));
  AOI211_X1 g0757(.A(new_n952), .B(new_n957), .C1(G116), .C2(new_n895), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n736), .A2(new_n337), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G50), .B2(new_n741), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n960), .B(new_n267), .C1(new_n278), .C2(new_n745), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n733), .A2(G68), .ZN(new_n962));
  INV_X1    g0762(.A(new_n753), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n354), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n793), .A2(new_n356), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n962), .A2(new_n896), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n961), .B(new_n966), .C1(G159), .C2(new_n728), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n716), .B1(new_n958), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n916), .B1(new_n240), .B2(new_n255), .ZN(new_n969));
  INV_X1    g0769(.A(new_n665), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n970), .B2(new_n712), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n282), .A2(KEYINPUT50), .A3(G50), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT50), .B1(new_n282), .B2(G50), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n485), .A4(new_n665), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G68), .B2(G77), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n971), .A2(new_n975), .B1(G107), .B2(new_n204), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n720), .B1(new_n976), .B2(new_n717), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n968), .B(new_n977), .C1(new_n656), .C2(new_n708), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n950), .A2(new_n951), .A3(new_n978), .ZN(G393));
  NAND2_X1  g0779(.A1(new_n939), .A2(new_n658), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n657), .B1(new_n935), .B2(new_n938), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n948), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n983), .B(new_n663), .C1(new_n948), .C2(new_n939), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n933), .A3(new_n981), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n895), .A2(G107), .B1(new_n759), .B2(G322), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n426), .B(new_n986), .C1(new_n788), .C2(new_n480), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n728), .A2(G317), .B1(G311), .B2(new_n741), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n988), .A2(new_n990), .B1(new_n767), .B2(new_n736), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n987), .B(new_n991), .C1(new_n988), .C2(new_n990), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n209), .B2(new_n751), .C1(new_n596), .C2(new_n803), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n727), .A2(new_n278), .B1(new_n746), .B2(new_n740), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT51), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n426), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n733), .A2(new_n354), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n804), .A2(G50), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n736), .A2(new_n331), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n798), .B(new_n999), .C1(G143), .C2(new_n759), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n751), .A2(new_n337), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n716), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n717), .B1(new_n220), .B2(new_n204), .C1(new_n248), .C2(new_n916), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n920), .A2(new_n708), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n721), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n984), .A2(new_n985), .A3(new_n1007), .ZN(G390));
  INV_X1    g0808(.A(KEYINPUT112), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n781), .A2(G330), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n870), .C1(new_n698), .C2(new_n841), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n871), .A2(new_n877), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n873), .B2(new_n875), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n858), .A2(new_n833), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n836), .A2(new_n837), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n677), .A2(new_n781), .B1(new_n867), .B2(new_n647), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n877), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1009), .B(new_n1011), .C1(new_n1013), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1011), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1010), .B(new_n870), .C1(new_n698), .C2(new_n700), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1013), .A2(new_n1017), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT112), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1018), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1010), .B1(new_n698), .B2(new_n700), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n1015), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n1011), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n869), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1010), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n697), .A2(KEYINPUT31), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n841), .B1(new_n1030), .B2(new_n839), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1015), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n1016), .A3(new_n1021), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n454), .B(G330), .C1(new_n698), .C2(new_n841), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n880), .A2(new_n1035), .A3(new_n622), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT113), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1024), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1024), .A2(new_n1039), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n663), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n426), .B1(new_n745), .B2(new_n480), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n737), .B(new_n1043), .C1(new_n728), .C2(G283), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n741), .A2(G116), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n804), .A2(G107), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n795), .B(new_n1002), .C1(new_n733), .C2(G97), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(G132), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n740), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(G128), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n727), .A2(new_n1051), .B1(new_n746), .B2(new_n751), .ZN(new_n1052));
  INV_X1    g0852(.A(G125), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n267), .B1(new_n745), .B2(new_n1053), .C1(new_n223), .C2(new_n754), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1050), .B(new_n1052), .C1(KEYINPUT115), .C2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT54), .B(G143), .Z(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(G137), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n788), .A2(new_n1057), .B1(new_n803), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT114), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1055), .B(new_n1060), .C1(KEYINPUT115), .C2(new_n1054), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n736), .A2(new_n278), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1048), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n716), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n721), .B(new_n1066), .C1(new_n876), .C2(new_n706), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n282), .B2(new_n812), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1024), .B2(new_n933), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1042), .A2(new_n1069), .ZN(G378));
  NOR2_X1   g0870(.A1(new_n751), .A2(new_n278), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1057), .A2(new_n736), .B1(new_n753), .B2(new_n1049), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n733), .C2(G137), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n1053), .B2(new_n727), .C1(new_n1051), .C2(new_n740), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT59), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n895), .A2(G159), .ZN(new_n1076));
  AOI21_X1  g0876(.A(G41), .B1(new_n759), .B2(G124), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1075), .A2(new_n257), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(KEYINPUT59), .B2(new_n1074), .ZN(new_n1079));
  AOI21_X1  g0879(.A(G50), .B1(new_n266), .B2(new_n258), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n895), .A2(G58), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n207), .B2(new_n740), .C1(new_n788), .C2(new_n357), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n959), .B(new_n1083), .C1(G97), .C2(new_n963), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n258), .B1(new_n751), .B2(new_n331), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n267), .B(new_n1085), .C1(G283), .C2(new_n759), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(new_n209), .C2(new_n727), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n786), .B1(new_n1081), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n720), .B1(new_n223), .B2(new_n812), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n294), .A2(new_n816), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n304), .B(new_n1095), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1094), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1093), .A3(new_n1099), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1090), .B(new_n1092), .C1(new_n1105), .C2(new_n705), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n834), .A2(new_n843), .A3(new_n845), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n842), .A2(new_n844), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n832), .B1(new_n1014), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(G330), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n879), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1105), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n873), .A2(new_n875), .A3(new_n877), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n860), .B(G330), .C1(new_n1113), .C2(new_n872), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1106), .B1(new_n1117), .B2(new_n933), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1105), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1111), .A2(new_n1114), .A3(new_n1112), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(KEYINPUT57), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1036), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n663), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1019), .A2(KEYINPUT112), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1022), .A2(KEYINPUT112), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1034), .C1(new_n1126), .C2(new_n1019), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1037), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT57), .B1(new_n1128), .B2(new_n1117), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1118), .B1(new_n1124), .B2(new_n1129), .ZN(G375));
  NAND3_X1  g0930(.A1(new_n1028), .A2(new_n1036), .A3(new_n1033), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1038), .A2(new_n945), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT121), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1082), .A2(new_n1133), .A3(new_n267), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n803), .B2(new_n1057), .C1(new_n788), .C2(new_n278), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n1082), .B2(new_n267), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n727), .A2(new_n1049), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n740), .A2(new_n1058), .B1(new_n736), .B2(new_n746), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n223), .B2(new_n751), .C1(new_n1051), .C2(new_n745), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n727), .A2(new_n480), .B1(new_n337), .B2(new_n754), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n426), .B1(new_n788), .B2(new_n207), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n965), .B1(new_n803), .B2(new_n209), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n745), .A2(new_n596), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n220), .B2(new_n736), .C1(new_n767), .C2(new_n740), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n786), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n720), .B(new_n1147), .C1(new_n331), .C2(new_n812), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1015), .A2(new_n705), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT120), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1034), .A2(new_n933), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1132), .A2(new_n1151), .ZN(G381));
  INV_X1    g0952(.A(new_n1106), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n933), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1115), .A2(new_n1116), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n664), .B1(new_n1158), .B2(new_n1128), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1123), .B2(new_n1154), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1042), .A2(new_n1069), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1163), .A2(G384), .A3(G381), .ZN(new_n1164));
  OR2_X1    g0964(.A1(G393), .A2(G396), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(G390), .A2(new_n1165), .A3(G387), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(G407));
  OAI211_X1 g0967(.A(G407), .B(G213), .C1(G343), .C2(new_n1163), .ZN(G409));
  XNOR2_X1  g0968(.A(G393), .B(G396), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT123), .ZN(new_n1170));
  AND2_X1   g0970(.A1(G390), .A2(G387), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(G390), .A2(G387), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(KEYINPUT124), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1170), .A2(new_n1173), .B1(new_n1176), .B2(KEYINPUT124), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT126), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(KEYINPUT126), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT61), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n641), .A2(G343), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1128), .A2(new_n1117), .A3(new_n945), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1042), .A2(new_n1118), .A3(new_n1184), .A4(new_n1069), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT60), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1131), .A2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1028), .A2(new_n1036), .A3(KEYINPUT60), .A4(new_n1033), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1188), .A2(new_n1038), .A3(new_n663), .A4(new_n1189), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1190), .A2(G384), .A3(new_n1151), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G384), .B1(new_n1190), .B2(new_n1151), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1186), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT62), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1181), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT122), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1190), .A2(new_n1151), .ZN(new_n1199));
  INV_X1    g0999(.A(G384), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT122), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1190), .A2(G384), .A3(new_n1151), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1182), .A2(G2897), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1198), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1193), .A2(new_n1202), .A3(G2897), .A4(new_n1182), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1186), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1210), .A2(new_n1193), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT62), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1179), .B(new_n1180), .C1(new_n1197), .C2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT63), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1214), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1216), .A2(new_n1217), .A3(KEYINPUT125), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT125), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1182), .B1(G375), .B2(G378), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n1185), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT63), .B1(new_n1195), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1181), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1214), .B2(new_n1211), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1219), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1213), .B1(new_n1218), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT127), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n1213), .C1(new_n1218), .C2(new_n1226), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(G405));
  NAND2_X1  g1031(.A1(new_n1163), .A2(new_n1210), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(new_n1193), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(new_n1178), .ZN(G402));
endmodule


