

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715;

  XOR2_X2 U366 ( .A(n582), .B(KEYINPUT38), .Z(n627) );
  INV_X2 U367 ( .A(G953), .ZN(n704) );
  XNOR2_X1 U368 ( .A(n367), .B(n576), .ZN(n366) );
  XNOR2_X1 U369 ( .A(n504), .B(n503), .ZN(n513) );
  XNOR2_X1 U370 ( .A(n465), .B(KEYINPUT22), .ZN(n527) );
  NOR2_X1 U371 ( .A1(n510), .A2(n524), .ZN(n357) );
  XNOR2_X1 U372 ( .A(n590), .B(n585), .ZN(n701) );
  NAND2_X1 U373 ( .A1(n366), .A2(n584), .ZN(n590) );
  XNOR2_X1 U374 ( .A(n398), .B(KEYINPUT74), .ZN(n397) );
  XNOR2_X1 U375 ( .A(n387), .B(n386), .ZN(n712) );
  AND2_X1 U376 ( .A1(n512), .A2(n511), .ZN(n387) );
  NOR2_X1 U377 ( .A1(n527), .A2(n498), .ZN(n500) );
  XNOR2_X1 U378 ( .A(n438), .B(KEYINPUT0), .ZN(n521) );
  INV_X1 U379 ( .A(n518), .ZN(n647) );
  BUF_X1 U380 ( .A(n536), .Z(n582) );
  XNOR2_X1 U381 ( .A(n476), .B(G472), .ZN(n518) );
  XNOR2_X1 U382 ( .A(n434), .B(n433), .ZN(n536) );
  XNOR2_X1 U383 ( .A(n450), .B(n449), .ZN(n524) );
  XNOR2_X1 U384 ( .A(n355), .B(n457), .ZN(n683) );
  XNOR2_X1 U385 ( .A(n454), .B(n392), .ZN(n430) );
  XNOR2_X1 U386 ( .A(n364), .B(KEYINPUT75), .ZN(n445) );
  XNOR2_X1 U387 ( .A(n406), .B(n345), .ZN(n426) );
  XNOR2_X1 U388 ( .A(n369), .B(G104), .ZN(n443) );
  XNOR2_X1 U389 ( .A(n442), .B(n441), .ZN(n481) );
  XNOR2_X1 U390 ( .A(n391), .B(G131), .ZN(n444) );
  XNOR2_X1 U391 ( .A(G101), .B(G104), .ZN(n466) );
  XOR2_X1 U392 ( .A(G146), .B(G125), .Z(n442) );
  XNOR2_X1 U393 ( .A(n700), .B(G146), .ZN(n473) );
  XNOR2_X1 U394 ( .A(n430), .B(n388), .ZN(n700) );
  XNOR2_X1 U395 ( .A(n444), .B(n389), .ZN(n388) );
  XNOR2_X1 U396 ( .A(n390), .B(KEYINPUT71), .ZN(n389) );
  INV_X1 U397 ( .A(G134), .ZN(n390) );
  INV_X1 U398 ( .A(n525), .ZN(n510) );
  XNOR2_X1 U399 ( .A(n357), .B(KEYINPUT105), .ZN(n630) );
  XNOR2_X1 U400 ( .A(n376), .B(n375), .ZN(n681) );
  XNOR2_X1 U401 ( .A(n348), .B(n481), .ZN(n375) );
  XNOR2_X1 U402 ( .A(n446), .B(n377), .ZN(n376) );
  NOR2_X1 U403 ( .A1(n701), .A2(n586), .ZN(n373) );
  XNOR2_X1 U404 ( .A(n403), .B(n402), .ZN(n401) );
  XNOR2_X1 U405 ( .A(n442), .B(n347), .ZN(n402) );
  XNOR2_X1 U406 ( .A(n429), .B(n430), .ZN(n403) );
  XNOR2_X1 U407 ( .A(n383), .B(n349), .ZN(n382) );
  NAND2_X1 U408 ( .A1(n685), .A2(G472), .ZN(n383) );
  NAND2_X1 U409 ( .A1(n685), .A2(G475), .ZN(n371) );
  NAND2_X1 U410 ( .A1(n385), .A2(n384), .ZN(n398) );
  NOR2_X1 U411 ( .A1(n513), .A2(KEYINPUT44), .ZN(n384) );
  INV_X1 U412 ( .A(n712), .ZN(n385) );
  NOR2_X1 U413 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U414 ( .A1(n515), .A2(n533), .ZN(n394) );
  XNOR2_X1 U415 ( .A(n514), .B(n396), .ZN(n395) );
  AND2_X1 U416 ( .A1(n575), .A2(n623), .ZN(n368) );
  XNOR2_X1 U417 ( .A(n419), .B(n407), .ZN(n420) );
  XNOR2_X1 U418 ( .A(G134), .B(G122), .ZN(n451) );
  NAND2_X1 U419 ( .A1(n413), .A2(n412), .ZN(n454) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n577) );
  INV_X1 U421 ( .A(KEYINPUT39), .ZN(n360) );
  NOR2_X1 U422 ( .A1(n553), .A2(n363), .ZN(n362) );
  XOR2_X1 U423 ( .A(n460), .B(n459), .Z(n525) );
  NOR2_X1 U424 ( .A1(n683), .A2(G902), .ZN(n460) );
  NOR2_X1 U425 ( .A1(n681), .A2(G902), .ZN(n450) );
  XNOR2_X1 U426 ( .A(n426), .B(n404), .ZN(n694) );
  AND2_X2 U427 ( .A1(n671), .A2(n592), .ZN(n685) );
  XOR2_X1 U428 ( .A(G107), .B(G110), .Z(n470) );
  INV_X1 U429 ( .A(KEYINPUT66), .ZN(n396) );
  INV_X1 U430 ( .A(KEYINPUT70), .ZN(n391) );
  NAND2_X1 U431 ( .A1(G234), .A2(G237), .ZN(n421) );
  XNOR2_X1 U432 ( .A(G137), .B(G116), .ZN(n416) );
  NAND2_X1 U433 ( .A1(n704), .A2(n365), .ZN(n364) );
  INV_X1 U434 ( .A(G237), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n447), .B(n408), .ZN(n377) );
  XOR2_X1 U436 ( .A(KEYINPUT11), .B(G140), .Z(n408) );
  XNOR2_X1 U437 ( .A(G113), .B(G143), .ZN(n439) );
  XNOR2_X1 U438 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n441) );
  XNOR2_X1 U439 ( .A(G137), .B(G140), .ZN(n479) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n392) );
  XNOR2_X1 U441 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U442 ( .A(n415), .B(n414), .ZN(n406) );
  XOR2_X1 U443 ( .A(KEYINPUT3), .B(KEYINPUT91), .Z(n415) );
  INV_X1 U444 ( .A(G122), .ZN(n369) );
  XNOR2_X1 U445 ( .A(KEYINPUT96), .B(KEYINPUT23), .ZN(n484) );
  XNOR2_X1 U446 ( .A(G119), .B(G128), .ZN(n482) );
  INV_X1 U447 ( .A(KEYINPUT85), .ZN(n585) );
  NOR2_X1 U448 ( .A1(n640), .A2(n378), .ZN(n497) );
  XNOR2_X1 U449 ( .A(n542), .B(n379), .ZN(n378) );
  INV_X1 U450 ( .A(KEYINPUT79), .ZN(n379) );
  XNOR2_X1 U451 ( .A(n518), .B(KEYINPUT6), .ZN(n542) );
  NAND2_X1 U452 ( .A1(n356), .A2(n508), .ZN(n465) );
  NOR2_X1 U453 ( .A1(n630), .A2(n505), .ZN(n464) );
  XNOR2_X1 U454 ( .A(n456), .B(n458), .ZN(n355) );
  XNOR2_X1 U455 ( .A(n400), .B(n344), .ZN(n399) );
  NOR2_X1 U456 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U457 ( .A1(n577), .A2(n615), .ZN(n554) );
  INV_X1 U458 ( .A(KEYINPUT35), .ZN(n386) );
  NAND2_X1 U459 ( .A1(n382), .A2(n381), .ZN(n380) );
  XNOR2_X1 U460 ( .A(n371), .B(n350), .ZN(n370) );
  XNOR2_X1 U461 ( .A(n677), .B(n358), .ZN(n680) );
  XNOR2_X1 U462 ( .A(n679), .B(n678), .ZN(n358) );
  XNOR2_X1 U463 ( .A(n594), .B(n597), .ZN(n344) );
  XNOR2_X1 U464 ( .A(G101), .B(KEYINPUT73), .ZN(n345) );
  XNOR2_X1 U465 ( .A(KEYINPUT16), .B(G110), .ZN(n346) );
  AND2_X1 U466 ( .A1(G224), .A2(n704), .ZN(n347) );
  AND2_X1 U467 ( .A1(G214), .A2(n445), .ZN(n348) );
  XOR2_X1 U468 ( .A(n475), .B(KEYINPUT62), .Z(n349) );
  XOR2_X1 U469 ( .A(n681), .B(n409), .Z(n350) );
  XNOR2_X1 U470 ( .A(n694), .B(n401), .ZN(n594) );
  NOR2_X1 U471 ( .A1(G952), .A2(n704), .ZN(n689) );
  INV_X1 U472 ( .A(n689), .ZN(n381) );
  XOR2_X1 U473 ( .A(n593), .B(KEYINPUT90), .Z(n351) );
  XOR2_X1 U474 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n352) );
  XOR2_X1 U475 ( .A(n599), .B(n598), .Z(n353) );
  XNOR2_X1 U476 ( .A(n354), .B(n352), .ZN(G60) );
  NAND2_X1 U477 ( .A1(n370), .A2(n381), .ZN(n354) );
  XNOR2_X1 U478 ( .A(n464), .B(KEYINPUT106), .ZN(n356) );
  XNOR2_X1 U479 ( .A(n359), .B(n353), .ZN(G51) );
  NAND2_X1 U480 ( .A1(n399), .A2(n381), .ZN(n359) );
  NAND2_X1 U481 ( .A1(n552), .A2(n551), .ZN(n571) );
  NAND2_X1 U482 ( .A1(n552), .A2(n362), .ZN(n361) );
  INV_X1 U483 ( .A(n551), .ZN(n363) );
  NAND2_X1 U484 ( .A1(n564), .A2(n368), .ZN(n367) );
  NAND2_X1 U485 ( .A1(n372), .A2(n588), .ZN(n592) );
  NAND2_X1 U486 ( .A1(n374), .A2(n373), .ZN(n372) );
  INV_X1 U487 ( .A(n667), .ZN(n374) );
  XNOR2_X1 U488 ( .A(n535), .B(n534), .ZN(n667) );
  XNOR2_X1 U489 ( .A(n500), .B(n499), .ZN(n713) );
  XNOR2_X1 U490 ( .A(n380), .B(n351), .ZN(G57) );
  NAND2_X1 U491 ( .A1(n397), .A2(n393), .ZN(n535) );
  NAND2_X1 U492 ( .A1(n685), .A2(G210), .ZN(n400) );
  XNOR2_X1 U493 ( .A(n405), .B(n346), .ZN(n404) );
  XNOR2_X1 U494 ( .A(n453), .B(n443), .ZN(n405) );
  NAND2_X1 U495 ( .A1(n513), .A2(KEYINPUT44), .ZN(n514) );
  XOR2_X1 U496 ( .A(n418), .B(n417), .Z(n407) );
  XNOR2_X1 U497 ( .A(KEYINPUT59), .B(KEYINPUT67), .ZN(n409) );
  XNOR2_X1 U498 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n642) );
  XNOR2_X1 U499 ( .A(n643), .B(n642), .ZN(n644) );
  INV_X1 U500 ( .A(KEYINPUT87), .ZN(n503) );
  XNOR2_X1 U501 ( .A(KEYINPUT52), .B(KEYINPUT120), .ZN(n655) );
  XNOR2_X1 U502 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U503 ( .A(n466), .B(KEYINPUT95), .ZN(n467) );
  XNOR2_X1 U504 ( .A(n467), .B(n479), .ZN(n469) );
  XNOR2_X1 U505 ( .A(n473), .B(n420), .ZN(n475) );
  XNOR2_X1 U506 ( .A(n448), .B(G475), .ZN(n449) );
  INV_X1 U507 ( .A(KEYINPUT63), .ZN(n593) );
  INV_X1 U508 ( .A(KEYINPUT32), .ZN(n499) );
  INV_X1 U509 ( .A(G128), .ZN(n410) );
  NAND2_X1 U510 ( .A1(G143), .A2(n410), .ZN(n413) );
  INV_X1 U511 ( .A(G143), .ZN(n411) );
  NAND2_X1 U512 ( .A1(n411), .A2(G128), .ZN(n412) );
  XNOR2_X1 U513 ( .A(G119), .B(G113), .ZN(n414) );
  INV_X1 U514 ( .A(n426), .ZN(n419) );
  NAND2_X1 U515 ( .A1(n445), .A2(G210), .ZN(n418) );
  XNOR2_X1 U516 ( .A(n416), .B(KEYINPUT5), .ZN(n417) );
  NOR2_X1 U517 ( .A1(G898), .A2(n704), .ZN(n696) );
  XNOR2_X1 U518 ( .A(KEYINPUT14), .B(n421), .ZN(n423) );
  NAND2_X1 U519 ( .A1(G902), .A2(n423), .ZN(n537) );
  INV_X1 U520 ( .A(n537), .ZN(n422) );
  NAND2_X1 U521 ( .A1(n696), .A2(n422), .ZN(n425) );
  NAND2_X1 U522 ( .A1(G952), .A2(n423), .ZN(n658) );
  NOR2_X1 U523 ( .A1(n658), .A2(G953), .ZN(n424) );
  XNOR2_X1 U524 ( .A(n424), .B(KEYINPUT93), .ZN(n540) );
  NAND2_X1 U525 ( .A1(n425), .A2(n540), .ZN(n437) );
  XOR2_X1 U526 ( .A(G116), .B(G107), .Z(n453) );
  XOR2_X1 U527 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n428) );
  XNOR2_X1 U528 ( .A(KEYINPUT89), .B(KEYINPUT78), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U530 ( .A(G902), .B(KEYINPUT15), .ZN(n586) );
  NAND2_X1 U531 ( .A1(n594), .A2(n586), .ZN(n434) );
  OR2_X1 U532 ( .A1(G237), .A2(G902), .ZN(n435) );
  NAND2_X1 U533 ( .A1(G210), .A2(n435), .ZN(n432) );
  INV_X1 U534 ( .A(KEYINPUT92), .ZN(n431) );
  NAND2_X1 U535 ( .A1(G214), .A2(n435), .ZN(n628) );
  NAND2_X1 U536 ( .A1(n536), .A2(n628), .ZN(n436) );
  XNOR2_X1 U537 ( .A(n436), .B(KEYINPUT19), .ZN(n566) );
  NAND2_X1 U538 ( .A1(n437), .A2(n566), .ZN(n438) );
  INV_X1 U539 ( .A(n521), .ZN(n508) );
  XOR2_X1 U540 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n440) );
  XNOR2_X1 U541 ( .A(n440), .B(n439), .ZN(n447) );
  XOR2_X1 U542 ( .A(n444), .B(n443), .Z(n446) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n448) );
  XOR2_X1 U544 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n452) );
  XNOR2_X1 U545 ( .A(n452), .B(n451), .ZN(n458) );
  XOR2_X1 U546 ( .A(n454), .B(n453), .Z(n457) );
  NAND2_X1 U547 ( .A1(G234), .A2(n704), .ZN(n455) );
  XOR2_X1 U548 ( .A(KEYINPUT8), .B(n455), .Z(n488) );
  NAND2_X1 U549 ( .A1(G217), .A2(n488), .ZN(n456) );
  XNOR2_X1 U550 ( .A(KEYINPUT103), .B(G478), .ZN(n459) );
  NAND2_X1 U551 ( .A1(n586), .A2(G234), .ZN(n462) );
  XNOR2_X1 U552 ( .A(KEYINPUT20), .B(KEYINPUT98), .ZN(n461) );
  XNOR2_X1 U553 ( .A(n462), .B(n461), .ZN(n492) );
  NAND2_X1 U554 ( .A1(n492), .A2(G221), .ZN(n463) );
  XOR2_X1 U555 ( .A(n463), .B(KEYINPUT21), .Z(n636) );
  XOR2_X1 U556 ( .A(n636), .B(KEYINPUT100), .Z(n505) );
  NAND2_X1 U557 ( .A1(G227), .A2(n704), .ZN(n468) );
  XNOR2_X1 U558 ( .A(n469), .B(n468), .ZN(n471) );
  XNOR2_X1 U559 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U560 ( .A(n473), .B(n472), .ZN(n679) );
  NOR2_X1 U561 ( .A1(n679), .A2(G902), .ZN(n474) );
  XOR2_X1 U562 ( .A(n474), .B(G469), .Z(n558) );
  XOR2_X1 U563 ( .A(KEYINPUT1), .B(n558), .Z(n640) );
  INV_X1 U564 ( .A(n640), .ZN(n579) );
  NOR2_X1 U565 ( .A1(n475), .A2(G902), .ZN(n476) );
  XOR2_X1 U566 ( .A(KEYINPUT76), .B(KEYINPUT25), .Z(n478) );
  XNOR2_X1 U567 ( .A(KEYINPUT99), .B(KEYINPUT97), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n478), .B(n477), .ZN(n496) );
  INV_X1 U569 ( .A(n479), .ZN(n480) );
  XOR2_X1 U570 ( .A(n481), .B(n480), .Z(n699) );
  XOR2_X1 U571 ( .A(KEYINPUT24), .B(G110), .Z(n483) );
  XNOR2_X1 U572 ( .A(n483), .B(n482), .ZN(n487) );
  XOR2_X1 U573 ( .A(KEYINPUT82), .B(KEYINPUT77), .Z(n485) );
  XNOR2_X1 U574 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U575 ( .A(n487), .B(n486), .Z(n490) );
  NAND2_X1 U576 ( .A1(G221), .A2(n488), .ZN(n489) );
  XNOR2_X1 U577 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U578 ( .A(n699), .B(n491), .ZN(n687) );
  NOR2_X1 U579 ( .A1(G902), .A2(n687), .ZN(n494) );
  NAND2_X1 U580 ( .A1(G217), .A2(n492), .ZN(n493) );
  XNOR2_X1 U581 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U582 ( .A(n496), .B(n495), .ZN(n528) );
  INV_X1 U583 ( .A(n528), .ZN(n637) );
  NAND2_X1 U584 ( .A1(n497), .A2(n528), .ZN(n498) );
  NOR2_X1 U585 ( .A1(n637), .A2(n527), .ZN(n502) );
  NOR2_X1 U586 ( .A1(n647), .A2(n579), .ZN(n501) );
  NAND2_X1 U587 ( .A1(n502), .A2(n501), .ZN(n607) );
  NAND2_X1 U588 ( .A1(n713), .A2(n607), .ZN(n504) );
  XOR2_X1 U589 ( .A(KEYINPUT108), .B(KEYINPUT33), .Z(n507) );
  NOR2_X1 U590 ( .A1(n528), .A2(n505), .ZN(n516) );
  INV_X1 U591 ( .A(n516), .ZN(n641) );
  NOR2_X1 U592 ( .A1(n640), .A2(n641), .ZN(n520) );
  NAND2_X1 U593 ( .A1(n520), .A2(n542), .ZN(n506) );
  XNOR2_X1 U594 ( .A(n507), .B(n506), .ZN(n660) );
  XOR2_X1 U595 ( .A(n508), .B(KEYINPUT94), .Z(n517) );
  NOR2_X1 U596 ( .A1(n660), .A2(n517), .ZN(n509) );
  XNOR2_X1 U597 ( .A(KEYINPUT34), .B(n509), .ZN(n512) );
  NAND2_X1 U598 ( .A1(n524), .A2(n510), .ZN(n570) );
  INV_X1 U599 ( .A(n570), .ZN(n511) );
  NAND2_X1 U600 ( .A1(n712), .A2(KEYINPUT44), .ZN(n515) );
  NAND2_X1 U601 ( .A1(n558), .A2(n516), .ZN(n550) );
  NOR2_X1 U602 ( .A1(n550), .A2(n517), .ZN(n519) );
  NAND2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n602) );
  NAND2_X1 U604 ( .A1(n647), .A2(n520), .ZN(n649) );
  NOR2_X1 U605 ( .A1(n649), .A2(n521), .ZN(n522) );
  XNOR2_X1 U606 ( .A(n522), .B(KEYINPUT31), .ZN(n618) );
  NAND2_X1 U607 ( .A1(n602), .A2(n618), .ZN(n526) );
  NAND2_X1 U608 ( .A1(n524), .A2(n525), .ZN(n523) );
  XNOR2_X1 U609 ( .A(n523), .B(KEYINPUT104), .ZN(n615) );
  OR2_X1 U610 ( .A1(n525), .A2(n524), .ZN(n619) );
  NAND2_X1 U611 ( .A1(n615), .A2(n619), .ZN(n568) );
  NAND2_X1 U612 ( .A1(n526), .A2(n568), .ZN(n531) );
  NOR2_X1 U613 ( .A1(n527), .A2(n579), .ZN(n530) );
  NOR2_X1 U614 ( .A1(n542), .A2(n528), .ZN(n529) );
  NAND2_X1 U615 ( .A1(n530), .A2(n529), .ZN(n600) );
  NAND2_X1 U616 ( .A1(n531), .A2(n600), .ZN(n532) );
  XNOR2_X1 U617 ( .A(KEYINPUT107), .B(n532), .ZN(n533) );
  XOR2_X1 U618 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n534) );
  INV_X1 U619 ( .A(n582), .ZN(n545) );
  NOR2_X1 U620 ( .A1(G900), .A2(n537), .ZN(n538) );
  NAND2_X1 U621 ( .A1(G953), .A2(n538), .ZN(n539) );
  NAND2_X1 U622 ( .A1(n540), .A2(n539), .ZN(n551) );
  NAND2_X1 U623 ( .A1(n551), .A2(n636), .ZN(n541) );
  NOR2_X1 U624 ( .A1(n637), .A2(n541), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n542), .A2(n628), .ZN(n543) );
  NOR2_X1 U626 ( .A1(n615), .A2(n543), .ZN(n544) );
  NAND2_X1 U627 ( .A1(n555), .A2(n544), .ZN(n578) );
  NOR2_X1 U628 ( .A1(n545), .A2(n578), .ZN(n546) );
  XNOR2_X1 U629 ( .A(n546), .B(KEYINPUT36), .ZN(n547) );
  NAND2_X1 U630 ( .A1(n547), .A2(n579), .ZN(n623) );
  NAND2_X1 U631 ( .A1(n647), .A2(n628), .ZN(n548) );
  XNOR2_X1 U632 ( .A(n548), .B(KEYINPUT30), .ZN(n549) );
  NOR2_X1 U633 ( .A1(n550), .A2(n549), .ZN(n552) );
  INV_X1 U634 ( .A(n627), .ZN(n553) );
  XNOR2_X1 U635 ( .A(n554), .B(KEYINPUT40), .ZN(n714) );
  NAND2_X1 U636 ( .A1(n647), .A2(n555), .ZN(n557) );
  XNOR2_X1 U637 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n556) );
  XNOR2_X1 U638 ( .A(n557), .B(n556), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n559), .A2(n558), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n628), .A2(n627), .ZN(n631) );
  NOR2_X1 U641 ( .A1(n631), .A2(n630), .ZN(n561) );
  XNOR2_X1 U642 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n560) );
  XNOR2_X1 U643 ( .A(n561), .B(n560), .ZN(n661) );
  NOR2_X1 U644 ( .A1(n565), .A2(n661), .ZN(n562) );
  XNOR2_X1 U645 ( .A(n562), .B(KEYINPUT42), .ZN(n715) );
  NOR2_X1 U646 ( .A1(n714), .A2(n715), .ZN(n563) );
  XNOR2_X1 U647 ( .A(n563), .B(KEYINPUT46), .ZN(n564) );
  INV_X1 U648 ( .A(n565), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n613) );
  INV_X1 U650 ( .A(n568), .ZN(n632) );
  NOR2_X1 U651 ( .A1(n613), .A2(n632), .ZN(n569) );
  XOR2_X1 U652 ( .A(KEYINPUT47), .B(n569), .Z(n574) );
  NOR2_X1 U653 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U654 ( .A1(n572), .A2(n582), .ZN(n612) );
  INV_X1 U655 ( .A(n612), .ZN(n573) );
  NOR2_X1 U656 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U657 ( .A(KEYINPUT48), .B(KEYINPUT72), .Z(n576) );
  OR2_X1 U658 ( .A1(n619), .A2(n577), .ZN(n625) );
  NOR2_X1 U659 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U660 ( .A(n580), .B(KEYINPUT43), .ZN(n581) );
  NOR2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n626) );
  INV_X1 U662 ( .A(n626), .ZN(n583) );
  AND2_X1 U663 ( .A1(n625), .A2(n583), .ZN(n584) );
  XOR2_X1 U664 ( .A(n586), .B(KEYINPUT84), .Z(n587) );
  NAND2_X1 U665 ( .A1(n587), .A2(KEYINPUT2), .ZN(n588) );
  INV_X1 U666 ( .A(KEYINPUT2), .ZN(n589) );
  OR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U668 ( .A1(n667), .A2(n591), .ZN(n671) );
  XOR2_X1 U669 ( .A(KEYINPUT88), .B(KEYINPUT80), .Z(n596) );
  XNOR2_X1 U670 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n595) );
  XNOR2_X1 U671 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT86), .B(KEYINPUT123), .ZN(n599) );
  INV_X1 U673 ( .A(KEYINPUT56), .ZN(n598) );
  XNOR2_X1 U674 ( .A(G101), .B(n600), .ZN(G3) );
  NOR2_X1 U675 ( .A1(n615), .A2(n602), .ZN(n601) );
  XOR2_X1 U676 ( .A(G104), .B(n601), .Z(G6) );
  NOR2_X1 U677 ( .A1(n602), .A2(n619), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n604) );
  XNOR2_X1 U679 ( .A(G107), .B(KEYINPUT111), .ZN(n603) );
  XNOR2_X1 U680 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n606), .B(n605), .ZN(G9) );
  XNOR2_X1 U682 ( .A(G110), .B(n607), .ZN(G12) );
  NOR2_X1 U683 ( .A1(n613), .A2(n619), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n609) );
  XNOR2_X1 U685 ( .A(G128), .B(KEYINPUT113), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n611), .B(n610), .ZN(G30) );
  XNOR2_X1 U688 ( .A(G143), .B(n612), .ZN(G45) );
  NOR2_X1 U689 ( .A1(n615), .A2(n613), .ZN(n614) );
  XOR2_X1 U690 ( .A(G146), .B(n614), .Z(G48) );
  NOR2_X1 U691 ( .A1(n615), .A2(n618), .ZN(n616) );
  XOR2_X1 U692 ( .A(KEYINPUT114), .B(n616), .Z(n617) );
  XNOR2_X1 U693 ( .A(G113), .B(n617), .ZN(G15) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U695 ( .A(G116), .B(n620), .Z(G18) );
  XOR2_X1 U696 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n622) );
  XNOR2_X1 U697 ( .A(G125), .B(KEYINPUT37), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(n624) );
  XOR2_X1 U699 ( .A(n624), .B(n623), .Z(G27) );
  XNOR2_X1 U700 ( .A(G134), .B(n625), .ZN(G36) );
  XOR2_X1 U701 ( .A(G140), .B(n626), .Z(G42) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U706 ( .A1(n660), .A2(n635), .ZN(n654) );
  OR2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n638), .B(KEYINPUT49), .ZN(n639) );
  XNOR2_X1 U709 ( .A(KEYINPUT117), .B(n639), .ZN(n645) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U712 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U713 ( .A(n648), .B(KEYINPUT119), .ZN(n650) );
  NAND2_X1 U714 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U715 ( .A(KEYINPUT51), .B(n651), .ZN(n652) );
  NOR2_X1 U716 ( .A1(n661), .A2(n652), .ZN(n653) );
  NOR2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n656) );
  NOR2_X1 U718 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U719 ( .A(KEYINPUT121), .B(n659), .Z(n663) );
  NOR2_X1 U720 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U721 ( .A(n664), .B(KEYINPUT122), .ZN(n665) );
  NAND2_X1 U722 ( .A1(n665), .A2(n704), .ZN(n675) );
  XNOR2_X1 U723 ( .A(KEYINPUT2), .B(KEYINPUT81), .ZN(n669) );
  NAND2_X1 U724 ( .A1(n701), .A2(n669), .ZN(n666) );
  XNOR2_X1 U725 ( .A(KEYINPUT83), .B(n666), .ZN(n673) );
  BUF_X1 U726 ( .A(n667), .Z(n668) );
  NAND2_X1 U727 ( .A1(n668), .A2(n669), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U729 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U730 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U731 ( .A(KEYINPUT53), .B(n676), .ZN(G75) );
  XOR2_X1 U732 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n678) );
  NAND2_X1 U733 ( .A1(n685), .A2(G469), .ZN(n677) );
  NOR2_X1 U734 ( .A1(n689), .A2(n680), .ZN(G54) );
  NAND2_X1 U735 ( .A1(G478), .A2(n685), .ZN(n682) );
  XNOR2_X1 U736 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U737 ( .A1(n689), .A2(n684), .ZN(G63) );
  NAND2_X1 U738 ( .A1(G217), .A2(n685), .ZN(n686) );
  XNOR2_X1 U739 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U740 ( .A1(n689), .A2(n688), .ZN(G66) );
  OR2_X1 U741 ( .A1(G953), .A2(n668), .ZN(n693) );
  NAND2_X1 U742 ( .A1(G953), .A2(G224), .ZN(n690) );
  XNOR2_X1 U743 ( .A(KEYINPUT61), .B(n690), .ZN(n691) );
  NAND2_X1 U744 ( .A1(n691), .A2(G898), .ZN(n692) );
  NAND2_X1 U745 ( .A1(n693), .A2(n692), .ZN(n698) );
  XOR2_X1 U746 ( .A(n694), .B(KEYINPUT124), .Z(n695) );
  NOR2_X1 U747 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U748 ( .A(n698), .B(n697), .ZN(G69) );
  XNOR2_X1 U749 ( .A(n700), .B(n699), .ZN(n707) );
  XOR2_X1 U750 ( .A(n707), .B(KEYINPUT125), .Z(n702) );
  XNOR2_X1 U751 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U752 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U753 ( .A(n705), .B(KEYINPUT126), .ZN(n711) );
  XOR2_X1 U754 ( .A(G227), .B(KEYINPUT127), .Z(n706) );
  XNOR2_X1 U755 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U756 ( .A1(n708), .A2(G900), .ZN(n709) );
  NAND2_X1 U757 ( .A1(n709), .A2(G953), .ZN(n710) );
  NAND2_X1 U758 ( .A1(n711), .A2(n710), .ZN(G72) );
  XOR2_X1 U759 ( .A(n712), .B(G122), .Z(G24) );
  XNOR2_X1 U760 ( .A(n713), .B(G119), .ZN(G21) );
  XOR2_X1 U761 ( .A(n714), .B(G131), .Z(G33) );
  XOR2_X1 U762 ( .A(G137), .B(n715), .Z(G39) );
endmodule

