

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747;

  OR2_X2 U371 ( .A1(n652), .A2(G902), .ZN(n421) );
  NOR2_X2 U372 ( .A1(n535), .A2(n696), .ZN(n536) );
  XNOR2_X2 U373 ( .A(n470), .B(KEYINPUT4), .ZN(n492) );
  AND2_X1 U374 ( .A1(n398), .A2(n397), .ZN(n606) );
  AND2_X1 U375 ( .A1(n368), .A2(n600), .ZN(n367) );
  NAND2_X1 U376 ( .A1(n575), .A2(n574), .ZN(n576) );
  OR2_X1 U377 ( .A1(n582), .A2(n565), .ZN(n567) );
  XNOR2_X1 U378 ( .A(n499), .B(n498), .ZN(n512) );
  OR2_X1 U379 ( .A1(n665), .A2(G902), .ZN(n507) );
  XNOR2_X1 U380 ( .A(G101), .B(KEYINPUT90), .ZN(n409) );
  XNOR2_X1 U381 ( .A(KEYINPUT16), .B(G122), .ZN(n494) );
  XNOR2_X1 U382 ( .A(G116), .B(G113), .ZN(n410) );
  XNOR2_X1 U383 ( .A(G110), .B(G107), .ZN(n493) );
  XNOR2_X2 U384 ( .A(n392), .B(n349), .ZN(n562) );
  NOR2_X2 U385 ( .A1(n649), .A2(n747), .ZN(n545) );
  XOR2_X1 U386 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n467) );
  AND2_X1 U387 ( .A1(n399), .A2(n400), .ZN(n398) );
  NOR2_X1 U388 ( .A1(n602), .A2(n401), .ZN(n400) );
  AND2_X1 U389 ( .A1(n405), .A2(n402), .ZN(n401) );
  XNOR2_X1 U390 ( .A(n425), .B(n424), .ZN(n426) );
  INV_X1 U391 ( .A(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U392 ( .A(G119), .B(G110), .ZN(n425) );
  AND2_X2 U393 ( .A1(n367), .A2(n364), .ZN(n601) );
  INV_X1 U394 ( .A(KEYINPUT36), .ZN(n373) );
  XNOR2_X1 U395 ( .A(n391), .B(n352), .ZN(n390) );
  XNOR2_X1 U396 ( .A(n381), .B(n437), .ZN(n438) );
  XNOR2_X1 U397 ( .A(n416), .B(KEYINPUT73), .ZN(n456) );
  INV_X1 U398 ( .A(KEYINPUT82), .ZN(n402) );
  INV_X1 U399 ( .A(KEYINPUT2), .ZN(n405) );
  NOR2_X1 U400 ( .A1(KEYINPUT76), .A2(G953), .ZN(n357) );
  NAND2_X1 U401 ( .A1(n358), .A2(KEYINPUT76), .ZN(n362) );
  INV_X1 U402 ( .A(G224), .ZN(n358) );
  XNOR2_X1 U403 ( .A(n436), .B(n382), .ZN(n440) );
  XNOR2_X1 U404 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n382) );
  XNOR2_X1 U405 ( .A(G143), .B(G104), .ZN(n454) );
  XOR2_X1 U406 ( .A(KEYINPUT12), .B(G122), .Z(n455) );
  XNOR2_X1 U407 ( .A(n492), .B(n408), .ZN(n739) );
  NAND2_X1 U408 ( .A1(n360), .A2(n359), .ZN(n395) );
  AND2_X1 U409 ( .A1(n362), .A2(n361), .ZN(n360) );
  NAND2_X1 U410 ( .A1(n357), .A2(G224), .ZN(n359) );
  NAND2_X1 U411 ( .A1(KEYINPUT76), .A2(G953), .ZN(n361) );
  XNOR2_X1 U412 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n394) );
  XNOR2_X1 U413 ( .A(n491), .B(n490), .ZN(n396) );
  XOR2_X1 U414 ( .A(KEYINPUT91), .B(KEYINPUT89), .Z(n491) );
  NAND2_X1 U415 ( .A1(n440), .A2(G217), .ZN(n381) );
  INV_X1 U416 ( .A(KEYINPUT83), .ZN(n378) );
  XOR2_X1 U417 ( .A(G122), .B(G107), .Z(n475) );
  XNOR2_X1 U418 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n466) );
  XNOR2_X1 U419 ( .A(n739), .B(G146), .ZN(n506) );
  OR2_X1 U420 ( .A1(n580), .A2(n678), .ZN(n581) );
  NAND2_X1 U421 ( .A1(n375), .A2(n374), .ZN(n580) );
  INV_X2 U422 ( .A(G953), .ZN(n711) );
  NAND2_X1 U423 ( .A1(n512), .A2(n511), .ZN(n392) );
  XNOR2_X1 U424 ( .A(n519), .B(n518), .ZN(n385) );
  XNOR2_X1 U425 ( .A(n427), .B(n426), .ZN(n431) );
  XNOR2_X1 U426 ( .A(n538), .B(n537), .ZN(n649) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n647) );
  INV_X1 U428 ( .A(KEYINPUT114), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n500), .B(n373), .ZN(n372) );
  NAND2_X1 U430 ( .A1(n390), .A2(n350), .ZN(n389) );
  XNOR2_X1 U431 ( .A(n380), .B(KEYINPUT28), .ZN(n379) );
  NOR2_X1 U432 ( .A1(n515), .A2(n587), .ZN(n380) );
  XOR2_X1 U433 ( .A(n513), .B(KEYINPUT66), .Z(n349) );
  XOR2_X1 U434 ( .A(n584), .B(KEYINPUT78), .Z(n350) );
  NAND2_X1 U435 ( .A1(n573), .A2(n376), .ZN(n351) );
  OR2_X1 U436 ( .A1(n570), .A2(n521), .ZN(n677) );
  INV_X1 U437 ( .A(n677), .ZN(n374) );
  XOR2_X1 U438 ( .A(n583), .B(KEYINPUT34), .Z(n352) );
  XOR2_X1 U439 ( .A(n741), .B(KEYINPUT126), .Z(n353) );
  XNOR2_X1 U440 ( .A(KEYINPUT15), .B(G902), .ZN(n602) );
  INV_X1 U441 ( .A(n602), .ZN(n404) );
  XOR2_X1 U442 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n354) );
  NAND2_X1 U443 ( .A1(n622), .A2(n602), .ZN(n499) );
  XNOR2_X1 U444 ( .A(n355), .B(n643), .ZN(n622) );
  XNOR2_X1 U445 ( .A(n356), .B(n492), .ZN(n355) );
  XNOR2_X1 U446 ( .A(n393), .B(n396), .ZN(n356) );
  INV_X1 U447 ( .A(n575), .ZN(n650) );
  XNOR2_X2 U448 ( .A(n363), .B(KEYINPUT32), .ZN(n575) );
  NAND2_X1 U449 ( .A1(n573), .A2(n406), .ZN(n363) );
  XNOR2_X2 U450 ( .A(n567), .B(n566), .ZN(n573) );
  NAND2_X1 U451 ( .A1(n365), .A2(n634), .ZN(n364) );
  NAND2_X1 U452 ( .A1(n366), .A2(n579), .ZN(n365) );
  NAND2_X1 U453 ( .A1(n586), .A2(n577), .ZN(n366) );
  NAND2_X1 U454 ( .A1(n369), .A2(KEYINPUT44), .ZN(n368) );
  NAND2_X1 U455 ( .A1(n586), .A2(n634), .ZN(n369) );
  NOR2_X1 U456 ( .A1(n647), .A2(n534), .ZN(n547) );
  NAND2_X1 U457 ( .A1(n372), .A2(n589), .ZN(n371) );
  NOR2_X1 U458 ( .A1(n376), .A2(n515), .ZN(n452) );
  INV_X1 U459 ( .A(n376), .ZN(n375) );
  AND2_X1 U460 ( .A1(n569), .A2(n376), .ZN(n406) );
  XNOR2_X2 U461 ( .A(n591), .B(KEYINPUT6), .ZN(n376) );
  NAND2_X1 U462 ( .A1(n377), .A2(n404), .ZN(n603) );
  INV_X1 U463 ( .A(n403), .ZN(n377) );
  AND2_X1 U464 ( .A1(n403), .A2(n354), .ZN(n670) );
  XNOR2_X1 U465 ( .A(n403), .B(n353), .ZN(n740) );
  XNOR2_X2 U466 ( .A(n607), .B(n378), .ZN(n403) );
  XNOR2_X2 U467 ( .A(n507), .B(G469), .ZN(n522) );
  AND2_X2 U468 ( .A1(n379), .A2(n522), .ZN(n732) );
  INV_X1 U469 ( .A(n591), .ZN(n587) );
  NAND2_X1 U470 ( .A1(n451), .A2(n570), .ZN(n515) );
  NAND2_X1 U471 ( .A1(n383), .A2(n555), .ZN(n607) );
  XNOR2_X1 U472 ( .A(n384), .B(n548), .ZN(n383) );
  NAND2_X1 U473 ( .A1(n546), .A2(n547), .ZN(n384) );
  NAND2_X1 U474 ( .A1(n386), .A2(n385), .ZN(n535) );
  NOR2_X1 U475 ( .A1(n677), .A2(n387), .ZN(n386) );
  NAND2_X1 U476 ( .A1(n522), .A2(n520), .ZN(n387) );
  NAND2_X1 U477 ( .A1(n374), .A2(n522), .ZN(n592) );
  XNOR2_X2 U478 ( .A(n388), .B(G143), .ZN(n470) );
  XNOR2_X2 U479 ( .A(G128), .B(KEYINPUT64), .ZN(n388) );
  NAND2_X1 U480 ( .A1(n591), .A2(n511), .ZN(n519) );
  XNOR2_X2 U481 ( .A(n421), .B(G472), .ZN(n591) );
  XNOR2_X2 U482 ( .A(n389), .B(n585), .ZN(n634) );
  NAND2_X1 U483 ( .A1(n710), .A2(n594), .ZN(n391) );
  INV_X1 U484 ( .A(n562), .ZN(n527) );
  XNOR2_X1 U485 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X1 U486 ( .A(G146), .B(G125), .ZN(n490) );
  NAND2_X1 U487 ( .A1(n635), .A2(n405), .ZN(n397) );
  XNOR2_X2 U488 ( .A(n601), .B(KEYINPUT45), .ZN(n635) );
  NAND2_X1 U489 ( .A1(n403), .A2(n405), .ZN(n399) );
  XNOR2_X1 U490 ( .A(n564), .B(n563), .ZN(n582) );
  INV_X1 U491 ( .A(KEYINPUT47), .ZN(n530) );
  INV_X1 U492 ( .A(G237), .ZN(n415) );
  NAND2_X1 U493 ( .A1(n711), .A2(n415), .ZN(n416) );
  INV_X1 U494 ( .A(KEYINPUT48), .ZN(n548) );
  INV_X1 U495 ( .A(KEYINPUT56), .ZN(n627) );
  INV_X1 U496 ( .A(KEYINPUT110), .ZN(n453) );
  XNOR2_X1 U497 ( .A(G134), .B(G131), .ZN(n407) );
  XNOR2_X1 U498 ( .A(n407), .B(G137), .ZN(n408) );
  XNOR2_X1 U499 ( .A(n410), .B(n409), .ZN(n412) );
  XNOR2_X1 U500 ( .A(KEYINPUT3), .B(G119), .ZN(n411) );
  XNOR2_X1 U501 ( .A(n412), .B(n411), .ZN(n496) );
  XNOR2_X1 U502 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n414) );
  XNOR2_X1 U503 ( .A(KEYINPUT72), .B(KEYINPUT98), .ZN(n413) );
  XNOR2_X1 U504 ( .A(n414), .B(n413), .ZN(n418) );
  AND2_X1 U505 ( .A1(n456), .A2(G210), .ZN(n417) );
  XNOR2_X1 U506 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U507 ( .A(n496), .B(n419), .ZN(n420) );
  XNOR2_X1 U508 ( .A(n506), .B(n420), .ZN(n652) );
  XOR2_X1 U509 ( .A(KEYINPUT95), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U510 ( .A(G128), .B(G137), .ZN(n422) );
  XNOR2_X1 U511 ( .A(n423), .B(n422), .ZN(n427) );
  NAND2_X1 U512 ( .A1(n711), .A2(G234), .ZN(n429) );
  XNOR2_X1 U513 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n428) );
  XNOR2_X1 U514 ( .A(n429), .B(n428), .ZN(n473) );
  NAND2_X1 U515 ( .A1(n473), .A2(G221), .ZN(n430) );
  XNOR2_X1 U516 ( .A(n431), .B(n430), .ZN(n435) );
  INV_X1 U517 ( .A(G140), .ZN(n432) );
  XNOR2_X1 U518 ( .A(n490), .B(n432), .ZN(n434) );
  XOR2_X1 U519 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n433) );
  XNOR2_X1 U520 ( .A(n434), .B(n433), .ZN(n738) );
  XNOR2_X1 U521 ( .A(n435), .B(n738), .ZN(n612) );
  INV_X1 U522 ( .A(G902), .ZN(n484) );
  NAND2_X1 U523 ( .A1(n612), .A2(n484), .ZN(n439) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n437) );
  NAND2_X1 U525 ( .A1(n602), .A2(G234), .ZN(n436) );
  XNOR2_X1 U526 ( .A(n439), .B(n438), .ZN(n570) );
  NAND2_X1 U527 ( .A1(n440), .A2(G221), .ZN(n442) );
  INV_X1 U528 ( .A(KEYINPUT21), .ZN(n441) );
  XNOR2_X1 U529 ( .A(n442), .B(n441), .ZN(n681) );
  XOR2_X1 U530 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n444) );
  NAND2_X1 U531 ( .A1(G234), .A2(G237), .ZN(n443) );
  XNOR2_X1 U532 ( .A(n444), .B(n443), .ZN(n448) );
  NAND2_X1 U533 ( .A1(G902), .A2(n448), .ZN(n556) );
  NOR2_X1 U534 ( .A1(G900), .A2(n556), .ZN(n445) );
  NAND2_X1 U535 ( .A1(G953), .A2(n445), .ZN(n447) );
  INV_X1 U536 ( .A(KEYINPUT109), .ZN(n446) );
  XNOR2_X1 U537 ( .A(n447), .B(n446), .ZN(n450) );
  NAND2_X1 U538 ( .A1(n448), .A2(G952), .ZN(n449) );
  XNOR2_X1 U539 ( .A(n449), .B(KEYINPUT93), .ZN(n707) );
  NAND2_X1 U540 ( .A1(n707), .A2(n711), .ZN(n560) );
  NAND2_X1 U541 ( .A1(n450), .A2(n560), .ZN(n520) );
  AND2_X1 U542 ( .A1(n681), .A2(n520), .ZN(n451) );
  XNOR2_X1 U543 ( .A(n453), .B(n452), .ZN(n489) );
  XNOR2_X1 U544 ( .A(n455), .B(n454), .ZN(n458) );
  NAND2_X1 U545 ( .A1(G214), .A2(n456), .ZN(n457) );
  XOR2_X1 U546 ( .A(n458), .B(n457), .Z(n461) );
  XNOR2_X1 U547 ( .A(G113), .B(G131), .ZN(n459) );
  XNOR2_X1 U548 ( .A(n459), .B(KEYINPUT11), .ZN(n460) );
  XNOR2_X1 U549 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U550 ( .A(n462), .B(n738), .Z(n616) );
  NOR2_X2 U551 ( .A1(n616), .A2(G902), .ZN(n464) );
  XNOR2_X1 U552 ( .A(KEYINPUT13), .B(G475), .ZN(n463) );
  XNOR2_X2 U553 ( .A(n464), .B(n463), .ZN(n540) );
  INV_X1 U554 ( .A(KEYINPUT100), .ZN(n465) );
  XNOR2_X1 U555 ( .A(n540), .B(n465), .ZN(n509) );
  INV_X1 U556 ( .A(n509), .ZN(n483) );
  XNOR2_X1 U557 ( .A(n467), .B(n466), .ZN(n469) );
  XOR2_X1 U558 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n468) );
  XNOR2_X1 U559 ( .A(n469), .B(n468), .ZN(n472) );
  INV_X1 U560 ( .A(n470), .ZN(n471) );
  XNOR2_X1 U561 ( .A(n472), .B(n471), .ZN(n479) );
  NAND2_X1 U562 ( .A1(n473), .A2(G217), .ZN(n477) );
  XNOR2_X1 U563 ( .A(G116), .B(G134), .ZN(n474) );
  XNOR2_X1 U564 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U565 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U566 ( .A(n479), .B(n478), .ZN(n659) );
  NOR2_X1 U567 ( .A1(n659), .A2(G902), .ZN(n480) );
  XNOR2_X1 U568 ( .A(n480), .B(G478), .ZN(n481) );
  XNOR2_X1 U569 ( .A(n481), .B(KEYINPUT105), .ZN(n539) );
  INV_X1 U570 ( .A(n539), .ZN(n482) );
  NAND2_X1 U571 ( .A1(n483), .A2(n482), .ZN(n730) );
  INV_X1 U572 ( .A(n730), .ZN(n487) );
  NAND2_X1 U573 ( .A1(n484), .A2(n415), .ZN(n497) );
  NAND2_X1 U574 ( .A1(n497), .A2(G214), .ZN(n486) );
  INV_X1 U575 ( .A(KEYINPUT92), .ZN(n485) );
  XNOR2_X1 U576 ( .A(n486), .B(n485), .ZN(n695) );
  INV_X1 U577 ( .A(n695), .ZN(n511) );
  NAND2_X1 U578 ( .A1(n487), .A2(n511), .ZN(n488) );
  NOR2_X2 U579 ( .A1(n489), .A2(n488), .ZN(n549) );
  XNOR2_X1 U580 ( .A(n493), .B(G104), .ZN(n503) );
  XNOR2_X1 U581 ( .A(n503), .B(n494), .ZN(n495) );
  XNOR2_X1 U582 ( .A(n496), .B(n495), .ZN(n643) );
  AND2_X1 U583 ( .A1(n497), .A2(G210), .ZN(n498) );
  BUF_X1 U584 ( .A(n512), .Z(n552) );
  NAND2_X1 U585 ( .A1(n549), .A2(n552), .ZN(n500) );
  XOR2_X1 U586 ( .A(G101), .B(G140), .Z(n502) );
  NAND2_X1 U587 ( .A1(G227), .A2(n711), .ZN(n501) );
  XNOR2_X1 U588 ( .A(n502), .B(n501), .ZN(n504) );
  XNOR2_X1 U589 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U590 ( .A(n506), .B(n505), .ZN(n665) );
  XNOR2_X1 U591 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n508) );
  XNOR2_X1 U592 ( .A(n522), .B(n508), .ZN(n678) );
  NAND2_X1 U593 ( .A1(n509), .A2(n539), .ZN(n510) );
  XNOR2_X2 U594 ( .A(n510), .B(KEYINPUT106), .ZN(n734) );
  NAND2_X1 U595 ( .A1(n734), .A2(n730), .ZN(n692) );
  NOR2_X1 U596 ( .A1(n692), .A2(KEYINPUT70), .ZN(n514) );
  XNOR2_X1 U597 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n513) );
  NAND2_X1 U598 ( .A1(n514), .A2(n562), .ZN(n517) );
  INV_X1 U599 ( .A(n732), .ZN(n516) );
  NOR2_X1 U600 ( .A1(n517), .A2(n516), .ZN(n526) );
  INV_X1 U601 ( .A(KEYINPUT30), .ZN(n518) );
  INV_X1 U602 ( .A(n681), .ZN(n521) );
  INV_X1 U603 ( .A(n535), .ZN(n525) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n584) );
  INV_X1 U605 ( .A(n552), .ZN(n523) );
  NOR2_X1 U606 ( .A1(n584), .A2(n523), .ZN(n524) );
  AND2_X1 U607 ( .A1(n525), .A2(n524), .ZN(n729) );
  NOR2_X1 U608 ( .A1(n526), .A2(n729), .ZN(n533) );
  NAND2_X1 U609 ( .A1(n692), .A2(KEYINPUT70), .ZN(n528) );
  NOR2_X1 U610 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U611 ( .A1(n529), .A2(n732), .ZN(n531) );
  XNOR2_X1 U612 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U613 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U614 ( .A(n552), .B(KEYINPUT38), .ZN(n696) );
  XNOR2_X1 U615 ( .A(n536), .B(KEYINPUT39), .ZN(n554) );
  NOR2_X1 U616 ( .A1(n554), .A2(n730), .ZN(n538) );
  XOR2_X1 U617 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n537) );
  NOR2_X1 U618 ( .A1(n696), .A2(n695), .ZN(n693) );
  NOR2_X1 U619 ( .A1(n540), .A2(n539), .ZN(n698) );
  NAND2_X1 U620 ( .A1(n693), .A2(n698), .ZN(n541) );
  XNOR2_X1 U621 ( .A(n541), .B(KEYINPUT41), .ZN(n709) );
  NAND2_X1 U622 ( .A1(n709), .A2(n732), .ZN(n544) );
  XNOR2_X1 U623 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n542) );
  XNOR2_X1 U624 ( .A(n542), .B(KEYINPUT42), .ZN(n543) );
  XNOR2_X1 U625 ( .A(n544), .B(n543), .ZN(n747) );
  XNOR2_X1 U626 ( .A(n545), .B(KEYINPUT46), .ZN(n546) );
  INV_X1 U627 ( .A(n549), .ZN(n550) );
  INV_X1 U628 ( .A(n678), .ZN(n589) );
  NOR2_X1 U629 ( .A1(n550), .A2(n589), .ZN(n551) );
  XNOR2_X1 U630 ( .A(n551), .B(KEYINPUT43), .ZN(n553) );
  NOR2_X1 U631 ( .A1(n553), .A2(n552), .ZN(n631) );
  NOR2_X1 U632 ( .A1(n554), .A2(n734), .ZN(n630) );
  NOR2_X1 U633 ( .A1(n631), .A2(n630), .ZN(n555) );
  INV_X1 U634 ( .A(n556), .ZN(n558) );
  NOR2_X1 U635 ( .A1(G898), .A2(n711), .ZN(n557) );
  XNOR2_X1 U636 ( .A(KEYINPUT94), .B(n557), .ZN(n642) );
  NAND2_X1 U637 ( .A1(n558), .A2(n642), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U639 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U640 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n563) );
  NAND2_X1 U641 ( .A1(n698), .A2(n681), .ZN(n565) );
  INV_X1 U642 ( .A(KEYINPUT22), .ZN(n566) );
  INV_X1 U643 ( .A(KEYINPUT108), .ZN(n568) );
  XNOR2_X1 U644 ( .A(n570), .B(n568), .ZN(n680) );
  NOR2_X1 U645 ( .A1(n678), .A2(n680), .ZN(n569) );
  AND2_X1 U646 ( .A1(n587), .A2(n570), .ZN(n571) );
  AND2_X1 U647 ( .A1(n678), .A2(n571), .ZN(n572) );
  AND2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n648) );
  INV_X1 U649 ( .A(n648), .ZN(n574) );
  XNOR2_X2 U650 ( .A(n576), .B(KEYINPUT86), .ZN(n578) );
  INV_X1 U651 ( .A(n578), .ZN(n586) );
  NOR2_X1 U652 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n578), .A2(KEYINPUT85), .ZN(n579) );
  XNOR2_X2 U654 ( .A(n581), .B(KEYINPUT33), .ZN(n710) );
  INV_X1 U655 ( .A(n582), .ZN(n594) );
  INV_X1 U656 ( .A(KEYINPUT69), .ZN(n583) );
  XNOR2_X1 U657 ( .A(KEYINPUT77), .B(KEYINPUT35), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n587), .A2(n677), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n687) );
  NOR2_X1 U660 ( .A1(n687), .A2(n582), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT31), .ZN(n735) );
  BUF_X1 U662 ( .A(n591), .Z(n683) );
  NOR2_X1 U663 ( .A1(n592), .A2(n683), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n722) );
  NAND2_X1 U665 ( .A1(n735), .A2(n722), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n595), .A2(n692), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n596), .B(KEYINPUT107), .ZN(n599) );
  XNOR2_X1 U668 ( .A(n351), .B(KEYINPUT84), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n678), .A2(n680), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n633) );
  NOR2_X1 U671 ( .A1(n599), .A2(n633), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n603), .A2(n635), .ZN(n604) );
  NOR2_X1 U673 ( .A1(n604), .A2(KEYINPUT82), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n611) );
  INV_X1 U675 ( .A(n607), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n608), .A2(KEYINPUT2), .ZN(n609) );
  NOR2_X1 U677 ( .A1(n635), .A2(n609), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n610), .B(KEYINPUT74), .ZN(n675) );
  NOR2_X2 U679 ( .A1(n611), .A2(n675), .ZN(n651) );
  BUF_X2 U680 ( .A(n651), .Z(n663) );
  NAND2_X1 U681 ( .A1(n663), .A2(G217), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n613), .B(n612), .ZN(n615) );
  INV_X1 U683 ( .A(G952), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n614), .A2(G953), .ZN(n661) );
  AND2_X1 U685 ( .A1(n615), .A2(n661), .ZN(G66) );
  NAND2_X1 U686 ( .A1(n651), .A2(G475), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n616), .B(KEYINPUT59), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n619), .A2(n661), .ZN(n621) );
  INV_X1 U690 ( .A(KEYINPUT60), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(G60) );
  NAND2_X1 U692 ( .A1(n651), .A2(G210), .ZN(n625) );
  XOR2_X1 U693 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n623) );
  XNOR2_X1 U694 ( .A(n622), .B(n623), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n626), .A2(n661), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(G51) );
  NOR2_X1 U698 ( .A1(n735), .A2(n730), .ZN(n629) );
  XOR2_X1 U699 ( .A(G113), .B(n629), .Z(G15) );
  XOR2_X1 U700 ( .A(G134), .B(n630), .Z(G36) );
  XOR2_X1 U701 ( .A(G140), .B(KEYINPUT119), .Z(n632) );
  XOR2_X1 U702 ( .A(n632), .B(n631), .Z(G42) );
  XOR2_X1 U703 ( .A(G101), .B(n633), .Z(G3) );
  XNOR2_X1 U704 ( .A(n634), .B(G122), .ZN(G24) );
  INV_X1 U705 ( .A(n635), .ZN(n671) );
  NAND2_X1 U706 ( .A1(n671), .A2(n711), .ZN(n641) );
  XOR2_X1 U707 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n637) );
  NAND2_X1 U708 ( .A1(G224), .A2(G953), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U710 ( .A(KEYINPUT124), .B(n638), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n639), .A2(G898), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n645) );
  NOR2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(G69) );
  XNOR2_X1 U715 ( .A(G125), .B(KEYINPUT37), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G27) );
  XOR2_X1 U717 ( .A(G110), .B(n648), .Z(G12) );
  XOR2_X1 U718 ( .A(G131), .B(n649), .Z(G33) );
  XOR2_X1 U719 ( .A(G119), .B(n650), .Z(G21) );
  NAND2_X1 U720 ( .A1(n651), .A2(G472), .ZN(n655) );
  BUF_X1 U721 ( .A(n652), .Z(n653) );
  XOR2_X1 U722 ( .A(KEYINPUT62), .B(n653), .Z(n654) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n656), .A2(n661), .ZN(n658) );
  XOR2_X1 U725 ( .A(KEYINPUT87), .B(KEYINPUT63), .Z(n657) );
  XNOR2_X1 U726 ( .A(n658), .B(n657), .ZN(G57) );
  NAND2_X1 U727 ( .A1(n663), .A2(G478), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n662) );
  INV_X1 U729 ( .A(n661), .ZN(n668) );
  NOR2_X1 U730 ( .A1(n662), .A2(n668), .ZN(G63) );
  NAND2_X1 U731 ( .A1(n663), .A2(G469), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(G54) );
  XNOR2_X1 U736 ( .A(n670), .B(KEYINPUT81), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n635), .A2(n354), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U739 ( .A(KEYINPUT79), .B(n674), .Z(n676) );
  NOR2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n716) );
  XNOR2_X1 U741 ( .A(KEYINPUT123), .B(KEYINPUT52), .ZN(n706) );
  NAND2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U743 ( .A(n679), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT49), .B(n682), .Z(n684) );
  NOR2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n688) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U749 ( .A(KEYINPUT51), .B(n689), .Z(n690) );
  NAND2_X1 U750 ( .A1(n709), .A2(n690), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n691), .B(KEYINPUT120), .ZN(n704) );
  NAND2_X1 U752 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U753 ( .A(KEYINPUT122), .B(n694), .ZN(n701) );
  NAND2_X1 U754 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U756 ( .A(KEYINPUT121), .B(n699), .Z(n700) );
  NAND2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U758 ( .A1(n702), .A2(n710), .ZN(n703) );
  NAND2_X1 U759 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U760 ( .A(n706), .B(n705), .Z(n708) );
  NAND2_X1 U761 ( .A1(n708), .A2(n707), .ZN(n714) );
  NAND2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n712) );
  AND2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U764 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U765 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n717), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U767 ( .A1(n722), .A2(n730), .ZN(n719) );
  XNOR2_X1 U768 ( .A(G104), .B(KEYINPUT115), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(G6) );
  XOR2_X1 U770 ( .A(KEYINPUT116), .B(KEYINPUT26), .Z(n721) );
  XNOR2_X1 U771 ( .A(G107), .B(KEYINPUT27), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n724) );
  NOR2_X1 U773 ( .A1(n722), .A2(n734), .ZN(n723) );
  XOR2_X1 U774 ( .A(n724), .B(n723), .Z(G9) );
  XOR2_X1 U775 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n727) );
  NOR2_X1 U776 ( .A1(n734), .A2(n527), .ZN(n725) );
  NAND2_X1 U777 ( .A1(n725), .A2(n732), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n727), .B(n726), .ZN(n728) );
  XOR2_X1 U779 ( .A(G128), .B(n728), .Z(G30) );
  XOR2_X1 U780 ( .A(G143), .B(n729), .Z(G45) );
  NOR2_X1 U781 ( .A1(n730), .A2(n527), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n733), .B(G146), .ZN(G48) );
  NOR2_X1 U784 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U785 ( .A(KEYINPUT118), .B(n736), .Z(n737) );
  XNOR2_X1 U786 ( .A(G116), .B(n737), .ZN(G18) );
  XNOR2_X1 U787 ( .A(n739), .B(n738), .ZN(n741) );
  NOR2_X1 U788 ( .A1(G953), .A2(n740), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n741), .B(G227), .ZN(n743) );
  NAND2_X1 U790 ( .A1(G900), .A2(G953), .ZN(n742) );
  NOR2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U792 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U793 ( .A(KEYINPUT127), .B(n746), .Z(G72) );
  XOR2_X1 U794 ( .A(G137), .B(n747), .Z(G39) );
endmodule

