//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1319, new_n1320, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1379, new_n1380;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n211), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n202), .A2(new_n203), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT64), .B(G68), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n213), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(new_n234));
  AND3_X1   g0034(.A1(new_n222), .A2(new_n232), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n201), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n254), .A2(new_n256), .A3(G232), .A4(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n254), .A2(new_n256), .A3(G226), .A4(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n257), .B(new_n259), .C1(new_n255), .C2(new_n206), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G238), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT67), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(new_n210), .C1(G41), .C2(G45), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n268), .A2(G274), .A3(new_n264), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n262), .A2(KEYINPUT13), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n267), .A2(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n260), .A2(new_n261), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(G200), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n217), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n210), .B2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT12), .ZN(new_n282));
  OAI21_X1  g0082(.A(G68), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n223), .A2(new_n211), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n282), .A2(new_n285), .A3(G1), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(G1), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n284), .A2(new_n286), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n211), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT71), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n211), .A3(G33), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(G77), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT64), .A2(G68), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT64), .A2(G68), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n297), .A2(new_n298), .A3(new_n211), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G50), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT11), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n302), .A2(new_n303), .A3(new_n280), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n302), .B2(new_n280), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n291), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT13), .B1(new_n262), .B2(new_n272), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n275), .A2(new_n274), .A3(new_n276), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G190), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n278), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(G169), .B1(new_n273), .B2(new_n277), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n308), .B2(new_n309), .ZN(new_n318));
  INV_X1    g0118(.A(new_n315), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n308), .A2(G179), .A3(new_n309), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n306), .B(KEYINPUT76), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n312), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT17), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT8), .B(G58), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT70), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OR3_X1    g0128(.A1(new_n327), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n288), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n330), .B2(new_n281), .ZN(new_n332));
  OAI21_X1  g0132(.A(G58), .B1(new_n297), .B2(new_n298), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT77), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(G58), .C1(new_n297), .C2(new_n298), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n219), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n300), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n254), .A2(new_n256), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n340), .B2(new_n211), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT3), .B(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n338), .A2(KEYINPUT16), .A3(new_n339), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n280), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n337), .A2(G20), .B1(G159), .B2(new_n300), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT78), .ZN(new_n349));
  OAI211_X1 g0149(.A(KEYINPUT7), .B(new_n211), .C1(new_n254), .C2(KEYINPUT78), .ZN(new_n350));
  AOI21_X1  g0150(.A(G20), .B1(new_n254), .B2(new_n256), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(KEYINPUT7), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n223), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT16), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n332), .B1(new_n347), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT79), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n264), .A2(G232), .A3(new_n265), .ZN(new_n357));
  INV_X1    g0157(.A(G87), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n255), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G223), .A2(G1698), .ZN(new_n360));
  INV_X1    g0160(.A(G226), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(G1698), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(new_n362), .B2(new_n342), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n271), .B(new_n357), .C1(new_n363), .C2(new_n264), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(G190), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n264), .A2(G232), .A3(new_n265), .ZN(new_n366));
  INV_X1    g0166(.A(G223), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n258), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n361), .A2(G1698), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n254), .A2(new_n368), .A3(new_n256), .A4(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n359), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n366), .B1(new_n372), .B2(new_n261), .ZN(new_n373));
  AOI21_X1  g0173(.A(G200), .B1(new_n373), .B2(new_n271), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n356), .B1(new_n365), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n261), .ZN(new_n378));
  INV_X1    g0178(.A(G190), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n271), .A4(new_n357), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(KEYINPUT79), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n325), .B1(new_n355), .B2(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n377), .A2(KEYINPUT79), .A3(new_n380), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT79), .B1(new_n377), .B2(new_n380), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n338), .A2(new_n353), .A3(new_n339), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n280), .A3(new_n346), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n390), .A4(new_n332), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n364), .A2(G169), .ZN(new_n394));
  INV_X1    g0194(.A(G179), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(new_n364), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n355), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n393), .B1(new_n355), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G238), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n254), .A2(new_n256), .A3(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT69), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT69), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n340), .B2(new_n258), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n342), .A2(G232), .A3(new_n258), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n207), .B2(new_n342), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n261), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n266), .A2(G244), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT72), .A3(new_n271), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n271), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n414), .A2(G179), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n281), .A2(G77), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G77), .B2(new_n288), .ZN(new_n417));
  INV_X1    g0217(.A(new_n326), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n300), .B1(G20), .B2(G77), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT15), .B(G87), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n292), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(new_n421), .B2(new_n280), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n414), .B2(new_n317), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n414), .A2(G200), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(new_n422), .C1(new_n379), .C2(new_n414), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n324), .A2(new_n392), .A3(new_n399), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n342), .A2(G222), .A3(new_n258), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT68), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n429), .A2(new_n430), .B1(G77), .B2(new_n340), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n430), .B2(new_n429), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n367), .B1(new_n402), .B2(new_n404), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n261), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n266), .A2(G226), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(new_n271), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(G179), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n279), .A2(new_n217), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n328), .A2(new_n329), .A3(new_n293), .A4(new_n295), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n300), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n288), .A2(G50), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(G50), .B2(new_n281), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(G169), .B1(new_n434), .B2(new_n436), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n438), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT10), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n434), .A2(G190), .A3(new_n436), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT9), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n442), .B2(new_n445), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n446), .A2(KEYINPUT9), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT74), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n376), .B1(new_n434), .B2(new_n436), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n450), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT73), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT10), .B1(new_n461), .B2(KEYINPUT74), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n450), .A2(KEYINPUT73), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n454), .A2(new_n453), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n451), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n449), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT80), .B1(new_n428), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n324), .A2(new_n427), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT74), .B1(new_n465), .B2(new_n451), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT10), .B1(new_n471), .B2(new_n458), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n448), .B1(new_n472), .B2(new_n466), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n355), .A2(new_n396), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT18), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n355), .A2(new_n393), .A3(new_n396), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n383), .A2(new_n391), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n470), .A2(new_n473), .A3(new_n474), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n469), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n254), .A2(new_n256), .A3(G244), .A4(new_n258), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n342), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n342), .A2(G250), .A3(G1698), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n261), .ZN(new_n491));
  INV_X1    g0291(.A(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(G1), .ZN(new_n493));
  AND2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G257), .A3(new_n264), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT5), .B(G41), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(G274), .A3(new_n264), .A4(new_n493), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n317), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT84), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n497), .B2(new_n499), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n497), .A2(new_n504), .A3(new_n499), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n491), .B(new_n395), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT81), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n208), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(G97), .A2(G107), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  OAI211_X1 g0315(.A(KEYINPUT81), .B(new_n509), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT82), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n518), .A2(G20), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n300), .A2(G77), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n340), .A2(new_n211), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT7), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT78), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n343), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT78), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n523), .A2(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n522), .B1(new_n529), .B2(new_n207), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n280), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  OR3_X1    g0331(.A1(new_n288), .A2(KEYINPUT83), .A3(G97), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT83), .B1(new_n288), .B2(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n210), .A2(G33), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n439), .A2(new_n288), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n532), .A2(new_n533), .B1(new_n535), .B2(G97), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n531), .A2(KEYINPUT86), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT86), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n352), .A2(G107), .B1(G77), .B2(new_n300), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n518), .A2(G20), .A3(new_n520), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n439), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n536), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n508), .B1(new_n537), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n491), .B1(new_n505), .B2(new_n506), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT85), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(G200), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n500), .B1(new_n490), .B2(new_n261), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G190), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n531), .A2(new_n536), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n546), .B1(new_n545), .B2(G200), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n544), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n288), .A2(G116), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n535), .B2(G116), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n488), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n280), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(KEYINPUT20), .A3(new_n280), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n317), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n261), .B1(new_n493), .B2(new_n498), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT90), .B1(new_n565), .B2(G270), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n496), .A2(new_n264), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT90), .ZN(new_n568));
  INV_X1    g0368(.A(G270), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n499), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n254), .A2(new_n256), .A3(G257), .A4(new_n258), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT91), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT91), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n342), .A2(new_n574), .A3(G257), .A4(new_n258), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n401), .A2(G264), .B1(G303), .B2(new_n340), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n264), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n564), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n577), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n261), .ZN(new_n583));
  INV_X1    g0383(.A(new_n499), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n565), .A2(KEYINPUT90), .A3(G270), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n555), .A2(new_n563), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n583), .A2(new_n587), .A3(new_n588), .A4(G179), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n583), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(KEYINPUT21), .A3(new_n564), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n581), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(G200), .B1(new_n571), .B2(new_n578), .ZN(new_n593));
  INV_X1    g0393(.A(new_n588), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n583), .A3(G190), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n598));
  AND2_X1   g0398(.A1(G33), .A2(G97), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n600));
  NOR2_X1   g0400(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n602), .B2(new_n211), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n254), .A2(new_n256), .A3(new_n211), .A4(G68), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n605));
  OR2_X1    g0405(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n606));
  NAND2_X1  g0406(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n280), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n288), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n420), .ZN(new_n612));
  INV_X1    g0412(.A(new_n420), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n535), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT88), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n610), .A2(new_n614), .A3(new_n617), .A4(new_n612), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n493), .A2(G274), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n210), .A2(G45), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G250), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n261), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n254), .A2(new_n256), .A3(G238), .A4(new_n258), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n254), .A2(new_n256), .A3(G244), .A4(G1698), .ZN(new_n624));
  NAND2_X1  g0424(.A1(G33), .A2(G116), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n622), .B1(new_n626), .B2(new_n261), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n395), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n261), .ZN(new_n629));
  INV_X1    g0429(.A(new_n622), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n317), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n616), .A2(new_n618), .A3(new_n628), .A4(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT89), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n631), .B2(new_n379), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n627), .A2(KEYINPUT89), .A3(G190), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n535), .A2(G87), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n610), .A2(new_n612), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n631), .A2(G200), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n635), .A2(new_n636), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n592), .A2(new_n597), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n254), .A2(new_n256), .A3(G257), .A4(G1698), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n254), .A2(new_n256), .A3(G250), .A4(new_n258), .ZN(new_n644));
  NAND2_X1  g0444(.A1(G33), .A2(G294), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT92), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT92), .A4(new_n645), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n261), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n565), .A2(G264), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n499), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT93), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n650), .A2(KEYINPUT93), .A3(new_n499), .A4(new_n651), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G169), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n395), .B2(new_n652), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n342), .A2(new_n211), .A3(G87), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT22), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT22), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n342), .A2(new_n660), .A3(new_n211), .A4(G87), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT23), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n211), .B2(G107), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n665));
  INV_X1    g0465(.A(new_n625), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n664), .A2(new_n665), .B1(new_n666), .B2(new_n211), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT24), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT24), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n662), .A2(new_n670), .A3(new_n667), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n439), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n611), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT25), .B1(new_n611), .B2(new_n207), .ZN(new_n675));
  INV_X1    g0475(.A(new_n535), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n674), .A2(new_n675), .B1(new_n676), .B2(new_n207), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n657), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(G190), .B1(new_n654), .B2(new_n655), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n652), .A2(new_n376), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n553), .A2(new_n642), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n483), .A2(new_n684), .ZN(G372));
  NAND3_X1  g0485(.A1(new_n631), .A2(KEYINPUT94), .A3(new_n317), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n627), .B2(G169), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n686), .A2(new_n688), .A3(new_n615), .A4(new_n628), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n537), .A2(new_n543), .ZN(new_n690));
  INV_X1    g0490(.A(new_n508), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n551), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n541), .A2(new_n542), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n547), .A4(new_n549), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n640), .A2(new_n689), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n683), .A2(new_n692), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n592), .B1(new_n657), .B2(new_n679), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n689), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT26), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n503), .B(new_n507), .C1(new_n541), .C2(new_n542), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n696), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT95), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n705), .B(new_n701), .C1(new_n696), .C2(new_n702), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n633), .A2(new_n640), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n544), .A2(new_n707), .A3(KEYINPUT26), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n704), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n482), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n321), .B1(new_n318), .B2(new_n319), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n313), .A2(new_n315), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n323), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n312), .B2(new_n424), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n392), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n399), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n472), .A2(new_n466), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n448), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(G369));
  INV_X1    g0520(.A(KEYINPUT98), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n287), .A2(new_n211), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT96), .ZN(new_n724));
  INV_X1    g0524(.A(G213), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n722), .B2(KEYINPUT27), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G343), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n594), .ZN(new_n730));
  OR3_X1    g0530(.A1(new_n592), .A2(new_n597), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT97), .B1(new_n592), .B2(new_n730), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n592), .A2(KEYINPUT97), .A3(new_n730), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n721), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(KEYINPUT98), .A3(G330), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n680), .B(new_n683), .C1(new_n678), .C2(new_n729), .ZN(new_n741));
  INV_X1    g0541(.A(new_n729), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n657), .A2(new_n679), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT99), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n743), .A3(KEYINPUT99), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n680), .A2(new_n742), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n592), .A2(new_n729), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n750), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(new_n753), .ZN(G399));
  INV_X1    g0554(.A(KEYINPUT100), .ZN(new_n755));
  INV_X1    g0555(.A(new_n214), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(G41), .ZN(new_n757));
  INV_X1    g0557(.A(G41), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n214), .A2(KEYINPUT100), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n598), .A2(new_n557), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n761), .A2(new_n210), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n221), .B2(new_n761), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT28), .Z(new_n765));
  INV_X1    g0565(.A(KEYINPUT29), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n766), .B(new_n729), .C1(new_n700), .C2(new_n709), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n544), .A2(new_n707), .A3(new_n701), .ZN(new_n769));
  OAI21_X1  g0569(.A(KEYINPUT26), .B1(new_n696), .B2(new_n702), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n771), .B(new_n689), .C1(new_n699), .C2(new_n698), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n766), .B1(new_n772), .B2(new_n729), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n680), .A2(new_n683), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n775), .A2(new_n553), .A3(new_n642), .A4(new_n729), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n571), .A2(new_n395), .A3(new_n578), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n650), .A2(new_n651), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n548), .A2(new_n627), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n777), .A2(KEYINPUT30), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT30), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n548), .A2(new_n651), .A3(new_n650), .A4(new_n627), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n587), .A2(new_n583), .A3(G179), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n627), .A2(G179), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n590), .A2(new_n652), .A3(new_n545), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n780), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n742), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT31), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT31), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n787), .A2(new_n790), .A3(new_n742), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n737), .B1(new_n776), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n765), .B1(new_n794), .B2(G1), .ZN(G364));
  INV_X1    g0595(.A(new_n740), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n285), .A2(G20), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n210), .B1(new_n797), .B2(G45), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n761), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n796), .B(new_n801), .C1(G330), .C2(new_n735), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n756), .A2(new_n340), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G355), .B1(new_n557), .B2(new_n756), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n756), .A2(new_n342), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G45), .B2(new_n220), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n251), .A2(new_n492), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n217), .B1(G20), .B2(new_n317), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n801), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n812), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n211), .A2(new_n379), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n395), .A2(new_n376), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G326), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n395), .A2(G200), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n211), .A2(G190), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n818), .A2(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G179), .A2(G200), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n211), .B1(new_n825), .B2(G190), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n824), .B1(G294), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT101), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n376), .A2(G179), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n821), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n342), .B1(new_n832), .B2(G283), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n816), .A2(new_n830), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n816), .A2(new_n820), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G303), .A2(new_n835), .B1(new_n837), .B2(G322), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n817), .A2(new_n821), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(KEYINPUT33), .B(G317), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n821), .A2(new_n825), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n840), .A2(new_n841), .B1(new_n843), .B2(G329), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n829), .A2(new_n833), .A3(new_n838), .A4(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT102), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n843), .A2(G159), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT32), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G68), .A2(new_n840), .B1(new_n835), .B2(G87), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n826), .A2(new_n206), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n340), .B1(new_n837), .B2(G58), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n831), .A2(new_n207), .ZN(new_n856));
  INV_X1    g0656(.A(G77), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n818), .A2(new_n201), .B1(new_n822), .B2(new_n857), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n850), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n847), .A2(new_n848), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n811), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n814), .B1(new_n815), .B2(new_n860), .C1(new_n735), .C2(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n802), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G396));
  AND2_X1   g0664(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(G283), .ZN(new_n869));
  INV_X1    g0669(.A(G294), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n836), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n340), .B1(new_n822), .B2(new_n557), .ZN(new_n872));
  INV_X1    g0672(.A(new_n818), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n871), .B(new_n872), .C1(G303), .C2(new_n873), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n834), .A2(new_n207), .B1(new_n842), .B2(new_n823), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G87), .B2(new_n832), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n869), .A2(new_n874), .A3(new_n853), .A4(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G137), .A2(new_n873), .B1(new_n840), .B2(G150), .ZN(new_n878));
  INV_X1    g0678(.A(new_n822), .ZN(new_n879));
  AOI22_X1  g0679(.A1(G143), .A2(new_n837), .B1(new_n879), .B2(G159), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT34), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n342), .B1(new_n831), .B2(new_n203), .ZN(new_n883));
  INV_X1    g0683(.A(G132), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n834), .A2(new_n201), .B1(new_n842), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n883), .B(new_n885), .C1(G58), .C2(new_n827), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n881), .A2(KEYINPUT34), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n877), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n815), .B1(new_n889), .B2(KEYINPUT104), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(KEYINPUT104), .B2(new_n889), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n815), .A2(new_n810), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n891), .B(new_n800), .C1(G77), .C2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT105), .Z(new_n894));
  NOR2_X1   g0694(.A1(new_n424), .A2(new_n742), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n426), .B1(new_n422), .B2(new_n729), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n424), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n810), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n710), .A2(new_n729), .ZN(new_n900));
  INV_X1    g0700(.A(new_n897), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n900), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n792), .B1(new_n684), .B2(new_n742), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n800), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(G384));
  NOR2_X1   g0708(.A1(new_n797), .A2(new_n210), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n727), .B(KEYINPUT107), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n355), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT109), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n383), .A2(new_n391), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n399), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n383), .B2(new_n391), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n390), .A2(new_n332), .A3(new_n375), .A4(new_n381), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n912), .A3(new_n475), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT37), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n919), .A2(new_n912), .A3(new_n475), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n918), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT16), .B1(new_n348), .B2(new_n345), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n332), .B1(new_n347), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n728), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n478), .B2(new_n479), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n396), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n919), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT37), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n923), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n930), .A2(new_n934), .A3(KEYINPUT38), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n910), .B1(new_n925), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n714), .A2(new_n742), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  INV_X1    g0738(.A(new_n332), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n346), .A2(new_n280), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n389), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n941), .A2(new_n386), .B1(new_n927), .B2(new_n728), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n922), .B1(new_n942), .B2(new_n931), .ZN(new_n943));
  AND4_X1   g0743(.A1(new_n922), .A2(new_n919), .A3(new_n912), .A4(new_n475), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n928), .B1(new_n392), .B2(new_n399), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n930), .A2(new_n934), .A3(KEYINPUT38), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(KEYINPUT39), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n936), .A2(new_n937), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n714), .A2(KEYINPUT106), .A3(new_n311), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n323), .A2(new_n742), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n952), .A2(new_n322), .A3(new_n312), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n714), .A2(new_n954), .A3(new_n311), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n951), .A2(new_n953), .B1(new_n955), .B2(new_n952), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n729), .B(new_n897), .C1(new_n700), .C2(new_n709), .ZN(new_n958));
  INV_X1    g0758(.A(new_n895), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT38), .B1(new_n930), .B2(new_n934), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n935), .A2(new_n961), .A3(KEYINPUT108), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT108), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n947), .B2(new_n948), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n960), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n399), .A2(new_n911), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n950), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n482), .B1(new_n768), .B2(new_n773), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(new_n719), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n968), .B(new_n970), .Z(new_n971));
  NAND4_X1  g0771(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n897), .A4(new_n956), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n918), .A2(new_n924), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n938), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n972), .B1(new_n948), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT110), .ZN(new_n976));
  INV_X1    g0776(.A(new_n791), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n790), .B1(new_n787), .B2(new_n742), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND4_X1   g0779(.A1(new_n680), .A2(new_n553), .A3(new_n642), .A4(new_n683), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n729), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n953), .A2(new_n951), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n955), .A2(new_n952), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n983), .A3(new_n897), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n976), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n903), .A2(KEYINPUT110), .A3(new_n897), .A4(new_n956), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n962), .C2(new_n964), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT40), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n975), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n483), .A2(new_n981), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n737), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n990), .B2(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n909), .B1(new_n971), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n971), .B2(new_n992), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n518), .A2(new_n520), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT35), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT35), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n997), .A2(new_n998), .A3(G116), .A4(new_n218), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT36), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n334), .A2(G77), .A3(new_n221), .A4(new_n336), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n247), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(G1), .A3(new_n285), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n994), .A2(new_n1000), .A3(new_n1003), .ZN(G367));
  INV_X1    g0804(.A(new_n805), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n813), .B1(new_n214), .B2(new_n420), .C1(new_n1005), .C2(new_n242), .ZN(new_n1006));
  INV_X1    g0806(.A(G150), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n202), .A2(new_n834), .B1(new_n836), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n340), .B(new_n1008), .C1(G143), .C2(new_n873), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n832), .A2(G77), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n201), .B2(new_n822), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G137), .B2(new_n843), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n827), .A2(G68), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n868), .A2(G159), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n834), .A2(new_n557), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n867), .C2(new_n870), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT116), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G303), .A2(new_n837), .B1(new_n879), .B2(G283), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G97), .A2(new_n832), .B1(new_n843), .B2(G317), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n340), .B1(new_n818), .B2(new_n823), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G107), .B2(new_n827), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1019), .A2(KEYINPUT116), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1015), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT47), .Z(new_n1028));
  OAI211_X1 g0828(.A(new_n800), .B(new_n1006), .C1(new_n1028), .C2(new_n815), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT117), .Z(new_n1030));
  OR2_X1    g0830(.A1(new_n729), .A2(new_n638), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n697), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n689), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1030), .B1(new_n861), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n794), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT115), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n740), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n738), .A2(KEYINPUT115), .A3(new_n739), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n747), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT99), .B1(new_n741), .B2(new_n743), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(KEYINPUT114), .A3(new_n751), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n751), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n748), .A2(new_n752), .ZN(new_n1046));
  OR3_X1    g0846(.A1(new_n1045), .A2(new_n1046), .A3(KEYINPUT114), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1040), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT115), .B1(new_n738), .B2(new_n739), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1049), .A3(new_n1044), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n794), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n694), .A2(new_n729), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n553), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT111), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n508), .B2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n753), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT112), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT112), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n753), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT45), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n753), .A2(new_n1058), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT44), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1060), .A2(KEYINPUT45), .A3(new_n1062), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT113), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1052), .B1(new_n1071), .B2(new_n749), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n749), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1069), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1036), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n760), .B(KEYINPUT41), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n798), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT42), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1045), .B2(new_n1058), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n544), .B2(new_n729), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1058), .B1(new_n1078), .B2(new_n750), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1081), .A2(new_n753), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1080), .A2(new_n1082), .B1(KEYINPUT43), .B2(new_n1033), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1033), .A2(KEYINPUT43), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1073), .A2(new_n1058), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1085), .A2(new_n1073), .A3(new_n1058), .A4(new_n1086), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1035), .B1(new_n1077), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G387));
  NAND2_X1  g0894(.A1(new_n1047), .A2(new_n1044), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n1036), .A3(new_n1050), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1052), .A2(new_n761), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n803), .A2(new_n762), .B1(new_n207), .B2(new_n756), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n239), .A2(new_n492), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n326), .A2(G50), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT50), .ZN(new_n1102));
  AOI211_X1 g0902(.A(G45), .B(new_n762), .C1(G68), .C2(G77), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n805), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1099), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n801), .B1(new_n1106), .B2(new_n813), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G50), .A2(new_n837), .B1(new_n879), .B2(G68), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n827), .A2(new_n613), .ZN(new_n1109));
  INV_X1    g0909(.A(G159), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(new_n1109), .C1(new_n1110), .C2(new_n818), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G77), .A2(new_n835), .B1(new_n843), .B2(G150), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n342), .C1(new_n206), .C2(new_n831), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT118), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1111), .B(new_n1114), .C1(new_n330), .C2(new_n840), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G317), .A2(new_n837), .B1(new_n879), .B2(G303), .ZN(new_n1116));
  INV_X1    g0916(.A(G322), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n818), .C1(new_n867), .C2(new_n823), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1119), .A2(KEYINPUT48), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(KEYINPUT48), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n835), .A2(G294), .B1(new_n827), .B2(G283), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1124), .A2(KEYINPUT49), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n340), .B1(new_n842), .B2(new_n819), .C1(new_n557), .C2(new_n831), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1124), .B2(KEYINPUT49), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1115), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1107), .B1(new_n1128), .B2(new_n815), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1043), .B2(new_n811), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1096), .A2(new_n1050), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n799), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1098), .A2(new_n1132), .ZN(G393));
  AOI21_X1  g0933(.A(new_n760), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1135), .A2(KEYINPUT119), .A3(new_n749), .A4(new_n1065), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1052), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1134), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1136), .A2(new_n1138), .A3(new_n799), .A4(new_n1139), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n813), .B1(new_n206), .B2(new_n214), .C1(new_n1005), .C2(new_n246), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n800), .A2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G317), .A2(new_n873), .B1(new_n837), .B2(G311), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT52), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n868), .A2(G303), .ZN(new_n1148));
  INV_X1    g0948(.A(G283), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n834), .A2(new_n1149), .B1(new_n842), .B2(new_n1117), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G294), .B2(new_n879), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n342), .B(new_n856), .C1(G116), .C2(new_n827), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n223), .A2(new_n835), .B1(new_n843), .B2(G143), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n342), .C1(new_n358), .C2(new_n831), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT120), .Z(new_n1156));
  OAI22_X1  g0956(.A1(new_n818), .A2(new_n1007), .B1(new_n836), .B2(new_n1110), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT51), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n826), .A2(new_n857), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n418), .B2(new_n879), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(new_n201), .C2(new_n867), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1153), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1162), .B2(new_n812), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1058), .B2(new_n861), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1143), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1142), .A2(new_n1165), .ZN(G390));
  NAND2_X1  g0966(.A1(new_n958), .A2(new_n959), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n904), .A2(new_n901), .A3(new_n957), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n956), .B1(new_n793), .B2(new_n897), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n957), .B1(new_n904), .B2(new_n901), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n793), .A2(new_n897), .A3(new_n956), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n896), .A2(new_n424), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n772), .A2(new_n729), .A3(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n959), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n482), .A2(new_n793), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n969), .A2(new_n719), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n937), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1167), .A2(new_n956), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1181), .A2(new_n1182), .B1(new_n936), .B2(new_n949), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n925), .B2(new_n935), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n957), .B1(new_n1174), .B2(new_n959), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1183), .A2(new_n1168), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT39), .B1(new_n974), .B2(new_n948), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n949), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1188), .A2(new_n1189), .B1(new_n937), .B2(new_n960), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1172), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1180), .B1(new_n1187), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1168), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1178), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1190), .A2(new_n1172), .A3(new_n1191), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n761), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(new_n1196), .A3(new_n799), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n809), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n800), .B1(new_n330), .B2(new_n892), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n342), .B(new_n1159), .C1(G87), .C2(new_n835), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n836), .A2(new_n557), .B1(new_n822), .B2(new_n206), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G283), .B2(new_n873), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n207), .C2(new_n867), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n831), .A2(new_n203), .B1(new_n842), .B2(new_n870), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT122), .Z(new_n1207));
  NOR2_X1   g1007(.A1(new_n834), .A2(new_n1007), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT53), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT54), .B(G143), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT121), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n879), .ZN(new_n1212));
  INV_X1    g1012(.A(G137), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1209), .B(new_n1212), .C1(new_n1213), .C2(new_n867), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G132), .A2(new_n837), .B1(new_n843), .B2(G125), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n340), .B1(new_n873), .B2(G128), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n832), .A2(G50), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n827), .A2(G159), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1205), .A2(new_n1207), .B1(new_n1214), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1201), .B1(new_n1220), .B2(new_n812), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1200), .A2(new_n1221), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1199), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1198), .A2(KEYINPUT123), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT123), .B1(new_n1198), .B2(new_n1223), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(G378));
  NAND2_X1  g1027(.A1(new_n987), .A2(new_n988), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n975), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(G330), .A3(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n473), .B1(new_n446), .B2(new_n727), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n446), .A2(new_n727), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n468), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1234), .B(new_n1236), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n950), .A2(new_n1237), .A3(new_n965), .A4(new_n967), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT108), .B1(new_n935), .B2(new_n961), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n947), .A2(new_n963), .A3(new_n948), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n966), .B1(new_n1241), .B2(new_n960), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1237), .B1(new_n1242), .B2(new_n950), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1230), .B1(new_n1238), .B2(new_n1243), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n737), .B(new_n975), .C1(new_n987), .C2(new_n988), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1237), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n968), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1242), .A2(new_n950), .A3(new_n1237), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n798), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n809), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n800), .B1(G50), .B2(new_n892), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n873), .A2(G125), .B1(new_n827), .B2(G150), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT124), .Z(new_n1254));
  NAND2_X1  g1054(.A1(new_n1211), .A2(new_n835), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n839), .A2(new_n884), .B1(new_n822), .B2(new_n1213), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G128), .B2(new_n837), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT59), .Z(new_n1259));
  NAND2_X1  g1059(.A1(new_n843), .A2(G124), .ZN(new_n1260));
  AOI211_X1 g1060(.A(G33), .B(G41), .C1(new_n832), .C2(G159), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(G41), .B(new_n342), .C1(new_n835), .C2(G77), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n832), .A2(G58), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n843), .A2(G283), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1263), .A2(new_n1013), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n818), .A2(new_n557), .B1(new_n822), .B2(new_n420), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n206), .A2(new_n839), .B1(new_n836), .B2(new_n207), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT58), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(KEYINPUT58), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n758), .B1(new_n253), .B2(new_n255), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n201), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1262), .A2(new_n1270), .A3(new_n1271), .A4(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1252), .B1(new_n1274), .B2(new_n812), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1251), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1250), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1197), .A2(new_n1179), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(KEYINPUT57), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n761), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT57), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1282), .B2(new_n1283), .ZN(G375));
  NOR2_X1   g1084(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1285), .A2(new_n1076), .A3(new_n1195), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT125), .Z(new_n1287));
  AOI22_X1  g1087(.A1(G283), .A2(new_n837), .B1(new_n843), .B2(G303), .ZN(new_n1288));
  AND4_X1   g1088(.A1(new_n340), .A2(new_n1288), .A3(new_n1010), .A4(new_n1109), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n822), .A2(new_n207), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n818), .A2(new_n870), .B1(new_n834), .B2(new_n206), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1290), .B(new_n1291), .C1(new_n868), .C2(G116), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(G159), .A2(new_n835), .B1(new_n879), .B2(G150), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n884), .B2(new_n818), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n868), .B2(new_n1211), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(G137), .A2(new_n837), .B1(new_n843), .B2(G128), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n342), .A3(new_n1264), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(G50), .B2(new_n827), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1289), .A2(new_n1292), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  OAI221_X1 g1099(.A(new_n800), .B1(G68), .B2(new_n892), .C1(new_n1299), .C2(new_n815), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n957), .B2(new_n809), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1176), .B2(new_n799), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1287), .A2(new_n1302), .ZN(G381));
  NOR3_X1   g1103(.A1(new_n1230), .A2(new_n1238), .A3(new_n1243), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1247), .A2(new_n1248), .B1(new_n989), .B2(G330), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n799), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1276), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1249), .A2(new_n1244), .B1(new_n1197), .B2(new_n1179), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n760), .B1(new_n1308), .B2(KEYINPUT57), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1283), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1307), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1198), .A2(new_n1223), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1098), .A2(new_n863), .A3(new_n1132), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1287), .A2(new_n907), .A3(new_n1302), .ZN(new_n1316));
  NOR4_X1   g1116(.A1(G390), .A2(new_n1314), .A3(new_n1315), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1093), .ZN(G407));
  NOR2_X1   g1118(.A1(new_n725), .A2(G343), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G407), .B(G213), .C1(new_n1314), .C2(new_n1320), .ZN(G409));
  NAND2_X1  g1121(.A1(G393), .A2(G396), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1315), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1142), .A2(new_n1323), .A3(new_n1165), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1142), .B2(new_n1165), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1076), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1074), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1073), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1052), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1326), .B1(new_n1329), .B2(new_n1036), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1091), .B1(new_n1330), .B2(new_n798), .ZN(new_n1331));
  OAI22_X1  g1131(.A1(new_n1324), .A2(new_n1325), .B1(new_n1331), .B2(new_n1035), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(G390), .A2(new_n1315), .A3(new_n1322), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1142), .A2(new_n1323), .A3(new_n1165), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1333), .A2(new_n1093), .A3(new_n1334), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1332), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1311), .A2(G378), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1306), .A2(KEYINPUT126), .A3(new_n1276), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT126), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(new_n1250), .B2(new_n1277), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1308), .A2(new_n1326), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1338), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1313), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1319), .B1(new_n1337), .B2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1285), .B1(KEYINPUT60), .B2(new_n1180), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1170), .A2(new_n1178), .A3(KEYINPUT60), .A4(new_n1175), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n761), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1302), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1348));
  OR2_X1    g1148(.A1(new_n1348), .A2(new_n907), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n907), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1344), .A2(KEYINPUT63), .A3(new_n1352), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1338), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT123), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1312), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1224), .ZN(new_n1357));
  OAI22_X1  g1157(.A1(new_n1354), .A2(new_n1312), .B1(G375), .B2(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1358), .A2(new_n1320), .A3(new_n1352), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT63), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(new_n1320), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1319), .A2(G2897), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1351), .B(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(KEYINPUT61), .B1(new_n1362), .B2(new_n1364), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1336), .A2(new_n1353), .A3(new_n1361), .A4(new_n1365), .ZN(new_n1366));
  AOI21_X1  g1166(.A(KEYINPUT62), .B1(new_n1344), .B2(new_n1352), .ZN(new_n1367));
  AOI22_X1  g1167(.A1(new_n1311), .A2(G378), .B1(new_n1342), .B2(new_n1313), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT62), .ZN(new_n1369));
  NOR4_X1   g1169(.A1(new_n1368), .A2(new_n1369), .A3(new_n1319), .A4(new_n1351), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1365), .B(KEYINPUT127), .C1(new_n1367), .C2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1332), .A2(new_n1335), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1359), .A2(new_n1369), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1344), .A2(KEYINPUT62), .A3(new_n1352), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  AOI21_X1  g1176(.A(KEYINPUT127), .B1(new_n1376), .B2(new_n1365), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1366), .B1(new_n1373), .B2(new_n1377), .ZN(G405));
  OAI21_X1  g1178(.A(new_n1337), .B1(new_n1312), .B2(new_n1311), .ZN(new_n1379));
  XNOR2_X1  g1179(.A(new_n1379), .B(new_n1352), .ZN(new_n1380));
  XNOR2_X1  g1180(.A(new_n1372), .B(new_n1380), .ZN(G402));
endmodule


