//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n216), .B2(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  AND2_X1   g0043(.A1(G1), .A2(G13), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n249), .B1(new_n250), .B2(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n246), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(new_n254), .B2(new_n253), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n244), .B2(new_n245), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT66), .B1(new_n258), .B2(new_n261), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n261), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(G226), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT69), .B(G179), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n203), .A2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(G150), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n214), .A2(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n272), .B1(new_n273), .B2(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n213), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n278), .A2(new_n280), .B1(new_n202), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n279), .A2(new_n213), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n282), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n283), .A2(new_n280), .A3(KEYINPUT68), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n284), .B1(new_n202), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n268), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n271), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n269), .A2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n256), .B2(new_n267), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n291), .B(KEYINPUT9), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n303), .A2(new_n296), .A3(new_n299), .A4(new_n300), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n295), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G68), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n283), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n309), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n250), .B2(new_n276), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n283), .A2(new_n280), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G68), .A3(new_n285), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n311), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT11), .B1(new_n313), .B2(new_n280), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G226), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n248), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n247), .B(new_n321), .C1(G232), .C2(new_n248), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n246), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n246), .A2(G274), .A3(new_n261), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT66), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n261), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT71), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n266), .A2(G238), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n330), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n325), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT13), .ZN(new_n336));
  INV_X1    g0136(.A(new_n332), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT71), .B1(new_n264), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n325), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n336), .A2(G190), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n336), .A2(new_n342), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT72), .B1(new_n344), .B2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT72), .ZN(new_n346));
  AOI211_X1 g0146(.A(new_n346), .B(new_n297), .C1(new_n336), .C2(new_n342), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n319), .B(new_n343), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n319), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n341), .B1(new_n340), .B2(new_n325), .ZN(new_n351));
  AOI211_X1 g0151(.A(KEYINPUT13), .B(new_n324), .C1(new_n338), .C2(new_n339), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(G169), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n336), .A2(G179), .A3(new_n342), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n350), .B1(new_n344), .B2(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n264), .B1(G244), .B2(new_n266), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n360));
  INV_X1    g0160(.A(G238), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n206), .B2(new_n247), .C1(new_n251), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n265), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G200), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n315), .A2(G77), .A3(new_n285), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G77), .B2(new_n282), .ZN(new_n367));
  INV_X1    g0167(.A(new_n277), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n276), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n367), .B1(new_n371), .B2(new_n280), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n365), .B(new_n372), .C1(new_n373), .C2(new_n364), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n364), .B2(new_n292), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n359), .A2(new_n270), .A3(new_n363), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n368), .A2(new_n283), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n315), .A2(new_n286), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT68), .B1(new_n283), .B2(new_n280), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n382), .A2(new_n383), .B1(new_n281), .B2(G20), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(new_n277), .ZN(new_n385));
  INV_X1    g0185(.A(G58), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n309), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n201), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n274), .A2(G159), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n391));
  INV_X1    g0191(.A(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G33), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n394), .A2(G33), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n214), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT16), .B(new_n390), .C1(new_n401), .C2(new_n309), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n280), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT73), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n393), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n400), .A2(G20), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n393), .B2(new_n404), .ZN(new_n407));
  AOI21_X1  g0207(.A(G20), .B1(new_n393), .B2(new_n395), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n405), .A2(new_n407), .B1(new_n408), .B2(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT16), .B1(new_n410), .B2(new_n390), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n385), .B1(new_n403), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n320), .A2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G223), .B2(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n393), .A2(new_n395), .ZN(new_n415));
  INV_X1    g0215(.A(G87), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n414), .A2(new_n415), .B1(new_n392), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n265), .B1(G232), .B2(new_n266), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n330), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(G190), .A3(new_n330), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n379), .B1(new_n412), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n380), .B1(new_n290), .B2(new_n368), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n388), .A2(new_n389), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n408), .A2(KEYINPUT7), .B1(new_n247), .B2(new_n391), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(G68), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n287), .B1(new_n427), .B2(KEYINPUT16), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT16), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n397), .A2(KEYINPUT73), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n406), .C1(new_n415), .C2(KEYINPUT73), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n400), .B1(new_n247), .B2(G20), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n309), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n429), .B1(new_n433), .B2(new_n425), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n424), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n417), .A2(new_n265), .ZN(new_n436));
  INV_X1    g0236(.A(new_n270), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n266), .A2(G232), .ZN(new_n438));
  AND4_X1   g0238(.A1(new_n330), .A2(new_n436), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n292), .B1(new_n418), .B2(new_n330), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT18), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n419), .A2(G169), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n418), .A2(new_n330), .A3(new_n437), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n412), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n418), .A2(G190), .A3(new_n330), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n297), .B1(new_n418), .B2(new_n330), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n435), .A2(new_n450), .A3(KEYINPUT17), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n423), .A2(new_n442), .A3(new_n447), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n378), .B1(new_n453), .B2(KEYINPUT74), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(KEYINPUT74), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n308), .A2(new_n358), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n393), .A2(new_n395), .A3(new_n214), .A4(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(KEYINPUT80), .A2(KEYINPUT22), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT81), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G116), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G20), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT23), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n214), .B2(G107), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n460), .B1(KEYINPUT81), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n462), .B(new_n468), .C1(new_n458), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT24), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n470), .A2(new_n458), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n462), .A4(new_n468), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n280), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT25), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n282), .B2(G107), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n282), .A2(new_n478), .A3(G107), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n281), .A2(G33), .ZN(new_n482));
  AND4_X1   g0282(.A1(new_n213), .A2(new_n282), .A3(new_n279), .A4(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n479), .A2(new_n481), .B1(new_n483), .B2(G107), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G257), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G1698), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G250), .B2(G1698), .ZN(new_n488));
  INV_X1    g0288(.A(G294), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n488), .A2(new_n415), .B1(new_n392), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n265), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n260), .A2(G1), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G264), .A3(new_n246), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n258), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n495), .A2(KEYINPUT82), .A3(G264), .A4(new_n246), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n491), .A2(new_n498), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n265), .A2(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(KEYINPUT83), .A3(new_n500), .A4(new_n501), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n506), .A3(G169), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n504), .A2(new_n506), .A3(new_n509), .A4(G169), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n491), .A2(new_n498), .A3(new_n501), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G179), .A3(new_n500), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n485), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NOR2_X1   g0315(.A1(G257), .A2(G1698), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n248), .A2(G264), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n247), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g0318(.A(KEYINPUT79), .B(G303), .Z(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n265), .C1(new_n247), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n495), .A2(G270), .A3(new_n246), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n500), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n283), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n287), .A2(new_n282), .A3(new_n482), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n524), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(KEYINPUT75), .A2(G33), .A3(G283), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(G20), .B1(new_n392), .B2(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n279), .A2(new_n213), .B1(G20), .B2(new_n524), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT20), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n535), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n527), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n515), .B1(new_n523), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n483), .A2(G116), .ZN(new_n541));
  INV_X1    g0341(.A(new_n538), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n525), .B(new_n541), .C1(new_n542), .C2(new_n536), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n543), .A2(KEYINPUT21), .A3(G169), .A4(new_n522), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n522), .A2(G200), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n520), .A2(G190), .A3(new_n500), .A4(new_n521), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  AND4_X1   g0347(.A1(G179), .A2(new_n520), .A3(new_n500), .A4(new_n521), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n543), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n540), .A2(new_n544), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n247), .A2(G244), .A3(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n393), .A2(new_n395), .A3(G238), .A4(new_n248), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n463), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n265), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n258), .A2(KEYINPUT77), .A3(new_n492), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n246), .A2(G274), .A3(new_n492), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT77), .ZN(new_n557));
  INV_X1    g0357(.A(G250), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n492), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n556), .A2(new_n557), .B1(new_n559), .B2(new_n246), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n292), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n554), .A2(new_n270), .A3(new_n555), .A4(new_n560), .ZN(new_n563));
  INV_X1    g0363(.A(new_n370), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n282), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n247), .A2(new_n214), .A3(G68), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n214), .B1(new_n323), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G87), .B2(new_n207), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n276), .B2(new_n205), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n565), .B1(new_n571), .B2(new_n280), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT78), .B1(new_n526), .B2(new_n370), .ZN(new_n573));
  OR3_X1    g0373(.A1(new_n526), .A2(KEYINPUT78), .A3(new_n370), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n562), .A2(new_n563), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n553), .A2(new_n265), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n556), .A2(new_n557), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n559), .A2(new_n246), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n555), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(G200), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  AOI221_X4 g0381(.A(new_n565), .B1(G87), .B2(new_n483), .C1(new_n571), .C2(new_n280), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n554), .A2(G190), .A3(new_n555), .A4(new_n560), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n550), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT6), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n587), .A2(new_n205), .A3(G107), .ZN(new_n588));
  XNOR2_X1  g0388(.A(G97), .B(G107), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n590), .A2(new_n214), .B1(new_n250), .B2(new_n275), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n206), .B1(new_n431), .B2(new_n432), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n280), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n282), .A2(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n483), .B2(G97), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n495), .A2(new_n246), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n500), .B1(new_n597), .B2(new_n486), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n393), .A2(new_n395), .A3(G244), .A4(new_n248), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT4), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n532), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n598), .B1(new_n604), .B2(new_n265), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(G190), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n598), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n604), .A2(KEYINPUT76), .A3(new_n265), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT76), .B1(new_n604), .B2(new_n265), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G200), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n270), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n604), .A2(new_n265), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n292), .A2(new_n614), .B1(new_n593), .B2(new_n595), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n606), .A2(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n504), .A2(new_n506), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n373), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n502), .A2(new_n297), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n485), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n514), .A2(new_n586), .A3(new_n616), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n457), .A2(new_n623), .ZN(G372));
  NAND2_X1  g0424(.A1(new_n423), .A2(new_n451), .ZN(new_n625));
  INV_X1    g0425(.A(new_n377), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n348), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n627), .B2(new_n357), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n442), .A2(new_n447), .ZN(new_n630));
  OR3_X1    g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n305), .A2(new_n306), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n628), .B2(new_n630), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n615), .A2(new_n612), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT26), .B1(new_n635), .B2(new_n585), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n580), .A2(KEYINPUT85), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n560), .A2(new_n638), .A3(new_n555), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n577), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n563), .B(new_n575), .C1(new_n640), .C2(G169), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n583), .B(new_n582), .C1(new_n640), .C2(new_n297), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(new_n612), .A4(new_n615), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n636), .B(new_n641), .C1(KEYINPUT26), .C2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n485), .B1(new_n618), .B2(new_n619), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n642), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n510), .A2(new_n512), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n621), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n544), .A2(new_n549), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n540), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n647), .B(new_n616), .C1(new_n650), .C2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n644), .B1(new_n653), .B2(KEYINPUT86), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n606), .A2(new_n611), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n635), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n656), .A2(new_n645), .A3(new_n646), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT86), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(new_n650), .C2(new_n652), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n456), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n634), .A2(new_n294), .A3(new_n661), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n281), .A2(new_n214), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n539), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n652), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n550), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT88), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n650), .A2(new_n677), .A3(new_n668), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT89), .B1(new_n514), .B2(new_n669), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n649), .A2(new_n512), .A3(new_n510), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n645), .B1(new_n485), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n485), .A2(new_n668), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n678), .A2(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n514), .A2(new_n668), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n677), .B1(new_n650), .B2(new_n668), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n514), .A2(KEYINPUT89), .A3(new_n669), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n652), .A2(new_n669), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n685), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n210), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n218), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT91), .B1(new_n623), .B2(new_n668), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n586), .A2(new_n616), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT91), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n681), .A4(new_n669), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n561), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n548), .A3(new_n511), .A4(new_n605), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT90), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(KEYINPUT90), .A3(new_n709), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n707), .A2(new_n511), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n605), .A4(new_n548), .ZN(new_n715));
  INV_X1    g0515(.A(new_n640), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n502), .A2(new_n270), .A3(new_n522), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n610), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n712), .A2(new_n713), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT31), .B1(new_n719), .B2(new_n668), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n715), .A2(new_n710), .A3(new_n718), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n668), .A2(KEYINPUT31), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n706), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT26), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n635), .B2(new_n585), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n727), .B(new_n728), .C1(new_n726), .C2(new_n643), .ZN(new_n729));
  INV_X1    g0529(.A(new_n646), .ZN(new_n730));
  INV_X1    g0530(.A(new_n635), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n729), .A2(new_n641), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT93), .B1(new_n650), .B2(new_n652), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n651), .A2(new_n540), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n514), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n657), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n668), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(KEYINPUT29), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT29), .B1(new_n660), .B2(new_n669), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n725), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n701), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n675), .A2(G330), .ZN(new_n745));
  INV_X1    g0545(.A(new_n673), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n674), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n673), .A2(KEYINPUT88), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n747), .A2(G330), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n214), .A2(G13), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n281), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n696), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n745), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n746), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n213), .B1(G20), .B2(new_n292), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n695), .A2(new_n415), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n210), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n695), .A2(new_n247), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G45), .B2(new_n218), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n242), .B2(G45), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n760), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n753), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n214), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT96), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n416), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n770), .A2(new_n373), .A3(new_n297), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n214), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G97), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(new_n373), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n206), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n415), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n780), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n437), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n373), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G200), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n776), .B(new_n788), .C1(new_n792), .C2(G77), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n297), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n790), .A2(G190), .A3(new_n297), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G68), .A2(new_n794), .B1(new_n796), .B2(G58), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n793), .B(new_n797), .C1(new_n202), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n777), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n247), .B1(new_n800), .B2(G329), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n785), .ZN(new_n803));
  INV_X1    g0603(.A(new_n792), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n775), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n803), .B(new_n806), .C1(G303), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  INV_X1    g0609(.A(new_n794), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(new_n809), .B2(new_n795), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n798), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G326), .B1(G294), .B2(new_n783), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT97), .Z(new_n815));
  OAI21_X1  g0615(.A(new_n799), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n769), .B1(new_n816), .B2(new_n759), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n754), .B1(new_n758), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n378), .A2(new_n669), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n654), .B2(new_n659), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n660), .A2(new_n669), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n374), .B1(new_n372), .B2(new_n669), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n377), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n626), .A2(new_n669), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n822), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n753), .B1(new_n830), .B2(new_n725), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n725), .B2(new_n830), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n794), .A2(KEYINPUT98), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n794), .A2(KEYINPUT98), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G283), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n796), .A2(G294), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n247), .B1(new_n800), .B2(G311), .ZN(new_n839));
  INV_X1    g0639(.A(new_n785), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G87), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n839), .A2(new_n784), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G107), .B2(new_n807), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G116), .A2(new_n792), .B1(new_n813), .B2(G303), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n837), .A2(new_n838), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G159), .A2(new_n792), .B1(new_n796), .B2(G143), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n798), .C1(new_n273), .C2(new_n810), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT99), .Z(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n415), .B1(new_n800), .B2(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n309), .B2(new_n785), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G58), .B2(new_n783), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n850), .B(new_n853), .C1(new_n202), .C2(new_n775), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n845), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n759), .ZN(new_n857));
  INV_X1    g0657(.A(new_n753), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n759), .A2(new_n755), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n250), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n829), .B2(new_n756), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n832), .B1(new_n857), .B2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(new_n590), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n524), .B(new_n216), .C1(new_n863), .C2(KEYINPUT35), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(KEYINPUT35), .B2(new_n863), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT36), .Z(new_n866));
  OR3_X1    g0666(.A1(new_n218), .A2(new_n250), .A3(new_n387), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n202), .A2(G68), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n281), .B(G13), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n630), .A2(new_n666), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n412), .A2(new_n445), .ZN(new_n873));
  INV_X1    g0673(.A(new_n666), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n412), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n428), .A2(new_n434), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n876), .A2(new_n385), .A3(new_n421), .A4(new_n420), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n873), .A2(new_n875), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n390), .B1(new_n401), .B2(new_n309), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n429), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n424), .B1(new_n428), .B2(new_n881), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n412), .A2(new_n422), .B1(new_n882), .B2(new_n441), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n666), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n879), .A2(new_n885), .B1(new_n452), .B2(new_n884), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT39), .B1(new_n886), .B2(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT101), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n873), .A2(new_n875), .A3(new_n877), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n879), .ZN(new_n891));
  INV_X1    g0691(.A(new_n875), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n452), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n888), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI211_X1 g0697(.A(KEYINPUT101), .B(new_n895), .C1(new_n891), .C2(new_n893), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n887), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n885), .A2(new_n879), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n452), .A2(new_n884), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(G169), .B1(new_n351), .B2(new_n352), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT14), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n354), .A3(new_n353), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n349), .A3(new_n669), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n872), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n343), .A2(new_n319), .ZN(new_n915));
  OAI21_X1  g0715(.A(G200), .B1(new_n351), .B2(new_n352), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n346), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n344), .A2(KEYINPUT72), .A3(G200), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n349), .B(new_n668), .C1(new_n919), .C2(new_n911), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n349), .A2(new_n668), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n348), .A2(new_n357), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n827), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n906), .B(new_n923), .C1(new_n821), .C2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT102), .B1(new_n914), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n905), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n894), .A2(new_n888), .A3(new_n896), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n890), .A2(new_n879), .B1(new_n452), .B2(new_n892), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT101), .B1(new_n930), .B2(new_n895), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n928), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n927), .B1(new_n904), .B2(new_n905), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n913), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND4_X1   g0734(.A1(KEYINPUT102), .A2(new_n925), .A3(new_n934), .A4(new_n871), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n741), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n739), .A2(KEYINPUT29), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(new_n456), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n634), .A3(new_n294), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n936), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n828), .B1(new_n920), .B2(new_n922), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n720), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n706), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n945), .A3(new_n906), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n905), .B1(new_n897), .B2(new_n898), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n949), .A2(KEYINPUT40), .A3(new_n945), .A4(new_n942), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n456), .A3(new_n945), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(G330), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n951), .B1(new_n456), .B2(new_n945), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n281), .B2(new_n750), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n941), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n870), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT103), .ZN(G367));
  NAND2_X1  g0760(.A1(new_n836), .A2(G159), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n783), .A2(G68), .ZN(new_n962));
  INV_X1    g0762(.A(G143), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n962), .B1(new_n798), .B2(new_n963), .C1(new_n273), .C2(new_n795), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT106), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n964), .A2(KEYINPUT106), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n840), .A2(G77), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n415), .B1(new_n800), .B2(G137), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n775), .C2(new_n386), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n792), .B2(G50), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n961), .A2(new_n965), .A3(new_n966), .A4(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n519), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n804), .A2(new_n802), .B1(new_n972), .B2(new_n795), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G311), .B2(new_n813), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n807), .A2(KEYINPUT46), .A3(G116), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT46), .B1(new_n807), .B2(G116), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n782), .A2(new_n206), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n415), .B1(new_n777), .B2(new_n978), .C1(new_n205), .C2(new_n785), .ZN(new_n979));
  NOR4_X1   g0779(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n974), .B(new_n980), .C1(new_n835), .C2(new_n489), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n971), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT47), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT47), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n759), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n760), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n695), .B2(new_n564), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n230), .A2(new_n765), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n858), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n757), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n582), .A2(new_n669), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n730), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n641), .B2(new_n991), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n985), .B(new_n989), .C1(new_n990), .C2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n669), .B1(new_n593), .B2(new_n595), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n656), .A2(new_n996), .B1(new_n635), .B2(new_n669), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n995), .B1(new_n693), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n678), .A2(new_n679), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n691), .B1(new_n1000), .B2(new_n687), .ZN(new_n1001));
  OAI211_X1 g0801(.A(KEYINPUT44), .B(new_n999), .C1(new_n1001), .C2(new_n686), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n686), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1005), .B(new_n997), .C1(new_n683), .C2(new_n691), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n684), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n683), .A2(new_n691), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n676), .B1(new_n1013), .B2(new_n1001), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n690), .A2(new_n692), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n749), .A2(new_n1015), .A3(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n742), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1003), .A2(new_n685), .A3(new_n1009), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1011), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n743), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n696), .B(KEYINPUT41), .Z(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n752), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT104), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n514), .B1(new_n611), .B2(new_n606), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n669), .B1(new_n1026), .B2(new_n731), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT42), .B1(new_n1001), .B2(new_n997), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT42), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n683), .A2(new_n1029), .A3(new_n999), .A4(new_n691), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1027), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1025), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1029), .B1(new_n1015), .B2(new_n999), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1001), .A2(KEYINPUT42), .A3(new_n997), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1036), .A2(KEYINPUT104), .A3(new_n1037), .A4(new_n1027), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n993), .B(KEYINPUT43), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1033), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n997), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n684), .A2(new_n997), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT105), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1041), .A2(new_n1045), .A3(new_n1044), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n994), .B1(new_n1024), .B2(new_n1049), .ZN(G387));
  OAI21_X1  g0850(.A(KEYINPUT107), .B1(new_n1017), .B2(new_n751), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1017), .A2(KEYINPUT107), .A3(new_n751), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n765), .B1(new_n235), .B2(new_n260), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n698), .B2(new_n762), .ZN(new_n1054));
  OR3_X1    g0854(.A1(new_n277), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1055));
  OAI21_X1  g0855(.A(KEYINPUT50), .B1(new_n277), .B2(G50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1055), .A2(new_n698), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1054), .A2(new_n1058), .B1(new_n206), .B2(new_n695), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n753), .B1(new_n1059), .B2(new_n986), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n783), .A2(new_n564), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n795), .B2(new_n202), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT109), .Z(new_n1063));
  NAND2_X1  g0863(.A1(new_n807), .A2(G77), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT108), .B(G150), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n415), .B1(new_n800), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(new_n205), .C2(new_n785), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n794), .B2(new_n368), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G68), .A2(new_n792), .B1(new_n813), .B2(G159), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1063), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n796), .B1(new_n813), .B2(G322), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n972), .B2(new_n804), .C1(new_n835), .C2(new_n805), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n775), .A2(new_n489), .B1(new_n802), .B2(new_n782), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT110), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n247), .B1(new_n800), .B2(G326), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n524), .C2(new_n785), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT49), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1070), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1060), .B1(new_n1082), .B2(new_n759), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n683), .A2(new_n757), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1051), .A2(new_n1052), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n937), .A2(new_n938), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1086), .A2(new_n725), .A3(new_n1016), .A4(new_n1014), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n742), .A2(new_n1017), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n696), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1085), .A2(new_n1089), .ZN(G393));
  AND3_X1   g0890(.A1(new_n1003), .A2(new_n685), .A3(new_n1009), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n685), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n999), .A2(new_n757), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n760), .B1(new_n205), .B2(new_n210), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n239), .B2(new_n765), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n273), .A2(new_n798), .B1(new_n795), .B2(new_n778), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n247), .B1(new_n777), .B2(new_n963), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G87), .B2(new_n840), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n250), .B2(new_n782), .C1(new_n309), .C2(new_n775), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n792), .B2(new_n368), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1098), .B(new_n1102), .C1(new_n202), .C2(new_n835), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n247), .B(new_n786), .C1(G116), .C2(new_n783), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n775), .A2(new_n802), .B1(new_n809), .B2(new_n777), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT111), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n804), .A2(new_n489), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n1106), .C2(new_n1105), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n972), .B2(new_n835), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n805), .A2(new_n795), .B1(new_n798), .B2(new_n978), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT52), .Z(new_n1112));
  OAI21_X1  g0912(.A(new_n1103), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n858), .B(new_n1096), .C1(new_n1113), .C2(new_n759), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1093), .A2(new_n752), .B1(new_n1094), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1087), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n1020), .A3(new_n696), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT112), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT112), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(G390));
  INV_X1    g0921(.A(new_n826), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n668), .B(new_n1122), .C1(new_n733), .C2(new_n738), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n923), .B1(new_n1123), .B2(new_n924), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT113), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n949), .A2(new_n912), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n920), .A2(new_n922), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n650), .A2(KEYINPUT93), .A3(new_n652), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n736), .B1(new_n514), .B2(new_n735), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n616), .A2(new_n730), .A3(new_n622), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n729), .A2(new_n641), .A3(new_n732), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n669), .B(new_n826), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1128), .B1(new_n1134), .B2(new_n827), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n949), .A2(new_n912), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT113), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n908), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n821), .A2(new_n924), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n912), .B1(new_n1139), .B2(new_n1128), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1127), .A2(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n945), .A2(G330), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n942), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1140), .A2(new_n1138), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n724), .A2(G330), .A3(new_n829), .A4(new_n923), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1125), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1135), .A2(new_n1136), .A3(KEYINPUT113), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1146), .B(new_n1147), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1143), .A2(new_n456), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n939), .A2(new_n634), .A3(new_n294), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1128), .B1(new_n1142), .B2(new_n828), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1156), .A2(new_n827), .A3(new_n1134), .A4(new_n1147), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n724), .A2(G330), .A3(new_n829), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1143), .A2(new_n942), .B1(new_n1158), .B2(new_n1128), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1139), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT114), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1152), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(KEYINPUT114), .B(new_n1161), .C1(new_n1145), .C2(new_n1151), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n696), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n804), .A2(new_n205), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n798), .A2(new_n802), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n415), .B1(new_n777), .B2(new_n489), .C1(new_n309), .C2(new_n785), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n776), .A4(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n795), .A2(new_n524), .B1(new_n250), .B2(new_n782), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT116), .Z(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n206), .C2(new_n835), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n813), .A2(G128), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n804), .A2(new_n1174), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G132), .C2(new_n796), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n807), .A2(new_n1065), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1177), .A2(KEYINPUT53), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(KEYINPUT53), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n782), .A2(new_n778), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n415), .B1(new_n800), .B2(G125), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n202), .B2(new_n785), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1176), .B(new_n1183), .C1(new_n847), .C2(new_n835), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1172), .B1(new_n1185), .B2(KEYINPUT115), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT115), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n759), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n858), .B1(new_n277), .B2(new_n859), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n908), .C2(new_n756), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1152), .B2(new_n752), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1165), .A2(new_n1193), .ZN(G378));
  OAI21_X1  g0994(.A(KEYINPUT119), .B1(new_n926), .B2(new_n935), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n925), .A2(new_n934), .A3(new_n871), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT102), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n914), .A2(KEYINPUT102), .A3(new_n925), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT119), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n948), .A2(G330), .A3(new_n950), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n291), .A2(new_n874), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT118), .Z(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n307), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1208));
  NAND2_X1  g1008(.A1(new_n307), .A2(new_n1205), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1208), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1204), .B(new_n295), .C1(new_n305), .C2(new_n306), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1202), .A2(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(G330), .A3(new_n948), .A4(new_n950), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1195), .A2(new_n1201), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT120), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1215), .B(new_n1217), .C1(new_n926), .C2(new_n935), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1195), .A2(new_n1218), .A3(new_n1201), .A4(KEYINPUT120), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1150), .B(new_n1160), .C1(new_n1141), .C2(new_n1144), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1155), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT121), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1226), .A2(KEYINPUT121), .A3(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1218), .A2(new_n936), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1227), .B1(new_n1232), .B2(new_n1221), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1225), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n696), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(new_n1231), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1222), .A2(new_n752), .A3(new_n1223), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G33), .A2(G41), .ZN(new_n1239));
  AOI211_X1 g1039(.A(G50), .B(new_n1239), .C1(new_n415), .C2(new_n259), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G97), .A2(new_n794), .B1(new_n796), .B2(G107), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n840), .A2(G58), .ZN(new_n1242));
  AOI211_X1 g1042(.A(G41), .B(new_n247), .C1(new_n800), .C2(G283), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1064), .A2(new_n962), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n792), .B2(new_n564), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1241), .B(new_n1245), .C1(new_n524), .C2(new_n798), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT58), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1240), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n775), .A2(new_n1174), .B1(new_n273), .B2(new_n782), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G125), .A2(new_n813), .B1(new_n796), .B2(G128), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n792), .A2(G137), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1249), .B(new_n1252), .C1(G132), .C2(new_n794), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT59), .ZN(new_n1255));
  INV_X1    g1055(.A(G124), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1239), .B1(new_n777), .B2(new_n1256), .C1(new_n778), .C2(new_n785), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT117), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT59), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1258), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1248), .B1(new_n1247), .B2(new_n1246), .C1(new_n1255), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n759), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n858), .B1(new_n202), .B2(new_n859), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n1216), .C2(new_n756), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1238), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1237), .A2(new_n1266), .ZN(G375));
  OR2_X1    g1067(.A1(new_n1159), .A2(new_n1139), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1161), .A2(new_n1269), .A3(new_n1023), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1128), .A2(new_n755), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n858), .B1(new_n309), .B2(new_n859), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT122), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n835), .A2(new_n1174), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G150), .A2(new_n792), .B1(new_n813), .B2(G132), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n415), .B1(new_n800), .B2(G128), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1276), .B(new_n1242), .C1(new_n202), .C2(new_n782), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G159), .B2(new_n807), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1275), .B(new_n1278), .C1(new_n847), .C2(new_n795), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n835), .A2(new_n524), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G283), .A2(new_n796), .B1(new_n813), .B2(G294), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n247), .B1(new_n800), .B2(G303), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1061), .A3(new_n967), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G97), .B2(new_n807), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1281), .B(new_n1284), .C1(new_n206), .C2(new_n804), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1274), .A2(new_n1279), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1273), .B1(new_n1286), .B2(new_n759), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1160), .A2(new_n752), .B1(new_n1271), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1270), .A2(new_n1288), .ZN(G381));
  AOI21_X1  g1089(.A(new_n1235), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1265), .B1(new_n1290), .B2(new_n1231), .ZN(new_n1291));
  INV_X1    g1091(.A(G378), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NOR4_X1   g1093(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1022), .B1(new_n1020), .B2(new_n743), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1047), .B(new_n1048), .C1(new_n1295), .C2(new_n752), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1294), .A2(new_n994), .A3(new_n1296), .A4(new_n1120), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT123), .ZN(G407));
  INV_X1    g1099(.A(new_n1293), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n667), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G407), .A2(G213), .A3(new_n1301), .ZN(G409));
  OAI211_X1 g1102(.A(new_n994), .B(new_n1296), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT126), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(G393), .B(G396), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1119), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT112), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(G387), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1304), .A2(new_n1305), .B1(new_n1303), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  AND4_X1   g1110(.A1(new_n1310), .A2(new_n1308), .A3(new_n1305), .A4(new_n1303), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1232), .A2(new_n1221), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n752), .ZN(new_n1314));
  AND4_X1   g1114(.A1(new_n1165), .A2(new_n1193), .A3(new_n1264), .A4(new_n1314), .ZN(new_n1315));
  OR2_X1    g1115(.A1(new_n1226), .A2(new_n1022), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n1315), .A2(new_n1316), .B1(G213), .B2(new_n667), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1268), .A2(KEYINPUT60), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1319), .B(new_n1320), .ZN(new_n1321));
  XOR2_X1   g1121(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n1322));
  NAND2_X1  g1122(.A1(new_n1269), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(new_n696), .A3(new_n1161), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1288), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(G384), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G384), .B(new_n1288), .C1(new_n1321), .C2(new_n1324), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n667), .A2(G213), .A3(G2897), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AOI211_X1 g1132(.A(KEYINPUT61), .B(new_n1312), .C1(new_n1318), .C2(new_n1332), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1317), .B(new_n1334), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1292), .B1(new_n1237), .B2(new_n1266), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n667), .A2(G213), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1344), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1334), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1333), .A2(new_n1337), .A3(new_n1339), .A4(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1335), .A2(KEYINPUT62), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1226), .A2(KEYINPUT121), .A3(new_n1227), .ZN(new_n1348));
  AOI21_X1  g1148(.A(KEYINPUT121), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1348), .A2(new_n1349), .A3(new_n1235), .ZN(new_n1350));
  OAI21_X1  g1150(.A(G378), .B1(new_n1350), .B2(new_n1265), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT62), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1351), .A2(new_n1352), .A3(new_n1317), .A4(new_n1334), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT61), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1332), .B1(new_n1340), .B2(new_n1343), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1347), .A2(new_n1353), .A3(new_n1354), .A4(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1312), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1346), .A2(new_n1357), .ZN(G405));
  OAI21_X1  g1158(.A(new_n1312), .B1(new_n1300), .B2(new_n1340), .ZN(new_n1359));
  OAI211_X1 g1159(.A(new_n1351), .B(new_n1293), .C1(new_n1311), .C2(new_n1309), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1334), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1359), .A2(new_n1334), .A3(new_n1360), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(G402));
endmodule


