//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n966, new_n967;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(G43gat), .A2(G50gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G43gat), .A2(G50gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(new_n208), .A3(KEYINPUT14), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT15), .B(new_n207), .C1(new_n211), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n213), .A2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(new_n206), .ZN(new_n219));
  NOR2_X1   g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT15), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n210), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n223));
  OAI21_X1  g022(.A(G36gat), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n205), .A2(new_n225), .A3(new_n206), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n218), .A2(new_n221), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT16), .ZN(new_n232));
  INV_X1    g031(.A(G15gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(G22gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G15gat), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(G1gat), .B1(new_n234), .B2(new_n236), .ZN(new_n238));
  OAI21_X1  g037(.A(G8gat), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n240));
  INV_X1    g039(.A(G8gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(G15gat), .B(G22gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n240), .B(new_n241), .C1(G1gat), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n217), .A2(new_n227), .A3(KEYINPUT17), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT90), .B1(new_n228), .B2(new_n244), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n230), .A2(KEYINPUT90), .A3(new_n245), .A4(new_n246), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n204), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n202), .B1(new_n251), .B2(KEYINPUT18), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n217), .A2(new_n227), .A3(KEYINPUT17), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT17), .B1(new_n217), .B2(new_n227), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(new_n244), .ZN(new_n255));
  INV_X1    g054(.A(new_n248), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n203), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT18), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT91), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n228), .B(new_n244), .Z(new_n261));
  XOR2_X1   g060(.A(new_n203), .B(KEYINPUT13), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n251), .B2(KEYINPUT18), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G141gat), .ZN(new_n266));
  INV_X1    g065(.A(G197gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT11), .B(G169gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  NAND4_X1  g071(.A1(new_n252), .A2(new_n260), .A3(new_n265), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n272), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n257), .A2(KEYINPUT18), .A3(new_n203), .ZN(new_n275));
  INV_X1    g074(.A(new_n264), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n251), .A2(KEYINPUT18), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G15gat), .B(G43gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(new_n291), .B2(new_n289), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n287), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n302), .B(KEYINPUT28), .Z(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n295), .A2(KEYINPUT26), .A3(new_n304), .ZN(new_n305));
  AOI211_X1 g104(.A(new_n289), .B(new_n305), .C1(KEYINPUT26), .C2(new_n304), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G113gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G120gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT66), .B(G113gat), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n315), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n313), .A2(G113gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n310), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G227gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n299), .A2(new_n307), .A3(new_n326), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n284), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(KEYINPUT32), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n333), .B(KEYINPUT32), .C1(new_n334), .C2(new_n284), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n328), .A2(new_n332), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT34), .B1(new_n341), .B2(new_n331), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT34), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n343), .C1(new_n329), .C2(new_n330), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n337), .A2(new_n342), .A3(new_n344), .A4(new_n338), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n351), .A3(new_n347), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT36), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n339), .A2(KEYINPUT68), .A3(new_n345), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G155gat), .B(G162gat), .Z(new_n357));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT73), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(G141gat), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT73), .A3(G148gat), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n362), .B(new_n364), .C1(new_n363), .C2(G148gat), .ZN(new_n365));
  INV_X1    g164(.A(G155gat), .ZN(new_n366));
  INV_X1    g165(.A(G162gat), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT2), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G155gat), .B(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT74), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n359), .A2(new_n365), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G141gat), .B(G148gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n357), .B1(KEYINPUT2), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G211gat), .B(G218gat), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G218gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n382), .A2(KEYINPUT69), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(KEYINPUT69), .B2(new_n382), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n382), .A2(new_n387), .A3(new_n390), .A4(new_n386), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n386), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT70), .B1(new_n392), .B2(new_n381), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n376), .A2(KEYINPUT81), .A3(new_n377), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n375), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n371), .A2(new_n373), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n391), .A2(new_n393), .B1(new_n381), .B2(new_n392), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n404));
  OR3_X1    g203(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT29), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n403), .B2(KEYINPUT29), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n375), .A3(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n407), .A2(new_n400), .B1(new_n395), .B2(new_n378), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n408), .B2(new_n398), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT82), .B1(new_n409), .B2(G22gat), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n402), .B(new_n235), .C1(new_n408), .C2(new_n398), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT31), .B(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(KEYINPUT82), .A3(G22gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n409), .A2(G22gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n411), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n414), .B(KEYINPUT79), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n416), .A2(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G1gat), .B(G29gat), .Z(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n327), .A2(new_n427), .A3(new_n374), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n374), .A2(new_n320), .A3(new_n325), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT4), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n430), .A3(KEYINPUT78), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n376), .A2(new_n326), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n434), .A3(KEYINPUT4), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT39), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n426), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n326), .A2(new_n400), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n429), .A3(new_n437), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT39), .B1(new_n443), .B2(new_n444), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  OR3_X1    g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n447), .B1(new_n445), .B2(new_n446), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n436), .A2(new_n438), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n441), .A2(new_n451), .A3(KEYINPUT40), .ZN(new_n452));
  INV_X1    g251(.A(new_n395), .ZN(new_n453));
  NAND2_X1  g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n454), .B(KEYINPUT71), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n308), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n299), .A2(new_n307), .A3(KEYINPUT72), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n455), .A2(KEYINPUT29), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n308), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n453), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n299), .A2(new_n307), .A3(new_n455), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n395), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G8gat), .B(G36gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G64gat), .B(G92gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n464), .A2(new_n467), .A3(new_n471), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n433), .A2(new_n437), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n428), .A2(new_n430), .A3(KEYINPUT75), .ZN(new_n477));
  OR3_X1    g276(.A1(new_n429), .A2(KEYINPUT75), .A3(KEYINPUT4), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n480));
  NAND2_X1  g279(.A1(new_n442), .A2(new_n429), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n438), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n476), .A2(new_n431), .A3(new_n480), .A4(new_n435), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n426), .ZN(new_n486));
  OR3_X1    g285(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n472), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n452), .A2(new_n475), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT40), .B1(new_n441), .B2(new_n451), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n421), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n464), .A2(new_n493), .A3(new_n467), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n395), .B1(new_n460), .B2(new_n463), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n465), .A2(new_n453), .A3(new_n466), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT37), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n471), .A2(KEYINPUT38), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n474), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n468), .A2(KEYINPUT37), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n472), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n493), .B1(new_n464), .B2(new_n467), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT86), .B1(new_n504), .B2(new_n471), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n505), .A3(new_n494), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n500), .B1(new_n506), .B2(KEYINPUT38), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508));
  INV_X1    g307(.A(new_n426), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n483), .A2(new_n509), .A3(new_n484), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n486), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n483), .B2(new_n484), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n507), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n356), .B1(new_n492), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n511), .A2(new_n513), .B1(new_n475), .B2(new_n487), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT82), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n418), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n411), .A2(new_n414), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n417), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n419), .A2(new_n420), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n519), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n475), .A2(new_n487), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n421), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n517), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n352), .A2(new_n354), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT87), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n352), .A2(new_n537), .A3(new_n354), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n526), .A2(new_n349), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n514), .A2(new_n530), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n281), .B1(new_n529), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G57gat), .B(G64gat), .Z(new_n545));
  NAND2_X1  g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT92), .A3(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n546), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n552), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(new_n545), .A3(KEYINPUT92), .A4(new_n548), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(KEYINPUT21), .ZN(new_n559));
  XOR2_X1   g358(.A(G127gat), .B(G155gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n244), .B1(new_n558), .B2(KEYINPUT21), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT93), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT94), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n563), .B(new_n570), .Z(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT95), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT7), .ZN(new_n579));
  AND2_X1   g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n577), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n575), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G99gat), .B(G106gat), .Z(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n586), .B(new_n575), .C1(new_n581), .C2(new_n582), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(KEYINPUT96), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n589), .A3(new_n584), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n588), .A2(new_n230), .A3(new_n246), .A4(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n253), .A2(new_n254), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n594), .A2(KEYINPUT97), .A3(new_n590), .A4(new_n588), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n588), .A2(new_n590), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n597), .A2(new_n228), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n601), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n596), .A2(new_n599), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n602), .A2(KEYINPUT98), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n605), .B(KEYINPUT98), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n596), .A2(new_n599), .A3(new_n607), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n596), .B2(new_n599), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n555), .A2(new_n557), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n588), .A2(new_n615), .A3(new_n590), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n558), .A2(new_n585), .A3(new_n587), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n558), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n622), .B1(new_n616), .B2(new_n618), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(KEYINPUT99), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n623), .B(new_n629), .C1(KEYINPUT99), .C2(new_n628), .ZN(new_n630));
  INV_X1    g429(.A(new_n622), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n619), .B2(new_n620), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n627), .B1(new_n632), .B2(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n571), .A2(new_n614), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n544), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n514), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n231), .ZN(G1324gat));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  INV_X1    g441(.A(new_n530), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G8gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n641), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n641), .B(new_n649), .C1(new_n644), .C2(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(G8gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(G1325gat));
  NAND2_X1  g451(.A1(new_n350), .A2(new_n355), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT102), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n233), .B1(new_n642), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n536), .A2(new_n538), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n638), .A2(G15gat), .A3(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n655), .A2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n638), .A2(new_n526), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(new_n571), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n635), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n614), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n544), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n514), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n209), .A4(new_n210), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT45), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n520), .B2(new_n526), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n541), .A2(new_n421), .A3(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n519), .A2(new_n673), .B1(new_n542), .B2(new_n539), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n669), .B1(new_n674), .B2(new_n614), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n614), .A2(new_n669), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n526), .B1(new_n488), .B2(new_n490), .ZN(new_n677));
  INV_X1    g476(.A(new_n517), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n514), .B2(new_n515), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n679), .B2(new_n507), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(new_n527), .A3(new_n356), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n539), .A2(new_n542), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n676), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n663), .A2(new_n281), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI22_X1  g485(.A1(new_n686), .A2(new_n514), .B1(new_n223), .B2(new_n222), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n668), .A2(new_n687), .ZN(G1328gat));
  NAND3_X1  g487(.A1(new_n665), .A2(new_n208), .A3(new_n643), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT46), .Z(new_n690));
  OAI21_X1  g489(.A(G36gat), .B1(new_n686), .B2(new_n530), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1329gat));
  OAI211_X1 g491(.A(KEYINPUT47), .B(G43gat), .C1(new_n686), .C2(new_n653), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n656), .A2(G43gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n544), .A2(new_n664), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n544), .A2(KEYINPUT104), .A3(new_n664), .A4(new_n694), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n697), .A2(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n697), .A2(new_n699), .A3(new_n698), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n675), .A2(new_n654), .A3(new_n683), .A4(new_n685), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n704), .A2(G43gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(G1330gat));
  NOR2_X1   g506(.A1(new_n526), .A2(G50gat), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT107), .Z(new_n709));
  NAND3_X1  g508(.A1(new_n544), .A2(new_n664), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT108), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n544), .A2(new_n712), .A3(new_n664), .A4(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n675), .A2(new_n421), .A3(new_n683), .A4(new_n685), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT106), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n714), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n715), .A2(KEYINPUT106), .A3(G50gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n716), .A2(new_n710), .A3(new_n718), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n719), .A2(new_n720), .B1(KEYINPUT48), .B2(new_n721), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n519), .A2(new_n673), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n543), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n609), .A2(new_n613), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n662), .A2(new_n725), .A3(new_n280), .A4(new_n635), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n666), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n530), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  AND2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n731), .B2(new_n732), .ZN(G1333gat));
  NAND3_X1  g534(.A1(new_n728), .A2(G71gat), .A3(new_n654), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n656), .B(KEYINPUT109), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT110), .B1(new_n727), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(G71gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n727), .A2(KEYINPUT110), .A3(new_n737), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n526), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT111), .B(G78gat), .Z(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n571), .A2(new_n280), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n635), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n684), .A2(new_n666), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n670), .A2(new_n672), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n680), .A2(new_n751), .A3(new_n356), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n725), .B(new_n747), .C1(new_n752), .C2(new_n682), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n666), .A2(new_n573), .A3(new_n634), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n750), .A2(new_n573), .B1(new_n756), .B2(new_n757), .ZN(G1336gat));
  NAND4_X1  g557(.A1(new_n675), .A2(new_n643), .A3(new_n683), .A4(new_n749), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n530), .A2(G92gat), .A3(new_n635), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n763), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n724), .A2(new_n725), .A3(new_n747), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n762), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n760), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI211_X1 g568(.A(KEYINPUT113), .B(new_n762), .C1(new_n764), .C2(new_n766), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT52), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(new_n755), .B2(new_n761), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n760), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1337gat));
  NOR3_X1   g573(.A1(new_n656), .A2(G99gat), .A3(new_n635), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n675), .A2(new_n654), .A3(new_n683), .A4(new_n749), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G99gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT114), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n776), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n526), .A2(G106gat), .A3(new_n635), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT53), .B1(new_n755), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n675), .A2(new_n421), .A3(new_n683), .A4(new_n749), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n785), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n764), .A2(new_n766), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n784), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n786), .A2(G106gat), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT53), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n619), .A2(new_n631), .A3(new_n620), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n623), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n626), .B1(new_n632), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n280), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n630), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(KEYINPUT116), .A3(new_n630), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n261), .A2(new_n263), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n257), .B2(new_n203), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n270), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n634), .A2(new_n273), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n614), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n808), .A2(new_n809), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n273), .A2(new_n813), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(new_n798), .B2(new_n800), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n614), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n571), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n636), .A2(new_n280), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n421), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n656), .A2(new_n514), .A3(new_n643), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n309), .B1(new_n827), .B2(new_n280), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n824), .A2(new_n514), .A3(new_n540), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n530), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n281), .A2(new_n312), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT117), .Z(G1340gat));
  INV_X1    g632(.A(new_n827), .ZN(new_n834));
  OAI21_X1  g633(.A(G120gat), .B1(new_n834), .B2(new_n635), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n634), .A2(new_n313), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT118), .Z(new_n837));
  NAND2_X1  g636(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(G1341gat));
  OAI21_X1  g638(.A(G127gat), .B1(new_n834), .B2(new_n662), .ZN(new_n840));
  INV_X1    g639(.A(G127gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n830), .A2(new_n841), .A3(new_n571), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1342gat));
  OAI21_X1  g642(.A(G134gat), .B1(new_n834), .B2(new_n614), .ZN(new_n844));
  INV_X1    g643(.A(G134gat), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n643), .A2(new_n614), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n844), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n851), .B(new_n421), .C1(new_n822), .C2(new_n823), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n356), .A2(new_n514), .A3(new_n643), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n279), .A2(new_n273), .B1(new_n801), .B2(new_n802), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n805), .A2(new_n630), .ZN(new_n855));
  INV_X1    g654(.A(new_n813), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n260), .A2(new_n252), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n277), .A2(new_n274), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n854), .A2(new_n855), .B1(new_n859), .B2(new_n634), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n805), .A2(KEYINPUT116), .A3(new_n630), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT116), .B1(new_n805), .B2(new_n630), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n725), .A2(new_n859), .A3(new_n803), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n860), .A2(new_n725), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n823), .B1(new_n865), .B2(new_n662), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n526), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n853), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G141gat), .B1(new_n868), .B2(new_n281), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n824), .A2(new_n514), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n654), .A2(new_n526), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n643), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n280), .A2(new_n363), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT58), .ZN(G1344gat));
  NAND4_X1  g676(.A1(new_n852), .A2(new_n634), .A3(new_n853), .A4(new_n867), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n361), .A2(KEYINPUT59), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n421), .B1(new_n822), .B2(new_n823), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n421), .A2(new_n851), .ZN(new_n886));
  INV_X1    g685(.A(new_n823), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n814), .B1(new_n804), .B2(new_n806), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n888), .A2(new_n614), .B1(new_n817), .B2(new_n820), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n571), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n893));
  AOI22_X1  g692(.A1(KEYINPUT57), .A2(new_n885), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n853), .A2(new_n634), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n361), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n884), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n892), .A2(new_n893), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n895), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G148gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n883), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n874), .A2(G148gat), .A3(new_n635), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT122), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT121), .B1(new_n902), .B2(KEYINPUT59), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n884), .B(new_n897), .C1(new_n901), .C2(G148gat), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n907), .A2(new_n908), .B1(new_n882), .B2(new_n881), .ZN(new_n909));
  INV_X1    g708(.A(new_n905), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n906), .A2(new_n912), .ZN(G1345gat));
  OAI21_X1  g712(.A(G155gat), .B1(new_n868), .B2(new_n662), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n571), .A2(new_n366), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n874), .B2(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n868), .B2(new_n614), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n846), .A2(new_n367), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n872), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n666), .A2(new_n530), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR4_X1   g720(.A1(new_n737), .A2(new_n824), .A3(new_n421), .A4(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n293), .B1(new_n922), .B2(new_n280), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n824), .A2(new_n666), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n540), .A2(new_n530), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(G169gat), .A3(new_n281), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT123), .ZN(G1348gat));
  OAI21_X1  g728(.A(new_n294), .B1(new_n926), .B2(new_n635), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT124), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n635), .A2(new_n294), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n922), .B2(new_n932), .ZN(G1349gat));
  NAND2_X1  g732(.A1(new_n922), .A2(new_n571), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  INV_X1    g734(.A(new_n926), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n300), .A3(new_n571), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(new_n939), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n301), .A3(new_n725), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n725), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n942), .A2(G190gat), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n942), .B2(G190gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  AND3_X1   g745(.A1(new_n924), .A2(new_n643), .A3(new_n871), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n280), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n654), .A2(new_n921), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n894), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n281), .A2(new_n267), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  INV_X1    g751(.A(new_n950), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n953), .B2(new_n635), .ZN(new_n954));
  INV_X1    g753(.A(G204gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n947), .A2(new_n955), .A3(new_n634), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n954), .B(new_n960), .C1(new_n958), .C2(new_n956), .ZN(G1353gat));
  AOI21_X1  g760(.A(new_n384), .B1(new_n950), .B2(new_n571), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT63), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n384), .A3(new_n571), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n953), .B2(new_n614), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n385), .A3(new_n725), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1355gat));
endmodule


