//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G197gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT86), .ZN(new_n209));
  OR2_X1    g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(KEYINPUT14), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT87), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n215));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n213), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n214), .A2(KEYINPUT15), .A3(new_n216), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT88), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n227), .B2(G1gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n229), .B(new_n230), .Z(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n233), .B1(new_n237), .B2(new_n232), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n223), .B(new_n231), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n239), .B(KEYINPUT13), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT18), .B1(new_n238), .B2(new_n239), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n207), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n238), .A2(new_n239), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n207), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n250), .A2(new_n240), .A3(new_n244), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G85gat), .A2(G92gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT7), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT8), .ZN(new_n256));
  AND2_X1   g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257));
  OAI221_X1 g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .C1(G85gat), .C2(G92gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(G99gat), .A2(G106gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT92), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n260), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT93), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT9), .ZN(new_n266));
  INV_X1    g065(.A(G57gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G64gat), .ZN(new_n268));
  INV_X1    g067(.A(G64gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G57gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n266), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G71gat), .ZN(new_n272));
  INV_X1    g071(.A(G78gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(G71gat), .A2(G78gat), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n271), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n276), .B(KEYINPUT90), .Z(new_n277));
  AOI21_X1  g076(.A(KEYINPUT91), .B1(new_n267), .B2(G64gat), .ZN(new_n278));
  MUX2_X1   g077(.A(KEYINPUT91), .B(new_n278), .S(new_n270), .Z(new_n279));
  AOI21_X1  g078(.A(new_n274), .B1(KEYINPUT9), .B2(new_n275), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT10), .ZN(new_n284));
  INV_X1    g083(.A(new_n282), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n263), .A3(new_n261), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT96), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT96), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n283), .A2(new_n289), .A3(new_n284), .A4(new_n286), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n265), .A2(new_n284), .A3(new_n282), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G230gat), .A2(G233gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT97), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT97), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n292), .B1(new_n288), .B2(new_n290), .ZN(new_n298));
  INV_X1    g097(.A(new_n295), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n295), .B1(new_n283), .B2(new_n286), .ZN(new_n301));
  XOR2_X1   g100(.A(G120gat), .B(G148gat), .Z(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT98), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT99), .ZN(new_n304));
  XOR2_X1   g103(.A(G176gat), .B(G204gat), .Z(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  NOR2_X1   g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n296), .A2(new_n300), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n298), .A2(new_n299), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n309), .B2(new_n301), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n253), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(KEYINPUT41), .ZN(new_n315));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n265), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n235), .B2(new_n236), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(KEYINPUT41), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(new_n223), .B2(new_n265), .ZN(new_n322));
  XNOR2_X1  g121(.A(G190gat), .B(G218gat), .ZN(new_n323));
  OR3_X1    g122(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n320), .B2(new_n322), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n318), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n326), .A2(KEYINPUT94), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(KEYINPUT94), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT95), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n329), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n330), .A2(new_n318), .A3(new_n324), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n335));
  INV_X1    g134(.A(G231gat), .ZN(new_n336));
  INV_X1    g135(.A(G233gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n285), .B2(KEYINPUT21), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT21), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n282), .B(new_n340), .C1(new_n336), .C2(new_n337), .ZN(new_n341));
  XNOR2_X1  g140(.A(G127gat), .B(G155gat), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n342), .B1(new_n339), .B2(new_n341), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n349));
  INV_X1    g148(.A(new_n335), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n231), .B1(new_n285), .B2(KEYINPUT21), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n353), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n345), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G183gat), .B(G211gat), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n354), .B2(new_n356), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n334), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G228gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(new_n337), .ZN(new_n365));
  XNOR2_X1  g164(.A(G197gat), .B(G204gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  INV_X1    g167(.A(G218gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G211gat), .B(G218gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n366), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G155gat), .B(G162gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(G141gat), .A2(G148gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT2), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n377), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n385));
  INV_X1    g184(.A(G141gat), .ZN(new_n386));
  INV_X1    g185(.A(G148gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n388), .A3(new_n378), .ZN(new_n389));
  XOR2_X1   g188(.A(G155gat), .B(G162gat), .Z(new_n390));
  OAI21_X1  g189(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n381), .A2(new_n377), .A3(KEYINPUT72), .A4(new_n383), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n384), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  INV_X1    g195(.A(new_n376), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(new_n397), .B2(KEYINPUT29), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n376), .A2(KEYINPUT81), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI221_X1 g200(.A(new_n365), .B1(new_n376), .B2(new_n395), .C1(new_n401), .C2(new_n393), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT3), .B1(new_n376), .B2(new_n399), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n395), .A2(new_n376), .B1(new_n393), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n365), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(KEYINPUT80), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT80), .B1(new_n404), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G22gat), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n402), .B(new_n411), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT79), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G78gat), .B(G106gat), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT78), .ZN(new_n415));
  XOR2_X1   g214(.A(KEYINPUT31), .B(G50gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n413), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT25), .ZN(new_n419));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT24), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT23), .ZN(new_n426));
  NAND2_X1  g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT23), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(G169gat), .B2(G176gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n419), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT64), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT64), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n419), .C1(new_n424), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n423), .A2(new_n420), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n421), .B2(new_n420), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n429), .A2(KEYINPUT25), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n426), .A2(new_n438), .A3(new_n427), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n426), .B2(new_n427), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n436), .B(new_n437), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(new_n434), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n425), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT26), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT26), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n425), .B1(new_n445), .B2(new_n427), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT27), .B(G183gat), .ZN(new_n447));
  INV_X1    g246(.A(G190gat), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n447), .A2(KEYINPUT28), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT28), .B1(new_n447), .B2(new_n448), .ZN(new_n450));
  OAI221_X1 g249(.A(new_n420), .B1(new_n444), .B2(new_n446), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G134gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G127gat), .ZN(new_n454));
  INV_X1    g253(.A(G127gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G134gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT66), .ZN(new_n458));
  INV_X1    g257(.A(G120gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G113gat), .ZN(new_n460));
  INV_X1    g259(.A(G113gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G120gat), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT1), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n453), .A2(KEYINPUT66), .A3(G127gat), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n458), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n454), .A2(new_n456), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n454), .B2(new_n456), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(new_n463), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n465), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G227gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(new_n337), .ZN(new_n476));
  OR3_X1    g275(.A1(new_n458), .A2(new_n463), .A3(new_n464), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n456), .A3(new_n466), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n471), .B1(new_n480), .B2(new_n463), .ZN(new_n481));
  INV_X1    g280(.A(new_n472), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n442), .A3(new_n451), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n474), .A2(new_n476), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT32), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G15gat), .B(G43gat), .Z(new_n489));
  XNOR2_X1  g288(.A(G71gat), .B(G99gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n491), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n485), .B(KEYINPUT32), .C1(new_n487), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n484), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT34), .B1(new_n497), .B2(new_n476), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n496), .B(new_n499), .C1(new_n475), .C2(new_n337), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n492), .A2(new_n498), .A3(new_n500), .A4(new_n494), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n495), .A2(KEYINPUT69), .A3(new_n501), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n418), .A2(new_n507), .A3(KEYINPUT35), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n452), .A2(new_n399), .ZN(new_n509));
  NAND2_X1  g308(.A1(G226gat), .A2(G233gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n442), .B2(new_n451), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n376), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n515));
  AOI211_X1 g314(.A(new_n515), .B(new_n510), .C1(new_n442), .C2(new_n451), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT29), .B1(new_n442), .B2(new_n451), .ZN(new_n517));
  INV_X1    g316(.A(new_n510), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT70), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n519), .B2(new_n513), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n514), .B1(new_n376), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G8gat), .B(G36gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(G64gat), .B(G92gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT30), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n397), .B(new_n516), .C1(new_n519), .C2(new_n513), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n528), .B2(new_n514), .ZN(new_n529));
  INV_X1    g328(.A(new_n516), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n515), .B1(new_n509), .B2(new_n510), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n376), .B(new_n530), .C1(new_n531), .C2(new_n512), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n513), .B1(new_n518), .B2(new_n517), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n397), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n532), .A2(KEYINPUT30), .A3(new_n534), .A4(new_n525), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n393), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT74), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n473), .A2(new_n540), .A3(new_n393), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(KEYINPUT4), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n473), .A2(new_n393), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  INV_X1    g347(.A(new_n393), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n473), .B1(KEYINPUT3), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(KEYINPUT3), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g350(.A1(G225gat), .A2(G233gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT5), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n546), .A2(new_n548), .A3(new_n551), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT75), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n483), .B2(new_n549), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n473), .A2(KEYINPUT75), .A3(new_n393), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n541), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n553), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT4), .B1(new_n539), .B2(new_n541), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n543), .B(new_n553), .C1(new_n473), .C2(new_n393), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n551), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n564), .A3(KEYINPUT5), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n555), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G1gat), .B(G29gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT0), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G85gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n566), .A2(KEYINPUT6), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n570), .A3(new_n565), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT6), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n555), .B2(new_n565), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n537), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT85), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n537), .A2(new_n577), .A3(KEYINPUT85), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n508), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n502), .A2(new_n505), .ZN(new_n583));
  INV_X1    g382(.A(new_n417), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n413), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n413), .A2(new_n584), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT77), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n574), .B(new_n573), .C1(new_n576), .C2(new_n588), .ZN(new_n589));
  AOI211_X1 g388(.A(KEYINPUT77), .B(new_n570), .C1(new_n555), .C2(new_n565), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n572), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n529), .A2(new_n535), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n592), .B1(new_n529), .B2(new_n535), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n593), .A2(new_n594), .A3(new_n526), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT35), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n524), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n397), .B(new_n530), .C1(new_n531), .C2(new_n512), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n533), .B2(new_n376), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT83), .B(KEYINPUT37), .Z(new_n605));
  NAND3_X1  g404(.A1(new_n532), .A2(new_n534), .A3(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n604), .A2(new_n606), .B1(new_n521), .B2(new_n525), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n572), .B(new_n607), .C1(new_n575), .C2(new_n576), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT84), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n566), .A2(new_n571), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(new_n574), .A3(new_n573), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n612), .A2(KEYINPUT84), .A3(new_n572), .A4(new_n607), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n606), .B(new_n524), .C1(new_n521), .C2(new_n602), .ZN(new_n614));
  INV_X1    g413(.A(new_n599), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n548), .A2(new_n551), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n547), .B1(new_n542), .B2(new_n544), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n553), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n559), .A2(new_n560), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n622), .B2(new_n552), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n621), .B(new_n553), .C1(new_n618), .C2(new_n619), .ZN(new_n625));
  AND4_X1   g424(.A1(KEYINPUT40), .A2(new_n624), .A3(new_n570), .A4(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n571), .B1(new_n620), .B2(new_n623), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT40), .B1(new_n627), .B2(new_n625), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n576), .B1(new_n527), .B2(new_n536), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n418), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n617), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n505), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n507), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n591), .A2(new_n595), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n636), .B2(new_n418), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  AOI211_X1 g437(.A(new_n313), .B(new_n363), .C1(new_n598), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n591), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  INV_X1    g441(.A(new_n537), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G8gat), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT42), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT16), .B(G8gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT100), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  MUX2_X1   g448(.A(KEYINPUT42), .B(new_n646), .S(new_n649), .Z(G1325gat));
  INV_X1    g449(.A(new_n507), .ZN(new_n651));
  AOI21_X1  g450(.A(G15gat), .B1(new_n639), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n635), .A2(G15gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT101), .Z(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n639), .B2(new_n654), .ZN(G1326gat));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n418), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT102), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT43), .B(G22gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  NAND2_X1  g458(.A1(new_n598), .A2(new_n638), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n333), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n313), .A2(new_n362), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n664), .A2(G29gat), .A3(new_n591), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT45), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(KEYINPUT44), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n632), .A2(new_n637), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n598), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n632), .B2(new_n637), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n333), .B(new_n668), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n663), .B(KEYINPUT103), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n591), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n666), .A2(new_n677), .ZN(G1328gat));
  NOR3_X1   g477(.A1(new_n664), .A2(G36gat), .A3(new_n537), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT46), .ZN(new_n680));
  OAI21_X1  g479(.A(G36gat), .B1(new_n676), .B2(new_n537), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1329gat));
  NAND4_X1  g481(.A1(new_n674), .A2(G43gat), .A3(new_n635), .A4(new_n675), .ZN(new_n683));
  INV_X1    g482(.A(G43gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n664), .B2(new_n507), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g486(.A1(new_n418), .A2(G50gat), .ZN(new_n688));
  INV_X1    g487(.A(new_n418), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n664), .A2(new_n689), .ZN(new_n690));
  OAI22_X1  g489(.A1(new_n676), .A2(new_n688), .B1(new_n690), .B2(G50gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g491(.A1(new_n671), .A2(new_n672), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n363), .A2(new_n253), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n311), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT106), .A4(new_n311), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n591), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n267), .ZN(G1332gat));
  AOI211_X1 g500(.A(new_n537), .B(new_n699), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1333gat));
  AND2_X1   g503(.A1(new_n697), .A2(new_n698), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(KEYINPUT107), .A3(new_n651), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n699), .B2(new_n507), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n272), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(G71gat), .A3(new_n635), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n709), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1334gat));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n689), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n273), .ZN(G1335gat));
  NAND3_X1  g515(.A1(new_n247), .A2(new_n361), .A3(new_n252), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n247), .A2(new_n361), .A3(new_n252), .A4(KEYINPUT109), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n333), .B(new_n721), .C1(new_n671), .C2(new_n672), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n312), .A2(G85gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n640), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n311), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT110), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n721), .A2(new_n729), .A3(new_n311), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n674), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G85gat), .B1(new_n732), .B2(new_n591), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT111), .ZN(G1336gat));
  NAND2_X1  g534(.A1(new_n722), .A2(KEYINPUT113), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n723), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n722), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n312), .A2(G92gat), .A3(new_n537), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT112), .Z(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G92gat), .B1(new_n732), .B2(new_n537), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n741), .A2(new_n742), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT52), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(new_n724), .B2(new_n739), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1337gat));
  INV_X1    g549(.A(new_n635), .ZN(new_n751));
  OAI21_X1  g550(.A(G99gat), .B1(new_n732), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n312), .A2(G99gat), .A3(new_n507), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n724), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1338gat));
  OR2_X1    g554(.A1(new_n312), .A2(G106gat), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT115), .B1(new_n756), .B2(new_n689), .ZN(new_n757));
  OR4_X1    g556(.A1(KEYINPUT115), .A2(new_n312), .A3(G106gat), .A4(new_n689), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n724), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n674), .A2(new_n731), .A3(new_n418), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G106gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n759), .A2(KEYINPUT116), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n757), .A2(new_n758), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n737), .A2(new_n738), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT117), .B1(new_n770), .B2(KEYINPUT53), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n772), .B(new_n763), .C1(new_n762), .C2(new_n769), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n764), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT118), .B(new_n764), .C1(new_n771), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1339gat));
  NAND2_X1  g577(.A1(new_n640), .A2(new_n537), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n294), .B2(new_n295), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n298), .A2(KEYINPUT119), .A3(new_n299), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(KEYINPUT54), .A3(new_n300), .A4(new_n296), .ZN(new_n785));
  INV_X1    g584(.A(new_n306), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n309), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n780), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n296), .A2(KEYINPUT54), .A3(new_n300), .ZN(new_n790));
  AND4_X1   g589(.A1(KEYINPUT119), .A2(new_n291), .A3(new_n293), .A4(new_n299), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT119), .B1(new_n298), .B2(new_n299), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n780), .B(new_n788), .C1(new_n790), .C2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n253), .B(new_n308), .C1(new_n789), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n241), .A2(new_n243), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n238), .A2(new_n239), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n206), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n252), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n311), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n333), .B1(new_n796), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n308), .B1(new_n789), .B2(new_n795), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n333), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n361), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n363), .A2(new_n253), .A3(new_n311), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n779), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n587), .ZN(new_n812));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n253), .ZN(new_n813));
  INV_X1    g612(.A(new_n811), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n689), .A2(new_n651), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n253), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n461), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n813), .B1(new_n816), .B2(new_n818), .ZN(G1340gat));
  AOI21_X1  g618(.A(G120gat), .B1(new_n812), .B2(new_n311), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n312), .A2(new_n459), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n816), .B2(new_n821), .ZN(G1341gat));
  NAND3_X1  g621(.A1(new_n812), .A2(new_n455), .A3(new_n362), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n814), .A2(new_n815), .A3(new_n361), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n455), .B2(new_n824), .ZN(G1342gat));
  NAND4_X1  g624(.A1(new_n811), .A2(new_n453), .A3(new_n587), .A4(new_n333), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n814), .A2(new_n815), .A3(new_n334), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n828), .A2(new_n829), .B1(new_n453), .B2(new_n830), .ZN(G1343gat));
  NOR2_X1   g630(.A1(new_n635), .A2(new_n689), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n811), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n386), .B1(new_n833), .B2(new_n817), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n751), .A2(new_n640), .A3(new_n537), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT121), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n689), .B1(new_n808), .B2(new_n810), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n809), .B1(new_n808), .B2(KEYINPUT122), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n841), .B(new_n361), .C1(new_n804), .C2(new_n807), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n689), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n843), .B2(new_n838), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n817), .A2(new_n386), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n834), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n834), .B(KEYINPUT58), .C1(new_n844), .C2(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1344gat));
  OAI21_X1  g650(.A(KEYINPUT59), .B1(new_n833), .B2(new_n312), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n387), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n311), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n808), .A2(new_n810), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n418), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n838), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n312), .A3(new_n836), .ZN(new_n861));
  NAND2_X1  g660(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n862));
  OAI221_X1 g661(.A(new_n853), .B1(new_n844), .B2(new_n855), .C1(new_n861), .C2(new_n862), .ZN(G1345gat));
  OAI21_X1  g662(.A(G155gat), .B1(new_n844), .B2(new_n361), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n361), .A2(G155gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n833), .B2(new_n865), .ZN(G1346gat));
  NAND2_X1  g665(.A1(new_n808), .A2(KEYINPUT122), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n810), .A3(new_n842), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n418), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n333), .A4(new_n839), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n333), .B(new_n839), .C1(new_n843), .C2(new_n838), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT123), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n874), .A3(G162gat), .ZN(new_n875));
  INV_X1    g674(.A(G162gat), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n811), .A2(new_n876), .A3(new_n333), .A4(new_n832), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n640), .A2(new_n537), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT124), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n815), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n204), .A3(new_n817), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n856), .A2(new_n587), .A3(new_n879), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n253), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n204), .ZN(G1348gat));
  INV_X1    g685(.A(G176gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n887), .A3(new_n311), .ZN(new_n888));
  OAI21_X1  g687(.A(G176gat), .B1(new_n882), .B2(new_n312), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1349gat));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n447), .A3(new_n362), .ZN(new_n891));
  OAI21_X1  g690(.A(G183gat), .B1(new_n882), .B2(new_n361), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n882), .B2(new_n334), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT61), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n884), .A2(new_n448), .A3(new_n333), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1351gat));
  AND2_X1   g698(.A1(new_n858), .A2(new_n859), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n880), .A2(new_n635), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G197gat), .B1(new_n902), .B2(new_n817), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n856), .A2(new_n879), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n817), .A2(G197gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n832), .A3(new_n905), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT126), .Z(new_n907));
  NAND2_X1  g706(.A1(new_n903), .A2(new_n907), .ZN(G1352gat));
  NAND3_X1  g707(.A1(new_n900), .A2(new_n311), .A3(new_n901), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G204gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n312), .A2(G204gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n832), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n904), .A2(KEYINPUT127), .A3(new_n832), .A4(new_n911), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n914), .A2(KEYINPUT62), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT62), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(G1353gat));
  AND2_X1   g717(.A1(new_n904), .A2(new_n832), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n368), .A3(new_n362), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n858), .A2(new_n362), .A3(new_n859), .A4(new_n901), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  OAI21_X1  g723(.A(G218gat), .B1(new_n902), .B2(new_n334), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n369), .A3(new_n333), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1355gat));
endmodule


