//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1349, new_n1350, new_n1351,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT65), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT67), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n207), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n202), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(new_n217), .A2(KEYINPUT1), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n219), .A2(new_n223), .A3(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT68), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT70), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT72), .ZN(new_n250));
  AND2_X1   g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(new_n224), .ZN(new_n252));
  AND2_X1   g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(KEYINPUT72), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(G223), .A3(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n259), .B(new_n260), .C1(new_n261), .C2(new_n257), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT71), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n256), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(new_n263), .B2(new_n262), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n253), .A2(new_n254), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(G274), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n265), .B(new_n270), .C1(new_n271), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n277), .B1(G200), .B2(new_n275), .ZN(new_n278));
  INV_X1    g0078(.A(G50), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT75), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT75), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(new_n272), .A3(G13), .A4(G20), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n224), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n281), .B2(new_n283), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n279), .B1(new_n272), .B2(G20), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n279), .A2(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT8), .A2(G58), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT73), .B(G58), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(KEYINPUT8), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G20), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n293), .A2(new_n295), .B1(G150), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n204), .A2(G20), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n298), .A2(KEYINPUT74), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(KEYINPUT74), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n290), .B1(new_n301), .B2(new_n286), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI211_X1 g0104(.A(KEYINPUT9), .B(new_n290), .C1(new_n301), .C2(new_n286), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n278), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n278), .B(new_n308), .C1(new_n304), .C2(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n302), .B1(new_n311), .B2(new_n275), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G179), .B2(new_n275), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n284), .A2(new_n209), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT12), .ZN(new_n316));
  INV_X1    g0116(.A(new_n296), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n279), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n225), .A2(G33), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n319), .A2(new_n261), .B1(new_n225), .B2(G68), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n286), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT11), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n272), .A2(G20), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n287), .A2(G68), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n316), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G226), .A2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G232), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(G1698), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n257), .B1(G33), .B2(G97), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT78), .B1(new_n330), .B2(new_n256), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(G1698), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G226), .B2(G1698), .ZN(new_n334));
  AND2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(KEYINPUT3), .A2(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n332), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n251), .A2(new_n250), .A3(new_n224), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT72), .B1(new_n253), .B2(new_n254), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT78), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n270), .B1(new_n274), .B2(new_n210), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n326), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI211_X1 g0147(.A(KEYINPUT13), .B(new_n345), .C1(new_n331), .C2(new_n343), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n325), .B1(new_n349), .B2(G190), .ZN(new_n350));
  INV_X1    g0150(.A(new_n343), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n342), .B1(new_n338), .B2(new_n341), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n344), .A2(new_n326), .A3(new_n346), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G200), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT8), .B(G58), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n359), .A2(new_n317), .B1(new_n225), .B2(new_n261), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT76), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n295), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n360), .B1(new_n368), .B2(KEYINPUT77), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(KEYINPUT77), .B2(new_n368), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n286), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n261), .B1(new_n272), .B2(G20), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n261), .A2(new_n284), .B1(new_n287), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n251), .A2(new_n224), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n269), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G244), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G232), .A2(G1698), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n258), .A2(G238), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n257), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(G107), .B2(new_n257), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n270), .B(new_n377), .C1(new_n381), .C2(new_n256), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(G179), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n311), .B2(new_n382), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n382), .A2(new_n276), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(G200), .B2(new_n382), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n371), .A2(new_n387), .A3(new_n373), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n358), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n202), .B1(new_n292), .B2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(G159), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n392), .A2(new_n225), .B1(new_n393), .B2(new_n317), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n257), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n209), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n391), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n337), .B2(new_n225), .ZN(new_n400));
  NOR4_X1   g0200(.A1(new_n335), .A2(new_n336), .A3(new_n395), .A4(G20), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(KEYINPUT73), .A2(G58), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT73), .A2(G58), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n227), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(G20), .B1(G159), .B2(new_n296), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n399), .A2(new_n286), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n281), .A2(new_n283), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n293), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n293), .A2(new_n323), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n287), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G274), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n253), .B2(new_n254), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n376), .A2(G232), .B1(new_n269), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n271), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G223), .B2(G1698), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n419), .A2(new_n337), .B1(new_n294), .B2(new_n211), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n341), .ZN(new_n421));
  INV_X1    g0221(.A(G179), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT79), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n417), .A2(new_n421), .A3(KEYINPUT79), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n421), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n425), .A2(new_n426), .B1(new_n311), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n414), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n414), .B2(new_n428), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n417), .A2(new_n421), .A3(new_n276), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n270), .B1(new_n274), .B2(new_n328), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n341), .B2(new_n420), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n435), .B2(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n409), .A2(new_n413), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n409), .A2(new_n436), .A3(KEYINPUT17), .A4(new_n413), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(G169), .C1(new_n347), .C2(new_n348), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n422), .B2(new_n356), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n356), .B2(G169), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n325), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n390), .A2(new_n432), .A3(new_n442), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n314), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT81), .ZN(new_n450));
  INV_X1    g0250(.A(G97), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n294), .A2(G1), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n287), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n410), .A2(new_n451), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n450), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n452), .B(new_n286), .C1(new_n281), .C2(new_n283), .ZN(new_n458));
  OAI211_X1 g0258(.A(KEYINPUT81), .B(new_n455), .C1(new_n458), .C2(new_n451), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  AND2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G97), .A2(G107), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n225), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n317), .A2(new_n261), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT80), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  INV_X1    g0270(.A(new_n468), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT6), .A2(G97), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G107), .ZN(new_n473));
  XNOR2_X1  g0273(.A(G97), .B(G107), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n461), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n470), .B(new_n471), .C1(new_n475), .C2(new_n225), .ZN(new_n476));
  OAI21_X1  g0276(.A(G107), .B1(new_n400), .B2(new_n401), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n469), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n286), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n460), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT85), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G41), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n272), .B(G45), .C1(new_n267), .C2(KEYINPUT5), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT82), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(G41), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT82), .A3(new_n272), .A4(G45), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n375), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n272), .A2(G45), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n486), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n484), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n493), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(G257), .A2(new_n490), .B1(new_n495), .B2(new_n416), .ZN(new_n496));
  OAI211_X1 g0296(.A(G244), .B(new_n258), .C1(new_n335), .C2(new_n336), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G250), .A2(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT4), .A2(G244), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G1698), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n501), .B1(new_n257), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n341), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n482), .B1(new_n496), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n487), .A2(new_n416), .A3(new_n489), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n493), .A2(new_n489), .A3(new_n494), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G257), .A3(new_n266), .ZN(new_n511));
  AND4_X1   g0311(.A1(new_n482), .A2(new_n507), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n311), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G179), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n460), .A2(new_n479), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n481), .A2(new_n513), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n511), .A2(new_n509), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n256), .B1(new_n499), .B2(new_n505), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT84), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n507), .A2(new_n482), .A3(new_n509), .A4(new_n511), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G190), .A3(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n457), .A2(new_n459), .B1(new_n478), .B2(new_n286), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n514), .A2(KEYINPUT83), .A3(G200), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT83), .B1(new_n514), .B2(G200), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n524), .B(new_n525), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n286), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n410), .A2(G116), .A3(new_n531), .A4(new_n453), .ZN(new_n532));
  INV_X1    g0332(.A(G116), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n281), .A2(new_n533), .A3(new_n283), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n285), .A2(new_n224), .B1(G20), .B2(new_n533), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n500), .B(new_n225), .C1(G33), .C2(new_n451), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT20), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n311), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT87), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n510), .A2(G270), .A3(new_n266), .ZN(new_n544));
  OAI211_X1 g0344(.A(G264), .B(G1698), .C1(new_n335), .C2(new_n336), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(new_n258), .C1(new_n335), .C2(new_n336), .ZN(new_n546));
  OR2_X1    g0346(.A1(KEYINPUT3), .A2(G33), .ZN(new_n547));
  NAND2_X1  g0347(.A1(KEYINPUT3), .A2(G33), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(G303), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n341), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n544), .A2(new_n551), .A3(new_n509), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT21), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(KEYINPUT21), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n532), .A2(new_n534), .ZN(new_n555));
  OAI21_X1  g0355(.A(G169), .B1(new_n555), .B2(new_n540), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT87), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n532), .B(new_n534), .C1(new_n539), .C2(new_n538), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n552), .B2(G200), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n276), .B2(new_n552), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n552), .A2(new_n559), .A3(G169), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT21), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n544), .A2(new_n551), .A3(G179), .A4(new_n509), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n562), .A2(new_n563), .B1(new_n565), .B2(new_n559), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n558), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n287), .A2(new_n364), .A3(new_n366), .A4(new_n453), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n364), .A2(new_n366), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n284), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n225), .B1(new_n332), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n463), .A2(new_n211), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n225), .B(G68), .C1(new_n335), .C2(new_n336), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n571), .B1(new_n319), .B2(new_n451), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n286), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n568), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT86), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n284), .A2(new_n569), .B1(new_n577), .B2(new_n286), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n568), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n272), .A2(new_n415), .A3(G45), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n212), .B1(new_n268), .B2(G1), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n266), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G244), .B(G1698), .C1(new_n335), .C2(new_n336), .ZN(new_n589));
  OAI211_X1 g0389(.A(G238), .B(new_n258), .C1(new_n335), .C2(new_n336), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G116), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n588), .B1(new_n592), .B2(new_n341), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n593), .A2(new_n422), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(G169), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G200), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n276), .B(new_n588), .C1(new_n592), .C2(new_n341), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n458), .A2(G87), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n581), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n584), .A2(new_n596), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n225), .B(G87), .C1(new_n335), .C2(new_n336), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT22), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n257), .A2(new_n606), .A3(new_n225), .A4(G87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT24), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT23), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n225), .B2(G107), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n465), .A2(KEYINPUT23), .A3(G20), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(new_n295), .B2(G116), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n608), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n286), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n410), .A2(G107), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n617), .A2(KEYINPUT25), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(KEYINPUT25), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n618), .A2(new_n619), .B1(G107), .B2(new_n458), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n257), .A2(G257), .A3(G1698), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G33), .A2(G294), .ZN(new_n623));
  OAI211_X1 g0423(.A(G250), .B(new_n258), .C1(new_n335), .C2(new_n336), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(G264), .A2(new_n490), .B1(new_n625), .B2(new_n341), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n422), .A3(new_n509), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n509), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n311), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(G200), .B1(new_n626), .B2(new_n509), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n625), .A2(new_n341), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n510), .A2(G264), .A3(new_n266), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n276), .A2(new_n632), .A3(new_n509), .A4(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n616), .B(new_n620), .C1(new_n631), .C2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n603), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n530), .A2(new_n567), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n449), .A2(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n374), .A2(new_n384), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n447), .B1(new_n358), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n442), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n425), .A2(new_n426), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n427), .A2(new_n311), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n413), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n402), .A2(new_n407), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n531), .B1(new_n646), .B2(new_n391), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n647), .B2(new_n408), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT18), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n414), .A2(new_n428), .A3(new_n429), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n310), .B1(new_n641), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n313), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n449), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n580), .A2(new_n583), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n592), .A2(new_n341), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n587), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT88), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n311), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT88), .B1(new_n593), .B2(G169), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n593), .A2(new_n422), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n513), .A2(new_n516), .A3(new_n480), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n600), .A2(new_n602), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n656), .B2(new_n663), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n522), .A2(new_n523), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n515), .B1(new_n671), .B2(new_n311), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n603), .A2(new_n672), .A3(new_n481), .A4(new_n518), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(new_n630), .ZN(new_n675));
  AOI22_X1  g0475(.A1(G270), .A2(new_n490), .B1(new_n495), .B2(new_n416), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n563), .B1(new_n676), .B2(new_n551), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n543), .B1(new_n677), .B2(new_n542), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n554), .A2(new_n556), .A3(KEYINPUT87), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n566), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT89), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT89), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n558), .A2(new_n682), .A3(new_n566), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n675), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n660), .A2(new_n662), .A3(new_n661), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n685), .A2(new_n584), .B1(new_n602), .B2(new_n600), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n519), .A2(new_n529), .A3(new_n635), .A4(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n670), .B(new_n674), .C1(new_n684), .C2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n654), .B1(new_n655), .B2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n681), .A2(new_n683), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n272), .A2(new_n225), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT90), .B(G343), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n559), .ZN(new_n701));
  MUX2_X1   g0501(.A(new_n692), .B(new_n567), .S(new_n701), .Z(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT91), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n691), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n630), .A2(new_n635), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n621), .A2(new_n700), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n630), .B2(new_n699), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n700), .B1(new_n558), .B2(new_n566), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n630), .A2(new_n700), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n220), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n573), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n228), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n687), .B1(new_n692), .B2(new_n630), .ZN(new_n724));
  INV_X1    g0524(.A(new_n664), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n686), .A2(new_n669), .A3(new_n672), .A4(new_n480), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n674), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n699), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT96), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT96), .B(new_n699), .C1(new_n724), .C2(new_n727), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT97), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n730), .A2(KEYINPUT97), .A3(new_n731), .A4(new_n732), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n680), .A2(new_n675), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n687), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n665), .B2(new_n667), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n740), .B(new_n725), .C1(KEYINPUT26), .C2(new_n673), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n699), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n460), .A2(new_n479), .A3(new_n517), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n517), .B1(new_n460), .B2(new_n479), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n524), .A2(new_n525), .ZN(new_n747));
  INV_X1    g0547(.A(new_n528), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n526), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n746), .A2(new_n672), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n567), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n603), .A2(new_n630), .A3(new_n635), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n699), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n508), .A2(new_n512), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT94), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n593), .A2(new_n632), .A3(new_n633), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n564), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT30), .A4(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n757), .A2(KEYINPUT30), .A3(new_n522), .A4(new_n523), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n552), .A2(new_n422), .A3(new_n658), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT93), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n628), .A2(new_n514), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n757), .A2(new_n522), .A3(new_n523), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT30), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT95), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n771), .A3(new_n768), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n761), .A2(new_n766), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n753), .A2(KEYINPUT31), .B1(new_n700), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT31), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n758), .A2(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n775), .B(new_n699), .C1(new_n776), .C2(new_n769), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n743), .A2(KEYINPUT98), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT98), .ZN(new_n781));
  INV_X1    g0581(.A(new_n742), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n735), .B2(new_n736), .ZN(new_n783));
  INV_X1    g0583(.A(new_n779), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n723), .B1(new_n786), .B2(G1), .ZN(G364));
  AND2_X1   g0587(.A1(new_n225), .A2(G13), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n272), .B1(new_n788), .B2(G45), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n717), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n705), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n703), .A2(new_n691), .A3(new_n704), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n703), .A2(new_n704), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n257), .A2(G355), .A3(new_n220), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G116), .B2(new_n220), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n716), .A2(new_n257), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n268), .B2(new_n229), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n243), .A2(G45), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n224), .B1(G20), .B2(new_n311), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n791), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n225), .A2(new_n276), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n597), .A2(G179), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n422), .A2(G200), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G322), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n225), .A2(G190), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n811), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G179), .A2(G200), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n814), .B(new_n821), .C1(G329), .C2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G190), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n276), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G326), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n815), .A2(new_n818), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n337), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n225), .B1(new_n822), .B2(G190), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(G294), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n825), .A2(new_n830), .A3(new_n832), .A4(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n816), .ZN(new_n840));
  INV_X1    g0640(.A(new_n833), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n292), .A2(new_n840), .B1(new_n841), .B2(G77), .ZN(new_n842));
  INV_X1    g0642(.A(new_n831), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n279), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT100), .Z(new_n845));
  OAI221_X1 g0645(.A(new_n257), .B1(new_n819), .B2(new_n465), .C1(new_n211), .C2(new_n812), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT101), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n828), .A2(G68), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n824), .A2(G159), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT32), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n836), .A2(new_n451), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n849), .B2(KEYINPUT32), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n847), .A2(new_n848), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n839), .B1(new_n845), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n809), .B1(new_n854), .B2(new_n806), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n798), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n794), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G396));
  NOR2_X1   g0658(.A1(new_n639), .A2(new_n700), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n374), .A2(new_n700), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n388), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n859), .B1(new_n639), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n699), .B(new_n862), .C1(new_n724), .C2(new_n727), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n730), .A2(new_n732), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n864), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n779), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT102), .Z(new_n867));
  AOI21_X1  g0667(.A(new_n791), .B1(new_n865), .B2(new_n779), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n806), .A2(new_n795), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n791), .B1(G77), .B2(new_n870), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n211), .A2(new_n819), .B1(new_n833), .B2(new_n533), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n812), .A2(new_n465), .B1(new_n823), .B2(new_n834), .ZN(new_n873));
  INV_X1    g0673(.A(G294), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n337), .B1(new_n816), .B2(new_n874), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n872), .A2(new_n873), .A3(new_n875), .A4(new_n851), .ZN(new_n876));
  INV_X1    g0676(.A(new_n828), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n820), .B2(new_n877), .C1(new_n813), .C2(new_n843), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G143), .A2(new_n840), .B1(new_n841), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G150), .ZN(new_n880));
  INV_X1    g0680(.A(G137), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n877), .B2(new_n880), .C1(new_n881), .C2(new_n843), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT34), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n257), .B1(new_n819), .B2(new_n209), .ZN(new_n885));
  INV_X1    g0685(.A(G132), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n812), .A2(new_n279), .B1(new_n823), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n885), .B(new_n887), .C1(new_n292), .C2(new_n837), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n882), .A2(new_n883), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n878), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n871), .B1(new_n891), .B2(new_n806), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n862), .B2(new_n796), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n869), .A2(new_n893), .ZN(G384));
  INV_X1    g0694(.A(new_n475), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(G116), .A4(new_n226), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  NAND3_X1  g0699(.A1(new_n229), .A2(G77), .A3(new_n405), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n201), .A2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n272), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n449), .A2(new_n742), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n653), .B1(new_n737), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n696), .B1(new_n409), .B2(new_n413), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n439), .A2(KEYINPUT107), .A3(new_n440), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n649), .A3(new_n650), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT107), .B1(new_n439), .B2(new_n440), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n414), .A2(new_n428), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n414), .A2(new_n697), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n437), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT106), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n908), .B1(new_n651), .B2(new_n441), .ZN(new_n922));
  XNOR2_X1  g0722(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n923), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n913), .A2(new_n914), .A3(new_n437), .A4(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n922), .A2(KEYINPUT38), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n907), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n447), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT104), .B(new_n325), .C1(new_n445), .C2(new_n446), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n700), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT38), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n914), .B1(new_n432), .B2(new_n442), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n926), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n929), .A2(new_n933), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n859), .B(KEYINPUT103), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n863), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n937), .A2(new_n927), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n325), .A2(new_n700), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n350), .B2(new_n357), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n931), .A2(new_n932), .A3(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n445), .A2(new_n446), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n944), .B1(new_n947), .B2(new_n358), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n942), .A2(new_n943), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n651), .A2(new_n696), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n939), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n906), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n699), .A2(new_n775), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n773), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n773), .A2(KEYINPUT108), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n753), .A2(KEYINPUT31), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n773), .A2(new_n700), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n915), .B(new_n917), .ZN(new_n964));
  INV_X1    g0764(.A(new_n911), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(new_n432), .A3(new_n909), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n908), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n927), .B1(new_n967), .B2(KEYINPUT38), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n861), .A2(new_n639), .ZN(new_n969));
  INV_X1    g0769(.A(new_n859), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n946), .B2(new_n948), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n963), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n957), .A2(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n949), .A2(new_n862), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT40), .B1(new_n937), .B2(new_n927), .ZN(new_n977));
  AOI22_X1  g0777(.A1(KEYINPUT40), .A2(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n655), .B2(new_n974), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n773), .A2(KEYINPUT108), .A3(new_n954), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT108), .B1(new_n773), .B2(new_n954), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n972), .B1(new_n982), .B2(new_n774), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n921), .A2(new_n928), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT40), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n963), .A2(new_n972), .A3(new_n977), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(new_n449), .A3(new_n963), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n979), .A2(new_n988), .A3(G330), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n953), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n272), .B2(new_n788), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n953), .A2(new_n989), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n903), .B1(new_n991), .B2(new_n992), .ZN(G367));
  OAI21_X1  g0793(.A(new_n257), .B1(new_n819), .B2(new_n261), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT113), .Z(new_n995));
  INV_X1    g0795(.A(new_n292), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n996), .A2(new_n812), .B1(new_n881), .B2(new_n823), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n816), .A2(new_n880), .B1(new_n833), .B2(new_n201), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n836), .A2(new_n209), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G143), .A2(new_n831), .B1(new_n828), .B2(G159), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT114), .Z(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n337), .B1(new_n823), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n812), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(G116), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT46), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1007), .A2(new_n1008), .B1(new_n465), .B2(new_n836), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1005), .B(new_n1009), .C1(new_n1008), .C2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n840), .A2(G303), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n819), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G97), .A2(new_n1012), .B1(new_n841), .B2(G283), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n874), .A2(new_n877), .B1(new_n843), .B2(new_n834), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1003), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n806), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n235), .A2(new_n802), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n808), .B1(new_n367), .B2(new_n716), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n717), .B(new_n790), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n797), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n602), .A2(new_n699), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n664), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n667), .B2(new_n1023), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1018), .B(new_n1021), .C1(new_n1022), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT111), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n709), .A2(new_n1027), .A3(new_n711), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n709), .B2(new_n711), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n712), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT112), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1030), .B1(new_n705), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n705), .A2(new_n1031), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n705), .A2(KEYINPUT110), .A3(new_n709), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n750), .B1(new_n525), .B2(new_n699), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n672), .A2(new_n480), .A3(new_n700), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1038), .A2(new_n714), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT44), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n714), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT45), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1035), .B(new_n1044), .Z(new_n1045));
  OAI21_X1  g0845(.A(new_n786), .B1(new_n1034), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n717), .B(KEYINPUT41), .Z(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n790), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n705), .A2(new_n709), .A3(new_n1038), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1038), .A2(new_n712), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT42), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1038), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n519), .B1(new_n1055), .B2(new_n630), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n699), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT109), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT109), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1054), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1025), .B(KEYINPUT43), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1025), .A2(KEYINPUT43), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1051), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n1050), .C1(new_n1065), .C2(new_n1062), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1026), .B1(new_n1049), .B2(new_n1070), .ZN(G387));
  XOR2_X1   g0871(.A(new_n1032), .B(new_n1033), .Z(new_n1072));
  NAND2_X1  g0872(.A1(new_n786), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1034), .A2(new_n780), .A3(new_n785), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n717), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n239), .A2(new_n268), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n359), .A2(G50), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT50), .Z(new_n1078));
  OAI211_X1 g0878(.A(new_n719), .B(new_n268), .C1(new_n209), .C2(new_n261), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n801), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n719), .A2(new_n337), .A3(new_n716), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n465), .B2(new_n716), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT115), .Z(new_n1084));
  OAI21_X1  g0884(.A(new_n807), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n791), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n709), .A2(new_n1022), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n841), .A2(G68), .B1(new_n824), .B2(G150), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n279), .B2(new_n816), .C1(new_n261), .C2(new_n812), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n337), .B(new_n1089), .C1(G97), .C2(new_n1012), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n367), .A2(new_n837), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G159), .A2(new_n831), .B1(new_n828), .B2(new_n293), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G311), .A2(new_n828), .B1(new_n831), .B2(G322), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1094), .A2(KEYINPUT116), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(KEYINPUT116), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G317), .A2(new_n840), .B1(new_n841), .B2(G303), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT48), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n812), .A2(new_n874), .B1(new_n836), .B2(new_n820), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(KEYINPUT49), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n257), .B1(new_n824), .B2(G326), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n533), .C2(new_n819), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT49), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1093), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1086), .B(new_n1087), .C1(new_n806), .C2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n1072), .B2(new_n790), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1075), .A2(new_n1109), .ZN(G393));
  XNOR2_X1  g0910(.A(new_n1035), .B(new_n1044), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n786), .A2(new_n1072), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1034), .B1(new_n785), .B2(new_n780), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1044), .B(new_n710), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n717), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1055), .A2(new_n797), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n248), .A2(new_n802), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n807), .B1(new_n451), .B2(new_n220), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n791), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n831), .A2(G317), .B1(G311), .B2(new_n840), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT52), .Z(new_n1121));
  OAI22_X1  g0921(.A1(new_n812), .A2(new_n820), .B1(new_n823), .B2(new_n817), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n337), .B1(new_n836), .B2(new_n533), .C1(new_n465), .C2(new_n819), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(G294), .C2(new_n841), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1124), .C1(new_n813), .C2(new_n877), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G68), .A2(new_n1006), .B1(new_n824), .B2(G143), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n257), .C1(new_n211), .C2(new_n819), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT118), .Z(new_n1128));
  OAI22_X1  g0928(.A1(new_n843), .A2(new_n880), .B1(new_n393), .B2(new_n816), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n836), .A2(new_n261), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n359), .B2(new_n833), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n201), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n828), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1128), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1125), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1119), .B1(new_n1140), .B2(new_n806), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1114), .A2(new_n790), .B1(new_n1116), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1115), .A2(new_n1142), .ZN(G390));
  OAI211_X1 g0943(.A(new_n699), .B(new_n969), .C1(new_n741), .C2(new_n739), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n970), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n949), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n912), .A2(new_n920), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n934), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n933), .B1(new_n1148), .B2(new_n927), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n778), .A2(G330), .A3(new_n862), .A4(new_n949), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n933), .B1(new_n942), .B2(new_n949), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n937), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n968), .B2(new_n907), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1150), .B(new_n1151), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1144), .A2(new_n970), .B1(new_n946), .B2(new_n948), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n933), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n921), .B2(new_n928), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n674), .A2(new_n725), .A3(new_n726), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n558), .A2(new_n682), .A3(new_n566), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n682), .B1(new_n558), .B2(new_n566), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n630), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND4_X1   g0963(.A1(new_n519), .A2(new_n529), .A3(new_n635), .A4(new_n686), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n700), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n940), .B1(new_n1166), .B2(new_n862), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n949), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1157), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n929), .A2(new_n938), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1159), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n963), .A2(G330), .A3(new_n972), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1155), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n732), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT96), .B1(new_n688), .B2(new_n699), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT97), .B1(new_n1176), .B2(new_n731), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n736), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n905), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n691), .B1(new_n959), .B2(new_n962), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n449), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n654), .A3(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(G330), .B(new_n862), .C1(new_n774), .C2(new_n777), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1168), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1167), .B1(new_n1172), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT119), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1186), .B(G330), .C1(new_n982), .C2(new_n774), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n862), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n963), .B2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1168), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n970), .B(new_n1144), .C1(new_n1183), .C2(new_n1168), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1185), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1173), .B1(new_n1182), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1155), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n863), .A2(new_n941), .B1(new_n946), .B2(new_n948), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1170), .B1(new_n1196), .B2(new_n933), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1172), .B1(new_n1197), .B2(new_n1150), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n904), .B1(new_n735), .B2(new_n736), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1181), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1200), .A2(new_n653), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n971), .B1(new_n1180), .B2(new_n1186), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT119), .B1(new_n974), .B2(new_n691), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n949), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1172), .A2(new_n1184), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1205), .A2(new_n1191), .B1(new_n1167), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1199), .A2(new_n1202), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1194), .A2(new_n1208), .A3(new_n717), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1170), .A2(new_n795), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n791), .B1(new_n293), .B2(new_n870), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1006), .A2(G150), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT53), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1212), .A2(KEYINPUT53), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G159), .C2(new_n837), .ZN(new_n1215));
  INV_X1    g1015(.A(G128), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n843), .C1(new_n881), .C2(new_n877), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n337), .B1(new_n1012), .B2(new_n1136), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT120), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT120), .ZN(new_n1220));
  INV_X1    g1020(.A(G125), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n816), .A2(new_n886), .B1(new_n823), .B2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT54), .B(G143), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1222), .B1(new_n841), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1219), .A2(new_n1220), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n828), .A2(G107), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n257), .B1(new_n1006), .B2(G87), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G116), .A2(new_n840), .B1(new_n841), .B2(G97), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1227), .A2(new_n1134), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n819), .A2(new_n209), .B1(new_n823), .B2(new_n874), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT121), .Z(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n820), .B2(new_n843), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1217), .A2(new_n1226), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1211), .B1(new_n1234), .B2(new_n806), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1210), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1173), .B2(new_n789), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1209), .A2(new_n1238), .ZN(G378));
  XOR2_X1   g1039(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n302), .A2(new_n696), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1242), .A2(KEYINPUT122), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(KEYINPUT122), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n310), .A3(new_n313), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n310), .B2(new_n313), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1241), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n314), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n1240), .A3(new_n1246), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1249), .A2(KEYINPUT123), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n939), .A2(new_n950), .A3(new_n951), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n987), .A2(G330), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n987), .B2(G330), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1254), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n952), .B1(new_n978), .B2(new_n691), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n987), .A2(G330), .A3(new_n1255), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1253), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1249), .A2(new_n795), .A3(new_n1252), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n791), .B1(new_n1136), .B2(new_n870), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n257), .A2(G41), .ZN(new_n1265));
  AOI211_X1 g1065(.A(G50), .B(new_n1265), .C1(new_n294), .C2(new_n267), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n261), .B2(new_n812), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n816), .A2(new_n465), .B1(new_n823), .B2(new_n820), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n996), .A2(new_n819), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n999), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G97), .A2(new_n828), .B1(new_n831), .B2(G116), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(new_n569), .C2(new_n833), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT58), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1266), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n833), .A2(new_n881), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1216), .A2(new_n816), .B1(new_n812), .B2(new_n1223), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1275), .B(new_n1276), .C1(G150), .C2(new_n837), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1277), .B1(new_n1221), .B2(new_n843), .C1(new_n886), .C2(new_n877), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT59), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n294), .B(new_n267), .C1(new_n819), .C2(new_n393), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G124), .B2(new_n824), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1278), .A2(KEYINPUT59), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n1274), .B1(new_n1273), .B2(new_n1272), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1264), .B1(new_n1284), .B2(new_n806), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1262), .A2(new_n790), .B1(new_n1263), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1182), .A2(KEYINPUT124), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n906), .A2(new_n1288), .A3(new_n1181), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1208), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT57), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n717), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT57), .B1(new_n1290), .B2(new_n1262), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1286), .B1(new_n1294), .B2(new_n1295), .ZN(G375));
  NOR2_X1   g1096(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1204), .A2(new_n862), .A3(new_n1187), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1191), .B1(new_n1299), .B2(new_n1168), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n906), .B(new_n1181), .C1(new_n1185), .C2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1301), .A3(new_n1048), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1168), .A2(new_n795), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n791), .B1(G68), .B2(new_n870), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(G116), .A2(new_n828), .B1(new_n831), .B2(G294), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n257), .B1(new_n1012), .B2(G77), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n816), .A2(new_n820), .B1(new_n833), .B2(new_n465), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n812), .A2(new_n451), .B1(new_n823), .B2(new_n813), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1305), .A2(new_n1091), .A3(new_n1306), .A4(new_n1309), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n337), .B(new_n1269), .C1(G50), .C2(new_n837), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n843), .B2(new_n886), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n828), .A2(new_n1224), .ZN(new_n1314));
  OAI22_X1  g1114(.A1(new_n812), .A2(new_n393), .B1(new_n833), .B2(new_n880), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n816), .A2(new_n881), .B1(new_n823), .B2(new_n1216), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1311), .A2(new_n1313), .A3(new_n1314), .A4(new_n1317), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n843), .A2(new_n1312), .A3(new_n886), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1310), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1304), .B1(new_n1320), .B2(new_n806), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1207), .A2(new_n790), .B1(new_n1303), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1302), .A2(new_n1322), .ZN(G381));
  INV_X1    g1123(.A(G384), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n718), .B1(new_n1301), .B2(new_n1173), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1237), .B1(new_n1325), .B2(new_n1208), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1324), .A2(new_n1326), .A3(new_n1322), .A4(new_n1302), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1075), .A2(new_n857), .A3(new_n1109), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1327), .A2(G390), .A3(new_n1328), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1072), .A2(new_n1111), .B1(new_n780), .B2(new_n785), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n789), .B1(new_n1330), .B2(new_n1047), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(new_n1069), .A3(new_n1067), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1259), .A2(new_n1253), .A3(new_n1260), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1253), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n790), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1263), .A2(new_n1285), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1182), .A2(new_n1173), .A3(new_n1193), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1262), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1291), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n718), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1337), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1329), .A2(new_n1026), .A3(new_n1332), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1347));
  OR2_X1    g1147(.A1(new_n1346), .A2(new_n1347), .ZN(G407));
  INV_X1    g1148(.A(G213), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n698), .A2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1343), .A2(new_n1326), .A3(new_n1350), .ZN(new_n1351));
  OAI211_X1 g1151(.A(G213), .B(new_n1351), .C1(new_n1346), .C2(new_n1347), .ZN(G409));
  INV_X1    g1152(.A(new_n1350), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT60), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1355), .A2(new_n1297), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1182), .A2(KEYINPUT60), .A3(new_n1193), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n717), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1322), .B1(new_n1356), .B2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1324), .ZN(new_n1360));
  OAI211_X1 g1160(.A(G384), .B(new_n1322), .C1(new_n1356), .C2(new_n1358), .ZN(new_n1361));
  AND2_X1   g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  AOI211_X1 g1162(.A(new_n1337), .B(new_n1326), .C1(new_n1341), .C2(new_n1342), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1290), .A2(new_n1048), .A3(new_n1262), .ZN(new_n1364));
  AOI21_X1  g1164(.A(G378), .B1(new_n1364), .B2(new_n1286), .ZN(new_n1365));
  OAI211_X1 g1165(.A(new_n1353), .B(new_n1362), .C1(new_n1363), .C2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(KEYINPUT62), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT61), .ZN(new_n1368));
  OAI211_X1 g1168(.A(G378), .B(new_n1286), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1365), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT62), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1371), .A2(new_n1372), .A3(new_n1353), .A4(new_n1362), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1350), .A2(G2897), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1360), .A2(new_n1361), .A3(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1374), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  AOI21_X1  g1178(.A(new_n1365), .B1(new_n1343), .B2(G378), .ZN(new_n1379));
  OAI211_X1 g1179(.A(new_n1375), .B(new_n1378), .C1(new_n1379), .C2(new_n1350), .ZN(new_n1380));
  NAND4_X1  g1180(.A1(new_n1367), .A2(new_n1368), .A3(new_n1373), .A4(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1328), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n857), .B1(new_n1075), .B2(new_n1109), .ZN(new_n1383));
  NOR2_X1   g1183(.A1(new_n1382), .A2(new_n1383), .ZN(new_n1384));
  AND2_X1   g1184(.A1(G387), .A2(G390), .ZN(new_n1385));
  NOR2_X1   g1185(.A1(G387), .A2(G390), .ZN(new_n1386));
  OAI211_X1 g1186(.A(KEYINPUT127), .B(new_n1384), .C1(new_n1385), .C2(new_n1386), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT127), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1388), .B1(new_n1382), .B2(new_n1383), .ZN(new_n1389));
  INV_X1    g1189(.A(new_n1383), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1390), .A2(KEYINPUT127), .A3(new_n1328), .ZN(new_n1391));
  NAND4_X1  g1191(.A1(new_n1332), .A2(new_n1026), .A3(new_n1115), .A4(new_n1142), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(G387), .A2(G390), .ZN(new_n1393));
  NAND4_X1  g1193(.A1(new_n1389), .A2(new_n1391), .A3(new_n1392), .A4(new_n1393), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1387), .A2(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1381), .A2(new_n1395), .ZN(new_n1396));
  AND2_X1   g1196(.A1(new_n1378), .A2(new_n1375), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1371), .A2(new_n1353), .ZN(new_n1398));
  AOI21_X1  g1198(.A(KEYINPUT61), .B1(new_n1397), .B2(new_n1398), .ZN(new_n1399));
  AND2_X1   g1199(.A1(new_n1387), .A2(new_n1394), .ZN(new_n1400));
  INV_X1    g1200(.A(KEYINPUT63), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1366), .A2(new_n1401), .ZN(new_n1402));
  NAND4_X1  g1202(.A1(new_n1371), .A2(KEYINPUT63), .A3(new_n1353), .A4(new_n1362), .ZN(new_n1403));
  NAND4_X1  g1203(.A1(new_n1399), .A2(new_n1400), .A3(new_n1402), .A4(new_n1403), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1396), .A2(new_n1404), .ZN(G405));
  NAND2_X1  g1205(.A1(G375), .A2(new_n1326), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1406), .A2(new_n1369), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1407), .A2(new_n1362), .ZN(new_n1408));
  NAND3_X1  g1208(.A1(new_n1406), .A2(new_n1369), .A3(new_n1376), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(new_n1408), .A2(new_n1409), .ZN(new_n1410));
  XNOR2_X1  g1210(.A(new_n1410), .B(new_n1395), .ZN(G402));
endmodule


