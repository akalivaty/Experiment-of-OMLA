//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT66), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  XOR2_X1   g041(.A(KEYINPUT3), .B(G2104), .Z(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  INV_X1    g047(.A(G136), .ZN(new_n473));
  AND2_X1   g048(.A1(G112), .A2(G2105), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n474), .B1(G100), .B2(new_n460), .ZN(new_n475));
  OAI22_X1  g050(.A1(new_n461), .A2(new_n473), .B1(new_n475), .B2(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n459), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n477), .B(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n476), .B1(new_n479), .B2(G124), .ZN(G162));
  NAND2_X1  g055(.A1(KEYINPUT4), .A2(G138), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n467), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(G102), .A2(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n460), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(G114), .A2(G2104), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n467), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n461), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n484), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  XNOR2_X1  g068(.A(KEYINPUT5), .B(G543), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n494), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n494), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(G166));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n494), .B(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n496), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(new_n494), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G89), .ZN(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n506), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT70), .B1(new_n499), .B2(new_n500), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n508), .A2(new_n519), .A3(new_n509), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G168));
  XOR2_X1   g098(.A(KEYINPUT5), .B(G543), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n504), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G64), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n496), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n521), .A2(G52), .B1(new_n512), .B2(G90), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(G68), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n525), .A2(new_n526), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n521), .A2(G43), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n512), .A2(G81), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT73), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT73), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n541), .B(new_n548), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n518), .A2(new_n520), .ZN(new_n560));
  AND4_X1   g135(.A1(new_n559), .A2(new_n560), .A3(G53), .A4(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n559), .B1(new_n521), .B2(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT70), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n519), .B1(new_n508), .B2(new_n509), .ZN(new_n565));
  OAI21_X1  g140(.A(G543), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n521), .A2(new_n559), .A3(G53), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(KEYINPUT75), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n524), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n512), .B2(G91), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n563), .A2(new_n570), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  XNOR2_X1  g151(.A(G166), .B(KEYINPUT76), .ZN(G303));
  OAI21_X1  g152(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n511), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n521), .A2(G49), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n580), .A2(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n494), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n496), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(G86), .B2(new_n512), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n538), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n496), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n521), .A2(G47), .B1(new_n512), .B2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n599), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT81), .B1(new_n511), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n510), .A2(new_n494), .A3(new_n607), .A4(G92), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n606), .B2(new_n608), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT82), .B(G66), .Z(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(new_n494), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n566), .A2(new_n612), .B1(new_n614), .B2(new_n496), .ZN(new_n615));
  NOR3_X1   g190(.A1(new_n610), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g194(.A(new_n618), .B1(G171), .B2(G868), .ZN(G321));
  MUX2_X1   g195(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g196(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n551), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n462), .A2(G135), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  MUX2_X1   g206(.A(G99), .B(G111), .S(G2105), .Z(new_n632));
  AOI22_X1  g207(.A1(new_n479), .A2(G123), .B1(G2104), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT84), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n462), .A2(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(new_n636), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n637), .A2(new_n641), .A3(new_n642), .ZN(G156));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT85), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT15), .B(G2435), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2438), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2427), .Z(new_n653));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n653), .B2(G2430), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(G2430), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g230(.A(G14), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n650), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT17), .Z(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n662), .ZN(new_n665));
  INV_X1    g240(.A(new_n658), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n661), .C1(new_n666), .C2(new_n662), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n660), .A3(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n636), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2100), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n675), .A2(new_n680), .A3(new_n678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n683));
  AOI211_X1 g258(.A(new_n679), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NOR2_X1   g267(.A1(G171), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G5), .B2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G1961), .ZN(new_n696));
  INV_X1    g271(.A(G140), .ZN(new_n697));
  AND2_X1   g272(.A1(G116), .A2(G2105), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G104), .B2(new_n460), .ZN(new_n699));
  OAI22_X1  g274(.A1(new_n461), .A2(new_n697), .B1(new_n699), .B2(new_n463), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n479), .B2(G128), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT92), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(G26), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2067), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n696), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n464), .A2(G103), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G139), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n712), .B(new_n713), .C1(new_n461), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT94), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n460), .B2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G33), .B(new_n718), .S(G29), .Z(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G2072), .Z(new_n720));
  INV_X1    g295(.A(G1348), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n616), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G4), .B2(G16), .ZN(new_n723));
  NOR2_X1   g298(.A1(G29), .A2(G35), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G162), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT29), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n720), .B1(new_n721), .B2(new_n723), .C1(G2090), .C2(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n695), .A2(G1961), .ZN(new_n728));
  NOR2_X1   g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(KEYINPUT24), .A2(G34), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G160), .B2(G29), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G2084), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G2084), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT31), .B(G11), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT30), .B(G28), .Z(new_n737));
  OAI211_X1 g312(.A(new_n735), .B(new_n736), .C1(G29), .C2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n734), .B(new_n738), .C1(G29), .C2(new_n635), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n692), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n692), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1966), .ZN(new_n742));
  NOR2_X1   g317(.A1(G27), .A2(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G164), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2078), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n702), .A2(G32), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n464), .A2(G105), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n749), .B(new_n750), .C1(new_n479), .C2(G129), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n462), .A2(G141), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT95), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(new_n702), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n723), .A2(new_n721), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n739), .A2(new_n746), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n709), .A2(new_n727), .A3(new_n728), .A4(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n692), .A2(KEYINPUT88), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n692), .A2(KEYINPUT88), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  MUX2_X1   g339(.A(G19), .B(new_n550), .S(new_n764), .Z(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  NAND3_X1  g341(.A1(new_n762), .A2(G20), .A3(new_n763), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT96), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G16), .B2(G299), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n726), .A2(G2090), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n761), .B(new_n766), .C1(KEYINPUT97), .C2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G25), .A2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G131), .ZN(new_n779));
  AND2_X1   g354(.A1(G107), .A2(G2105), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G95), .B2(new_n460), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n461), .A2(new_n779), .B1(new_n781), .B2(new_n463), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n479), .B2(G119), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT35), .B(G1991), .Z(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n603), .A2(new_n764), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G24), .B2(new_n764), .ZN(new_n788));
  INV_X1    g363(.A(G1986), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G23), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G288), .B2(new_n692), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT33), .B(G1976), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G6), .B(G305), .S(G16), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n764), .A2(G22), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n764), .ZN(new_n800));
  INV_X1    g375(.A(G1971), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n795), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI221_X1 g379(.A(new_n790), .B1(new_n789), .B2(new_n788), .C1(KEYINPUT34), .C2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n803), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(KEYINPUT91), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n810), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n777), .B1(new_n811), .B2(new_n812), .ZN(G311));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(new_n776), .ZN(G150));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n566), .A2(new_n816), .B1(new_n817), .B2(new_n511), .ZN(new_n818));
  INV_X1    g393(.A(G67), .ZN(new_n819));
  INV_X1    g394(.A(G80), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n538), .A2(new_n819), .B1(new_n820), .B2(new_n517), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n496), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI221_X1 g398(.A(KEYINPUT98), .B1(new_n820), .B2(new_n517), .C1(new_n538), .C2(new_n819), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(G860), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n616), .A2(G559), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT38), .Z(new_n830));
  AND2_X1   g405(.A1(new_n823), .A2(new_n824), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n547), .B(new_n549), .C1(new_n831), .C2(new_n818), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n825), .A2(new_n546), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n830), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(new_n826), .C1(new_n836), .C2(new_n835), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n828), .B1(new_n839), .B2(new_n840), .ZN(G145));
  XNOR2_X1  g416(.A(new_n718), .B(new_n754), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n701), .B(new_n492), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n639), .B(new_n783), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n479), .A2(G130), .ZN(new_n846));
  MUX2_X1   g421(.A(G106), .B(G118), .S(G2105), .Z(new_n847));
  AOI22_X1  g422(.A1(new_n462), .A2(G142), .B1(G2104), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n845), .B(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n844), .A2(new_n850), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(KEYINPUT100), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(KEYINPUT100), .B2(new_n852), .ZN(new_n854));
  XNOR2_X1  g429(.A(G160), .B(G162), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n635), .B(new_n855), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  INV_X1    g433(.A(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n851), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g437(.A1(new_n825), .A2(new_n626), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n834), .B(new_n625), .Z(new_n864));
  OR2_X1    g439(.A1(G299), .A2(new_n616), .ZN(new_n865));
  AND3_X1   g440(.A1(G299), .A2(KEYINPUT101), .A3(new_n616), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT101), .B1(G299), .B2(new_n616), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(G299), .A2(new_n616), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(G299), .A2(KEYINPUT101), .A3(new_n616), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n865), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n873), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(new_n878), .B2(new_n865), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n869), .B2(new_n874), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT104), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n872), .A2(KEYINPUT102), .A3(new_n873), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n881), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n879), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(new_n864), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n877), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n580), .A2(new_n581), .ZN(new_n892));
  INV_X1    g467(.A(new_n602), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n600), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n603), .A2(new_n892), .ZN(new_n896));
  XNOR2_X1  g471(.A(G305), .B(G166), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n601), .A2(G288), .A3(new_n602), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n891), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n863), .B1(new_n909), .B2(G868), .ZN(G295));
  AOI21_X1  g485(.A(new_n863), .B1(new_n909), .B2(G868), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  NAND2_X1  g487(.A1(G301), .A2(G286), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n531), .A2(new_n534), .A3(G168), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n833), .A3(new_n832), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n834), .A2(new_n913), .A3(new_n914), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n875), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n917), .A2(new_n916), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n919), .B(new_n902), .C1(new_n889), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n858), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n916), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT41), .B1(new_n886), .B2(new_n865), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n880), .B1(new_n872), .B2(new_n873), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n918), .B1(new_n926), .B2(KEYINPUT107), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n902), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n879), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n887), .B1(new_n886), .B2(new_n881), .ZN(new_n933));
  AOI211_X1 g508(.A(KEYINPUT104), .B(new_n880), .C1(new_n884), .C2(new_n885), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n918), .B1(new_n935), .B2(new_n923), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n936), .B2(new_n902), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n919), .B1(new_n889), .B2(new_n920), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n903), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n912), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n937), .B2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n925), .B1(new_n875), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n945), .B2(new_n920), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n929), .A3(new_n919), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n903), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n937), .A2(new_n948), .A3(new_n940), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n937), .A2(new_n948), .A3(KEYINPUT108), .A4(new_n940), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI211_X1 g528(.A(KEYINPUT109), .B(new_n942), .C1(new_n953), .C2(new_n912), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  INV_X1    g530(.A(new_n943), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n922), .A2(new_n930), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT108), .B1(new_n957), .B2(new_n940), .ZN(new_n958));
  INV_X1    g533(.A(new_n952), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n912), .B(new_n956), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n942), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n954), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n492), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT110), .B(G40), .Z(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n465), .A2(new_n470), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n701), .B(G2067), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n755), .B2(new_n973), .ZN(new_n974));
  OR3_X1    g549(.A1(new_n972), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT46), .B1(new_n972), .B2(G1996), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n754), .A2(G1996), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n973), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n783), .B(new_n785), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n971), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n971), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  INV_X1    g564(.A(G2067), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n701), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n783), .A2(new_n785), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n982), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n978), .B(new_n989), .C1(new_n971), .C2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(G305), .A2(G1981), .ZN(new_n995));
  INV_X1    g570(.A(new_n587), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT112), .B(G86), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n511), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(G1981), .B1(new_n998), .B2(new_n584), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n1000), .A2(KEYINPUT49), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n492), .A2(new_n964), .ZN(new_n1002));
  INV_X1    g577(.A(new_n970), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n995), .A2(KEYINPUT49), .A3(new_n999), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1001), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n892), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(new_n995), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1007), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n492), .A2(KEYINPUT50), .A3(new_n964), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT50), .B1(new_n492), .B2(new_n964), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1003), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1016), .A2(G2090), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n970), .B1(new_n965), .B2(new_n966), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n801), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1006), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT55), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n892), .A2(new_n1026), .A3(G1976), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT111), .B1(G288), .B2(new_n1010), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1007), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n892), .A2(G1976), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n1029), .A2(KEYINPUT52), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1009), .A3(new_n1032), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1012), .A2(new_n1013), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1016), .A2(G2084), .ZN(new_n1036));
  INV_X1    g611(.A(G1966), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1020), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1006), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1039), .A2(G168), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(KEYINPUT63), .A3(new_n1025), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1033), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT113), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1025), .A3(new_n1040), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT63), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT114), .B(new_n1035), .C1(new_n1047), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1046), .A2(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1053), .B2(new_n1034), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(G301), .B(KEYINPUT54), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1016), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT116), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1016), .A2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT125), .B(G1961), .Z(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1020), .B2(G2078), .ZN(new_n1065));
  XOR2_X1   g640(.A(new_n465), .B(KEYINPUT126), .Z(new_n1066));
  NAND2_X1  g641(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1067));
  AOI211_X1 g642(.A(G2078), .B(new_n1067), .C1(new_n469), .C2(G2105), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(new_n967), .A3(new_n1019), .A4(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1057), .A2(new_n1063), .A3(new_n1065), .A4(new_n1069), .ZN(new_n1070));
  OR3_X1    g645(.A1(new_n1020), .A2(new_n1064), .A3(G2078), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1063), .A2(new_n1065), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(new_n1057), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT123), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1036), .A2(new_n1077), .A3(new_n1038), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1006), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT124), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G168), .A2(new_n1006), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1079), .A2(KEYINPUT124), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT51), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1039), .A2(KEYINPUT51), .A3(new_n1081), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1081), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1074), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1059), .A2(new_n721), .A3(new_n1061), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1005), .A2(new_n990), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n617), .A2(KEYINPUT60), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  INV_X1    g674(.A(G1956), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1098), .A2(new_n1099), .B1(new_n1016), .B2(new_n1100), .ZN(new_n1101));
  AND2_X1   g676(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1102));
  INV_X1    g677(.A(new_n574), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT57), .B(new_n1103), .C1(new_n568), .C2(new_n569), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT61), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1016), .A2(new_n1100), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1107), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1097), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1105), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1113), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1096), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1093), .A2(new_n617), .A3(new_n1094), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n617), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT60), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n967), .A2(new_n979), .A3(new_n1003), .A4(new_n1019), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1018), .A2(KEYINPUT117), .A3(new_n979), .A4(new_n1019), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1004), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n550), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT118), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1122), .A2(new_n1123), .B1(new_n1004), .B2(new_n1125), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1130), .B(KEYINPUT59), .C1(new_n1131), .C2(new_n550), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1128), .A3(new_n551), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1127), .A2(KEYINPUT119), .A3(new_n1128), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1116), .B(new_n1119), .C1(new_n1133), .C2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1118), .B1(new_n1112), .B2(new_n1111), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1109), .B(KEYINPUT115), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1092), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1146), .ZN(new_n1148));
  AOI211_X1 g723(.A(KEYINPUT122), .B(new_n1148), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1091), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1079), .A2(KEYINPUT124), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1081), .B1(new_n1079), .B2(KEYINPUT124), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1090), .B1(new_n1154), .B2(new_n1086), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT62), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(new_n1090), .C1(new_n1154), .C2(new_n1086), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1156), .A2(G171), .A3(new_n1072), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1150), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1043), .A2(new_n1025), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1055), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n982), .B(new_n983), .C1(G290), .C2(G1986), .ZN(new_n1164));
  INV_X1    g739(.A(new_n985), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n972), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n994), .B1(new_n1163), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g742(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n672), .A2(G319), .ZN(new_n1171));
  NOR3_X1   g745(.A1(new_n1171), .A2(G401), .A3(G229), .ZN(new_n1172));
  NAND4_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n861), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n861), .A2(new_n1172), .ZN(new_n1174));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(new_n953), .B2(new_n1174), .ZN(new_n1175));
  AND2_X1   g749(.A1(new_n1173), .A2(new_n1175), .ZN(G308));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(G225));
endmodule


