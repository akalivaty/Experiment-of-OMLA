//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT13), .Z(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G1gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G1gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n215), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n217), .A2(new_n211), .A3(G8gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n221));
  NOR3_X1   g020(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT91), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G29gat), .ZN(new_n228));
  INV_X1    g027(.A(G36gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n227), .A2(KEYINPUT92), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n227), .A2(KEYINPUT92), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n221), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n223), .ZN(new_n233));
  OAI22_X1  g032(.A1(new_n220), .A2(KEYINPUT15), .B1(new_n233), .B2(new_n222), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n228), .A2(new_n229), .ZN(new_n235));
  OR3_X1    g034(.A1(new_n234), .A2(new_n221), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n219), .B1(new_n232), .B2(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n208), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n219), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT17), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n232), .A2(new_n244), .A3(new_n236), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n241), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT18), .A3(new_n207), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n240), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n232), .A2(new_n244), .A3(new_n236), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n244), .B1(new_n232), .B2(new_n236), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n219), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n207), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n239), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT18), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n206), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT18), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n239), .A2(new_n257), .A3(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n247), .A2(new_n237), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n258), .A2(new_n252), .B1(new_n259), .B2(new_n208), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n247), .A2(new_n207), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n257), .B1(new_n246), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n206), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n264), .A3(KEYINPUT93), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G211gat), .A2(G218gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274));
  AND2_X1   g073(.A1(G197gat), .A2(G204gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G211gat), .B(G218gat), .Z(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G197gat), .B(G204gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n280), .A3(new_n273), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(KEYINPUT24), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT67), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n285), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(G183gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n284), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n289), .A2(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT69), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT23), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(KEYINPUT25), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n313), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n309), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n304), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n318), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n292), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n289), .A2(new_n296), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n317), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n312), .A2(new_n314), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT65), .B(G176gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n313), .A2(G169gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n324), .A3(new_n327), .A4(new_n308), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT68), .B(G190gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT27), .B(G183gat), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n335), .A2(KEYINPUT28), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n308), .B1(new_n311), .B2(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n286), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n335), .B2(KEYINPUT28), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n331), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n331), .B2(new_n342), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n283), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n342), .A3(new_n343), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n316), .A2(new_n330), .B1(new_n336), .B2(new_n341), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n348), .B(new_n282), .C1(new_n349), .C2(new_n345), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(KEYINPUT75), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n344), .A2(new_n346), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n282), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n351), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(KEYINPUT30), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n355), .A2(new_n363), .A3(new_n358), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  INV_X1    g167(.A(G155gat), .ZN(new_n369));
  INV_X1    g168(.A(G162gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G141gat), .B(G148gat), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n368), .B(new_n371), .C1(new_n372), .C2(KEYINPUT2), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374));
  INV_X1    g173(.A(G148gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(G141gat), .ZN(new_n376));
  INV_X1    g175(.A(G141gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(G141gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n369), .A3(new_n370), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n368), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n373), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT71), .ZN(new_n386));
  INV_X1    g185(.A(G134gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(G127gat), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n387), .A2(G127gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n390), .B2(new_n393), .ZN(new_n395));
  INV_X1    g194(.A(G120gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G113gat), .ZN(new_n397));
  INV_X1    g196(.A(G113gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G120gat), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT1), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n394), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G127gat), .B(G134gat), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n385), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n406));
  INV_X1    g205(.A(G127gat), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT72), .B1(new_n408), .B2(new_n392), .ZN(new_n409));
  INV_X1    g208(.A(new_n400), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n403), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n375), .A2(G141gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n377), .A2(G148gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n381), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n371), .A2(new_n368), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n416), .A2(new_n417), .B1(new_n380), .B2(new_n383), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n412), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n367), .B1(new_n404), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n366), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n412), .A2(new_n413), .A3(new_n418), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n418), .B1(new_n412), .B2(new_n413), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT78), .B(KEYINPUT5), .C1(new_n425), .C2(new_n367), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT73), .B1(new_n401), .B2(new_n403), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT73), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n428), .A3(new_n413), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT77), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n373), .A2(new_n384), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(new_n373), .B2(new_n384), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(KEYINPUT4), .A3(new_n429), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n367), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n373), .A2(new_n384), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n373), .B2(new_n384), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n412), .A2(new_n413), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n437), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n434), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n422), .A2(new_n426), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n439), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n390), .A2(new_n393), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n400), .B1(new_n449), .B2(KEYINPUT72), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n403), .B1(new_n450), .B2(new_n411), .ZN(new_n451));
  OAI22_X1  g250(.A1(new_n448), .A2(new_n451), .B1(new_n419), .B2(new_n435), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(new_n435), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n437), .A2(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G1gat), .B(G29gat), .Z(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G57gat), .B(G85gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT80), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n462), .B2(new_n464), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n446), .B2(new_n456), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n464), .B(new_n461), .C1(new_n446), .C2(new_n456), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n365), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G15gat), .B(G43gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(G71gat), .B(G99gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G227gat), .A2(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n349), .A2(new_n427), .A3(new_n429), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n427), .A2(new_n429), .B1(new_n331), .B2(new_n342), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT69), .B1(new_n302), .B2(new_n303), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n329), .B1(G169gat), .B2(G176gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n324), .A2(new_n307), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n484), .A2(new_n304), .B1(new_n329), .B2(new_n328), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n336), .A2(new_n341), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT73), .B(new_n403), .C1(new_n450), .C2(new_n411), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n428), .B1(new_n412), .B2(new_n413), .ZN(new_n488));
  OAI22_X1  g287(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n349), .A2(new_n427), .A3(new_n429), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n474), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT34), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n489), .A2(new_n490), .A3(new_n493), .A4(new_n474), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n490), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT33), .B1(new_n497), .B2(new_n475), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n492), .B(new_n494), .C1(new_n498), .C2(new_n473), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n496), .B2(new_n499), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G78gat), .B(G106gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G50gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(KEYINPUT81), .Z(new_n507));
  INV_X1    g306(.A(G22gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n385), .A2(KEYINPUT77), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n418), .A2(new_n430), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n276), .A2(new_n277), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n279), .B1(new_n273), .B2(new_n280), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n510), .A2(new_n511), .B1(new_n515), .B2(new_n438), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n282), .B1(new_n439), .B2(new_n512), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT29), .B1(new_n278), .B2(new_n281), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n385), .B1(new_n519), .B2(KEYINPUT3), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT82), .ZN(new_n521));
  INV_X1    g320(.A(new_n509), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT82), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n385), .C1(new_n519), .C2(KEYINPUT3), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT29), .B1(new_n418), .B2(new_n438), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT83), .B1(new_n526), .B2(new_n282), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT83), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n517), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n508), .B(new_n518), .C1(new_n525), .C2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n509), .B1(new_n520), .B2(KEYINPUT82), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(new_n524), .A3(new_n527), .A4(new_n529), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n508), .B1(new_n534), .B2(new_n518), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n507), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n506), .B(new_n531), .C1(new_n535), .C2(KEYINPUT84), .ZN(new_n537));
  INV_X1    g336(.A(new_n517), .ZN(new_n538));
  OAI22_X1  g337(.A1(new_n431), .A2(new_n432), .B1(new_n519), .B2(KEYINPUT3), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n522), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n527), .A2(new_n529), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT84), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n543), .A2(new_n544), .A3(new_n508), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n536), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT85), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n536), .B(new_n548), .C1(new_n537), .C2(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n503), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT35), .B1(new_n470), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n503), .A2(new_n550), .A3(new_n365), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n462), .A2(new_n464), .ZN(new_n557));
  OAI22_X1  g356(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n467), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n556), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT40), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT39), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n425), .B2(new_n367), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n454), .B2(new_n367), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n487), .A2(new_n488), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT4), .B1(new_n568), .B2(new_n433), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n565), .B(new_n437), .C1(new_n569), .C2(new_n452), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n570), .A3(new_n461), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n467), .B1(new_n564), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n567), .A2(new_n570), .A3(KEYINPUT40), .A4(new_n461), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n362), .A3(new_n364), .A4(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n575));
  AOI21_X1  g374(.A(KEYINPUT37), .B1(new_n351), .B2(new_n354), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n360), .B1(new_n355), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT89), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(KEYINPUT89), .B(new_n360), .C1(new_n355), .C2(new_n577), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n360), .A2(new_n575), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT86), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT37), .B1(new_n350), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n347), .A2(new_n584), .A3(new_n350), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n355), .A2(new_n577), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n588), .A2(new_n589), .B1(new_n355), .B2(new_n358), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n469), .A2(KEYINPUT88), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n446), .A2(new_n456), .ZN(new_n592));
  INV_X1    g391(.A(new_n461), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(new_n464), .A3(new_n462), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n590), .A2(new_n560), .A3(new_n591), .A4(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n550), .B(new_n574), .C1(new_n582), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n550), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n466), .A2(new_n467), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n469), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n365), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT74), .B1(new_n501), .B2(new_n502), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(KEYINPUT74), .B(KEYINPUT36), .C1(new_n501), .C2(new_n502), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n597), .A2(new_n603), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n270), .B1(new_n563), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT8), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n615));
  OR2_X1    g414(.A1(G85gat), .A2(G92gat), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n612), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  AND2_X1   g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G99gat), .ZN(new_n624));
  INV_X1    g423(.A(G106gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(KEYINPUT96), .A3(new_n613), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n619), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n628), .B(new_n612), .C1(new_n617), .C2(new_n618), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G57gat), .B(G64gat), .Z(new_n633));
  INV_X1    g432(.A(G71gat), .ZN(new_n634));
  INV_X1    g433(.A(G78gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G71gat), .A2(G78gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT9), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G57gat), .B(G64gat), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n637), .B(new_n636), .C1(new_n642), .C2(new_n639), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n631), .B2(KEYINPUT98), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n632), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n630), .B(new_n631), .C1(KEYINPUT98), .C2(new_n644), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT10), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n632), .A2(new_n649), .A3(new_n644), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n610), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n646), .A2(new_n647), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(G230gat), .A3(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n610), .B(KEYINPUT99), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n648), .B2(new_n650), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n653), .ZN(new_n662));
  INV_X1    g461(.A(new_n656), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI211_X1 g463(.A(KEYINPUT100), .B(new_n656), .C1(new_n661), .C2(new_n653), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n657), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G190gat), .B(G218gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n632), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n243), .B2(new_n245), .ZN(new_n670));
  AND2_X1   g469(.A1(G232gat), .A2(G233gat), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n242), .A2(new_n669), .B1(KEYINPUT41), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n668), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n632), .B1(new_n250), .B2(new_n251), .ZN(new_n676));
  INV_X1    g475(.A(new_n668), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n672), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n671), .A2(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g478(.A(G134gat), .B(G162gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n674), .A2(new_n675), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(KEYINPUT97), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n684), .A2(new_n681), .B1(new_n674), .B2(new_n678), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT21), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n644), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G127gat), .B(G155gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n219), .B1(new_n687), .B2(new_n644), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(G231gat), .A2(G233gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT94), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(G183gat), .B(G211gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n692), .B(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n667), .A2(new_n686), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n609), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n557), .A2(KEYINPUT80), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n594), .A3(new_n600), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n555), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n213), .ZN(G1324gat));
  INV_X1    g508(.A(new_n704), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT16), .B(G8gat), .Z(new_n711));
  NAND4_X1  g510(.A1(new_n710), .A2(KEYINPUT42), .A3(new_n602), .A4(new_n711), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n704), .A2(KEYINPUT102), .A3(new_n365), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT102), .B1(new_n704), .B2(new_n365), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(G8gat), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n711), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n713), .B2(new_n714), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n712), .B(new_n715), .C1(new_n717), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g517(.A1(new_n606), .A2(new_n607), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G15gat), .B1(new_n704), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n503), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(G15gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n704), .B2(new_n723), .ZN(G1326gat));
  NOR2_X1   g523(.A1(new_n704), .A2(new_n550), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT103), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  NAND2_X1  g527(.A1(new_n667), .A2(new_n699), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n686), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT104), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n609), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n707), .A2(G29gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n265), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n729), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n686), .B1(new_n563), .B2(new_n608), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n683), .B2(new_n685), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n684), .A2(new_n681), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n674), .A2(new_n678), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(KEYINPUT106), .A3(new_n682), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  AOI211_X1 g550(.A(KEYINPUT44), .B(new_n751), .C1(new_n563), .C2(new_n608), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n741), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G29gat), .B1(new_n753), .B2(new_n707), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n735), .A2(KEYINPUT45), .A3(new_n736), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n754), .A3(new_n755), .ZN(G1328gat));
  OAI21_X1  g555(.A(G36gat), .B1(new_n753), .B2(new_n365), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n732), .A2(new_n229), .A3(new_n602), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n757), .B(new_n761), .C1(new_n759), .C2(new_n758), .ZN(G1329gat));
  OAI21_X1  g561(.A(G43gat), .B1(new_n753), .B2(new_n720), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n722), .A2(G43gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n609), .A2(new_n731), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT109), .ZN(new_n767));
  OR2_X1    g566(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n763), .A2(new_n766), .A3(new_n768), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n764), .A2(new_n769), .B1(new_n770), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g570(.A(G50gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n732), .A2(new_n772), .A3(new_n598), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n598), .B(new_n741), .C1(new_n744), .C2(new_n752), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n775), .B2(new_n772), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1331gat));
  NAND2_X1  g577(.A1(new_n563), .A2(new_n608), .ZN(new_n779));
  INV_X1    g578(.A(new_n686), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n667), .A2(new_n780), .A3(new_n265), .A4(new_n699), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n601), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g584(.A1(new_n782), .A2(new_n365), .ZN(new_n786));
  NOR2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  AND2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n786), .B2(new_n787), .ZN(G1333gat));
  OAI21_X1  g589(.A(G71gat), .B1(new_n782), .B2(new_n720), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n503), .A2(new_n634), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1334gat));
  NOR2_X1   g594(.A1(new_n782), .A2(new_n550), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(new_n635), .ZN(G1335gat));
  NOR3_X1   g596(.A1(new_n707), .A2(G85gat), .A3(new_n667), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n571), .A2(new_n564), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n594), .A3(new_n573), .ZN(new_n801));
  INV_X1    g600(.A(new_n549), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n544), .B1(new_n543), .B2(new_n508), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n531), .A2(new_n506), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n548), .B1(new_n806), .B2(new_n536), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n365), .A2(new_n801), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n580), .A2(new_n581), .ZN(new_n809));
  INV_X1    g608(.A(new_n575), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n347), .A2(new_n584), .A3(new_n350), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n360), .B(new_n575), .C1(new_n812), .C2(new_n585), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n359), .B1(new_n813), .B2(new_n576), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n469), .A2(KEYINPUT88), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n558), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n808), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n550), .B1(new_n707), .B2(new_n365), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n719), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n707), .A2(new_n503), .A3(new_n550), .A4(new_n365), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n820), .A2(KEYINPUT35), .B1(new_n553), .B2(new_n561), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT112), .B(new_n780), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n700), .A2(new_n265), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT112), .B1(new_n779), .B2(new_n780), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n799), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n823), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n742), .B2(KEYINPUT112), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n780), .B1(new_n819), .B2(new_n821), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n831), .A3(KEYINPUT51), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n826), .A2(KEYINPUT113), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT113), .B1(new_n826), .B2(new_n832), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n798), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n823), .A2(new_n666), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT111), .Z(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n744), .B2(new_n752), .ZN(new_n838));
  OAI21_X1  g637(.A(G85gat), .B1(new_n838), .B2(new_n707), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(G1336gat));
  NAND2_X1  g639(.A1(new_n602), .A2(new_n666), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(G92gat), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n824), .A2(new_n799), .A3(new_n825), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT51), .B1(new_n828), .B2(new_n831), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n602), .B(new_n837), .C1(new_n744), .C2(new_n752), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n847), .A2(G92gat), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n845), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(G1337gat));
  NOR3_X1   g650(.A1(new_n722), .A2(G99gat), .A3(new_n667), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n833), .B2(new_n834), .ZN(new_n853));
  OAI21_X1  g652(.A(G99gat), .B1(new_n838), .B2(new_n720), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1338gat));
  OAI211_X1 g654(.A(new_n598), .B(new_n837), .C1(new_n744), .C2(new_n752), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n625), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n550), .A2(G106gat), .A3(new_n667), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n826), .B2(new_n832), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT53), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n843), .B2(new_n844), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n863), .B(new_n864), .C1(new_n625), .C2(new_n857), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1339gat));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n660), .C1(new_n648), .C2(new_n650), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(new_n663), .ZN(new_n869));
  INV_X1    g668(.A(new_n650), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n659), .C1(new_n652), .C2(KEYINPUT10), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(KEYINPUT54), .A3(new_n651), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n869), .A2(KEYINPUT55), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT55), .B1(new_n869), .B2(new_n872), .ZN(new_n874));
  INV_X1    g673(.A(new_n657), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n207), .B1(new_n252), .B2(new_n247), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n259), .A2(new_n208), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n205), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n264), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n876), .A2(new_n750), .A3(new_n746), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n869), .A2(new_n872), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n869), .A2(KEYINPUT55), .A3(new_n872), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n884), .A2(new_n265), .A3(new_n657), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n666), .A2(new_n880), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n751), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n881), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n701), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n890), .A2(new_n699), .B1(new_n740), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n707), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n553), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n398), .A3(new_n265), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n892), .A2(new_n598), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n707), .A2(new_n602), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n503), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G113gat), .B1(new_n899), .B2(new_n270), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(G1340gat));
  NAND3_X1  g702(.A1(new_n895), .A2(new_n396), .A3(new_n666), .ZN(new_n904));
  OAI21_X1  g703(.A(G120gat), .B1(new_n899), .B2(new_n667), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT116), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT116), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1341gat));
  NAND3_X1  g707(.A1(new_n895), .A2(new_n407), .A3(new_n700), .ZN(new_n909));
  OAI21_X1  g708(.A(G127gat), .B1(new_n899), .B2(new_n699), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1342gat));
  NOR4_X1   g710(.A1(new_n894), .A2(new_n406), .A3(new_n405), .A4(new_n686), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT56), .ZN(new_n913));
  OAI21_X1  g712(.A(G134gat), .B1(new_n899), .B2(new_n686), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(KEYINPUT117), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(KEYINPUT117), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1343gat));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n719), .A2(new_n550), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n893), .A2(new_n365), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n270), .A2(G141gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n720), .A2(new_n898), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n550), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n874), .A2(new_n875), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n256), .A2(new_n264), .A3(KEYINPUT93), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT93), .B1(new_n256), .B2(new_n264), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n928), .B(new_n885), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n780), .B1(new_n931), .B2(new_n887), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n880), .A3(new_n885), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n751), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n927), .B(new_n699), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n891), .A2(new_n740), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n269), .A2(new_n876), .B1(new_n666), .B2(new_n880), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n881), .B1(new_n938), .B2(new_n780), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n927), .B1(new_n939), .B2(new_n699), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n926), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n925), .B1(new_n892), .B2(new_n550), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n924), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(new_n269), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n918), .B(new_n923), .C1(new_n944), .C2(new_n377), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  INV_X1    g745(.A(new_n924), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n265), .A3(new_n947), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n948), .A2(G141gat), .B1(new_n921), .B2(new_n922), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(KEYINPUT119), .A3(new_n918), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n951));
  AOI211_X1 g750(.A(new_n740), .B(new_n924), .C1(new_n941), .C2(new_n942), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n923), .B1(new_n952), .B2(new_n377), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(KEYINPUT58), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n945), .B1(new_n950), .B2(new_n954), .ZN(G1344gat));
  NAND3_X1  g754(.A1(new_n921), .A2(new_n375), .A3(new_n666), .ZN(new_n956));
  XNOR2_X1  g755(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n703), .A2(new_n270), .ZN(new_n958));
  INV_X1    g757(.A(new_n932), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n780), .A2(new_n876), .A3(new_n880), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n700), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n925), .B(new_n598), .C1(new_n958), .C2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT57), .B1(new_n892), .B2(new_n550), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n666), .A3(new_n947), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n957), .B1(new_n965), .B2(G148gat), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT59), .B(new_n375), .C1(new_n943), .C2(new_n666), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n956), .B1(new_n966), .B2(new_n967), .ZN(G1345gat));
  NAND3_X1  g767(.A1(new_n921), .A2(new_n369), .A3(new_n700), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n943), .A2(new_n700), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(new_n369), .ZN(G1346gat));
  AOI21_X1  g770(.A(G162gat), .B1(new_n921), .B2(new_n780), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n751), .A2(new_n370), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n943), .B2(new_n973), .ZN(G1347gat));
  NAND3_X1  g773(.A1(new_n707), .A2(new_n602), .A3(new_n503), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT121), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n897), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n977), .A2(new_n305), .A3(new_n270), .ZN(new_n978));
  NOR4_X1   g777(.A1(new_n892), .A2(new_n601), .A3(new_n365), .A4(new_n551), .ZN(new_n979));
  AOI21_X1  g778(.A(G169gat), .B1(new_n979), .B2(new_n265), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n978), .A2(new_n980), .ZN(G1348gat));
  OR3_X1    g780(.A1(new_n977), .A2(new_n325), .A3(new_n667), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(KEYINPUT122), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(KEYINPUT122), .ZN(new_n984));
  AOI21_X1  g783(.A(G176gat), .B1(new_n979), .B2(new_n666), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(G1349gat));
  AND2_X1   g785(.A1(new_n700), .A2(new_n334), .ZN(new_n987));
  AOI22_X1  g786(.A1(new_n979), .A2(new_n987), .B1(KEYINPUT123), .B2(KEYINPUT60), .ZN(new_n988));
  OAI21_X1  g787(.A(G183gat), .B1(new_n977), .B2(new_n699), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g789(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n990), .B(new_n991), .Z(G1350gat));
  NAND3_X1  g791(.A1(new_n979), .A2(new_n333), .A3(new_n889), .ZN(new_n993));
  OAI21_X1  g792(.A(G190gat), .B1(new_n977), .B2(new_n686), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(G1351gat));
  NOR2_X1   g796(.A1(new_n892), .A2(new_n601), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(new_n919), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n999), .A2(new_n365), .ZN(new_n1000));
  XNOR2_X1  g799(.A(KEYINPUT124), .B(G197gat), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n740), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n719), .A2(new_n601), .A3(new_n365), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n964), .A2(new_n269), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT125), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(G1352gat));
  NOR3_X1   g808(.A1(new_n999), .A2(G204gat), .A3(new_n841), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT62), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n964), .A2(new_n666), .A3(new_n1004), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(G204gat), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1011), .A2(new_n1013), .ZN(G1353gat));
  NOR4_X1   g813(.A1(new_n999), .A2(G211gat), .A3(new_n365), .A4(new_n699), .ZN(new_n1015));
  XOR2_X1   g814(.A(new_n1015), .B(KEYINPUT126), .Z(new_n1016));
  NAND3_X1  g815(.A1(new_n964), .A2(new_n700), .A3(new_n1004), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(G211gat), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(KEYINPUT63), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT63), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1017), .A2(new_n1020), .A3(G211gat), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1016), .A2(new_n1019), .A3(new_n1021), .ZN(G1354gat));
  INV_X1    g821(.A(G218gat), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1000), .A2(new_n1023), .A3(new_n889), .ZN(new_n1024));
  NAND4_X1  g823(.A1(new_n962), .A2(new_n780), .A3(new_n963), .A4(new_n1004), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1025), .A2(G218gat), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g826(.A(new_n1027), .B(KEYINPUT127), .Z(G1355gat));
endmodule


