

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n711), .A2(G1996), .ZN(n683) );
  NOR2_X1 U550 ( .A1(n690), .A2(n1008), .ZN(n689) );
  XOR2_X1 U551 ( .A(KEYINPUT98), .B(n726), .Z(n516) );
  AND2_X1 U552 ( .A1(n687), .A2(n686), .ZN(n690) );
  INV_X1 U553 ( .A(KEYINPUT96), .ZN(n688) );
  XNOR2_X1 U554 ( .A(n689), .B(n688), .ZN(n696) );
  AND2_X1 U555 ( .A1(G160), .A2(n682), .ZN(n711) );
  XNOR2_X1 U556 ( .A(n550), .B(KEYINPUT13), .ZN(n551) );
  NOR2_X1 U557 ( .A1(n628), .A2(n538), .ZN(n638) );
  XNOR2_X1 U558 ( .A(n552), .B(n551), .ZN(n555) );
  XOR2_X1 U559 ( .A(KEYINPUT17), .B(n523), .Z(n983) );
  OR2_X1 U560 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X2 U561 ( .A1(n528), .A2(n527), .ZN(G160) );
  INV_X1 U562 ( .A(G2104), .ZN(n519) );
  NOR2_X4 U563 ( .A1(n519), .A2(G2105), .ZN(n984) );
  NAND2_X1 U564 ( .A1(n984), .A2(G101), .ZN(n517) );
  XNOR2_X1 U565 ( .A(n517), .B(KEYINPUT65), .ZN(n518) );
  XNOR2_X1 U566 ( .A(n518), .B(KEYINPUT23), .ZN(n521) );
  AND2_X1 U567 ( .A1(n519), .A2(G2105), .ZN(n980) );
  NAND2_X1 U568 ( .A1(G125), .A2(n980), .ZN(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U570 ( .A(KEYINPUT66), .B(n522), .ZN(n528) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  AND2_X1 U572 ( .A1(n983), .A2(G137), .ZN(n526) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n979) );
  NAND2_X1 U574 ( .A1(G113), .A2(n979), .ZN(n524) );
  XNOR2_X1 U575 ( .A(KEYINPUT67), .B(n524), .ZN(n525) );
  XNOR2_X1 U576 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U577 ( .A1(G138), .A2(n983), .ZN(n533) );
  AND2_X1 U578 ( .A1(G102), .A2(n984), .ZN(n532) );
  NAND2_X1 U579 ( .A1(G114), .A2(n979), .ZN(n530) );
  NAND2_X1 U580 ( .A1(G126), .A2(n980), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n679) );
  AND2_X1 U583 ( .A1(n533), .A2(n679), .ZN(G164) );
  AND2_X1 U584 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U585 ( .A(G132), .ZN(G219) );
  INV_X1 U586 ( .A(G120), .ZN(G236) );
  INV_X1 U587 ( .A(G69), .ZN(G235) );
  INV_X1 U588 ( .A(G108), .ZN(G238) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NOR2_X1 U590 ( .A1(G651), .A2(n628), .ZN(n641) );
  NAND2_X1 U591 ( .A1(G52), .A2(n641), .ZN(n536) );
  INV_X1 U592 ( .A(G651), .ZN(n538) );
  NOR2_X1 U593 ( .A1(G543), .A2(n538), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n534), .Z(n644) );
  NAND2_X1 U595 ( .A1(G64), .A2(n644), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n640) );
  NAND2_X1 U598 ( .A1(n640), .A2(G90), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT69), .B(n537), .Z(n540) );
  NAND2_X1 U600 ( .A1(n638), .A2(G77), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U603 ( .A1(n543), .A2(n542), .ZN(G171) );
  NAND2_X1 U604 ( .A1(G7), .A2(G661), .ZN(n544) );
  XOR2_X1 U605 ( .A(n544), .B(KEYINPUT10), .Z(n1020) );
  NAND2_X1 U606 ( .A1(n1020), .A2(G567), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT11), .B(n545), .Z(G234) );
  NAND2_X1 U608 ( .A1(n644), .A2(G56), .ZN(n546) );
  XNOR2_X1 U609 ( .A(KEYINPUT14), .B(n546), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n640), .A2(G81), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(KEYINPUT12), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G68), .A2(n638), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n552) );
  XNOR2_X1 U614 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n550) );
  NAND2_X1 U615 ( .A1(G43), .A2(n641), .ZN(n553) );
  XNOR2_X1 U616 ( .A(KEYINPUT75), .B(n553), .ZN(n554) );
  NOR2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n1007) );
  INV_X1 U619 ( .A(G860), .ZN(n591) );
  OR2_X1 U620 ( .A1(n1007), .A2(n591), .ZN(G153) );
  NAND2_X1 U621 ( .A1(G92), .A2(n640), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G66), .A2(n644), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G79), .A2(n638), .ZN(n561) );
  NAND2_X1 U625 ( .A1(G54), .A2(n641), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT15), .B(n564), .Z(n1008) );
  NOR2_X1 U629 ( .A1(n1008), .A2(G868), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT76), .ZN(n567) );
  INV_X1 U631 ( .A(G868), .ZN(n658) );
  NOR2_X1 U632 ( .A1(n658), .A2(G171), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT77), .B(n568), .ZN(G284) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G65), .A2(n644), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT70), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G78), .A2(n638), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G91), .A2(n640), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G53), .A2(n641), .ZN(n572) );
  XNOR2_X1 U642 ( .A(KEYINPUT71), .B(n572), .ZN(n573) );
  NOR2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(G299) );
  NAND2_X1 U645 ( .A1(G89), .A2(n640), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n577), .B(KEYINPUT4), .ZN(n578) );
  XNOR2_X1 U647 ( .A(n578), .B(KEYINPUT78), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G76), .A2(n638), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U650 ( .A(n581), .B(KEYINPUT5), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G51), .A2(n641), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G63), .A2(n644), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT6), .B(n584), .Z(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n587), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U657 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U658 ( .A(G299), .ZN(n703) );
  NAND2_X1 U659 ( .A1(n703), .A2(n658), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n588), .B(KEYINPUT79), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n658), .A2(G286), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U663 ( .A1(n591), .A2(G559), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n592), .A2(n1008), .ZN(n593) );
  XNOR2_X1 U665 ( .A(n593), .B(KEYINPUT16), .ZN(n594) );
  XNOR2_X1 U666 ( .A(KEYINPUT80), .B(n594), .ZN(G148) );
  NOR2_X1 U667 ( .A1(G868), .A2(n1007), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G868), .A2(n1008), .ZN(n595) );
  NOR2_X1 U669 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U671 ( .A1(n980), .A2(G123), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n598), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G99), .A2(n984), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G111), .A2(n979), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G135), .A2(n983), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n998) );
  XNOR2_X1 U679 ( .A(n998), .B(G2096), .ZN(n605) );
  INV_X1 U680 ( .A(G2100), .ZN(n959) );
  NAND2_X1 U681 ( .A1(n605), .A2(n959), .ZN(G156) );
  NAND2_X1 U682 ( .A1(G55), .A2(n641), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G67), .A2(n644), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U685 ( .A(KEYINPUT83), .B(n608), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n638), .A2(G80), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G93), .A2(n640), .ZN(n609) );
  AND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n657) );
  NAND2_X1 U690 ( .A1(G559), .A2(n1008), .ZN(n613) );
  XOR2_X1 U691 ( .A(n1007), .B(n613), .Z(n655) );
  XNOR2_X1 U692 ( .A(KEYINPUT81), .B(n655), .ZN(n614) );
  NOR2_X1 U693 ( .A1(G860), .A2(n614), .ZN(n615) );
  XOR2_X1 U694 ( .A(n657), .B(n615), .Z(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT82), .ZN(G145) );
  NAND2_X1 U696 ( .A1(G85), .A2(n640), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G60), .A2(n644), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G72), .A2(n638), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G47), .A2(n641), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT68), .B(n623), .Z(G290) );
  NAND2_X1 U704 ( .A1(G49), .A2(n641), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U707 ( .A(KEYINPUT84), .B(n626), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n644), .A2(n627), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G75), .A2(n638), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G50), .A2(n641), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G88), .A2(n640), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G62), .A2(n644), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U718 ( .A(n637), .B(KEYINPUT86), .Z(G303) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  NAND2_X1 U720 ( .A1(n638), .A2(G73), .ZN(n639) );
  XNOR2_X1 U721 ( .A(n639), .B(KEYINPUT2), .ZN(n649) );
  NAND2_X1 U722 ( .A1(G86), .A2(n640), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G48), .A2(n641), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G61), .A2(n644), .ZN(n645) );
  XNOR2_X1 U726 ( .A(KEYINPUT85), .B(n645), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U729 ( .A(G290), .B(KEYINPUT19), .ZN(n651) );
  XOR2_X1 U730 ( .A(G288), .B(G166), .Z(n650) );
  XNOR2_X1 U731 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U732 ( .A(n657), .B(n652), .Z(n654) );
  XOR2_X1 U733 ( .A(G305), .B(G299), .Z(n653) );
  XNOR2_X1 U734 ( .A(n654), .B(n653), .ZN(n1006) );
  XNOR2_X1 U735 ( .A(n655), .B(n1006), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n664), .A2(G2072), .ZN(n665) );
  XOR2_X1 U744 ( .A(KEYINPUT87), .B(n665), .Z(G158) );
  XOR2_X1 U745 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U746 ( .A1(G235), .A2(G236), .ZN(n666) );
  XOR2_X1 U747 ( .A(KEYINPUT88), .B(n666), .Z(n667) );
  NOR2_X1 U748 ( .A1(G238), .A2(n667), .ZN(n668) );
  NAND2_X1 U749 ( .A1(G57), .A2(n668), .ZN(n946) );
  NAND2_X1 U750 ( .A1(G567), .A2(n946), .ZN(n669) );
  XNOR2_X1 U751 ( .A(n669), .B(KEYINPUT89), .ZN(n674) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n670) );
  XNOR2_X1 U753 ( .A(KEYINPUT22), .B(n670), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n671), .A2(G96), .ZN(n672) );
  OR2_X1 U755 ( .A1(G218), .A2(n672), .ZN(n947) );
  AND2_X1 U756 ( .A1(G2106), .A2(n947), .ZN(n673) );
  NOR2_X1 U757 ( .A1(n674), .A2(n673), .ZN(G319) );
  INV_X1 U758 ( .A(G319), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U760 ( .A1(n676), .A2(n675), .ZN(n823) );
  NAND2_X1 U761 ( .A1(n823), .A2(G36), .ZN(G176) );
  INV_X1 U762 ( .A(G1384), .ZN(n677) );
  AND2_X1 U763 ( .A1(G138), .A2(n677), .ZN(n678) );
  NAND2_X1 U764 ( .A1(n983), .A2(n678), .ZN(n681) );
  OR2_X1 U765 ( .A1(G1384), .A2(n679), .ZN(n680) );
  NAND2_X1 U766 ( .A1(n681), .A2(n680), .ZN(n774) );
  AND2_X1 U767 ( .A1(n774), .A2(G40), .ZN(n682) );
  XOR2_X1 U768 ( .A(KEYINPUT26), .B(n683), .Z(n687) );
  INV_X1 U769 ( .A(n711), .ZN(n727) );
  NAND2_X1 U770 ( .A1(n727), .A2(G1341), .ZN(n685) );
  INV_X1 U771 ( .A(n1007), .ZN(n684) );
  AND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n1008), .A2(n690), .ZN(n694) );
  XNOR2_X1 U774 ( .A(n711), .B(KEYINPUT94), .ZN(n698) );
  NAND2_X1 U775 ( .A1(G2067), .A2(n698), .ZN(n692) );
  NAND2_X1 U776 ( .A1(G1348), .A2(n727), .ZN(n691) );
  NAND2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n696), .A2(n695), .ZN(n702) );
  NAND2_X1 U780 ( .A1(G2072), .A2(n698), .ZN(n697) );
  XNOR2_X1 U781 ( .A(n697), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U782 ( .A(n698), .ZN(n710) );
  AND2_X1 U783 ( .A1(n710), .A2(G1956), .ZN(n699) );
  NOR2_X1 U784 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U785 ( .A1(n703), .A2(n704), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n702), .A2(n701), .ZN(n708) );
  NOR2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n706) );
  XNOR2_X1 U788 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n705) );
  XNOR2_X1 U789 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U790 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U791 ( .A(n709), .B(KEYINPUT29), .ZN(n715) );
  XOR2_X1 U792 ( .A(G2078), .B(KEYINPUT25), .Z(n837) );
  NOR2_X1 U793 ( .A1(n837), .A2(n710), .ZN(n713) );
  NOR2_X1 U794 ( .A1(n711), .A2(G1961), .ZN(n712) );
  NOR2_X1 U795 ( .A1(n713), .A2(n712), .ZN(n720) );
  NOR2_X1 U796 ( .A1(G301), .A2(n720), .ZN(n714) );
  NOR2_X1 U797 ( .A1(n715), .A2(n714), .ZN(n725) );
  XNOR2_X1 U798 ( .A(KEYINPUT97), .B(KEYINPUT30), .ZN(n718) );
  NAND2_X1 U799 ( .A1(G8), .A2(n727), .ZN(n798) );
  NOR2_X1 U800 ( .A1(G1966), .A2(n798), .ZN(n736) );
  NOR2_X1 U801 ( .A1(G2084), .A2(n727), .ZN(n735) );
  NOR2_X1 U802 ( .A1(n736), .A2(n735), .ZN(n716) );
  NAND2_X1 U803 ( .A1(n716), .A2(G8), .ZN(n717) );
  XOR2_X1 U804 ( .A(n718), .B(n717), .Z(n719) );
  NOR2_X1 U805 ( .A1(G168), .A2(n719), .ZN(n722) );
  AND2_X1 U806 ( .A1(G301), .A2(n720), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U808 ( .A(n723), .B(KEYINPUT31), .ZN(n724) );
  NOR2_X1 U809 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U810 ( .A1(G286), .A2(n516), .ZN(n732) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n798), .ZN(n729) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U814 ( .A1(n730), .A2(G303), .ZN(n731) );
  NAND2_X1 U815 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U816 ( .A1(n733), .A2(G8), .ZN(n734) );
  XNOR2_X1 U817 ( .A(KEYINPUT32), .B(n734), .ZN(n790) );
  NAND2_X1 U818 ( .A1(G8), .A2(n735), .ZN(n739) );
  XNOR2_X1 U819 ( .A(n516), .B(KEYINPUT99), .ZN(n737) );
  NOR2_X1 U820 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U821 ( .A1(n739), .A2(n738), .ZN(n791) );
  INV_X1 U822 ( .A(n798), .ZN(n740) );
  NAND2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n883) );
  AND2_X1 U824 ( .A1(n740), .A2(n883), .ZN(n742) );
  AND2_X1 U825 ( .A1(n791), .A2(n742), .ZN(n741) );
  NAND2_X1 U826 ( .A1(n790), .A2(n741), .ZN(n746) );
  INV_X1 U827 ( .A(n742), .ZN(n744) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U829 ( .A1(G303), .A2(G1971), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n749), .A2(n743), .ZN(n887) );
  OR2_X1 U831 ( .A1(n744), .A2(n887), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U833 ( .A(n747), .B(KEYINPUT64), .ZN(n748) );
  NOR2_X1 U834 ( .A1(KEYINPUT33), .A2(n748), .ZN(n753) );
  NAND2_X1 U835 ( .A1(KEYINPUT33), .A2(n749), .ZN(n750) );
  XNOR2_X1 U836 ( .A(KEYINPUT100), .B(n750), .ZN(n751) );
  NOR2_X1 U837 ( .A1(n798), .A2(n751), .ZN(n752) );
  NOR2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n789) );
  XNOR2_X1 U839 ( .A(KEYINPUT101), .B(G1981), .ZN(n754) );
  XNOR2_X1 U840 ( .A(n754), .B(G305), .ZN(n889) );
  XOR2_X1 U841 ( .A(G1986), .B(G290), .Z(n880) );
  XOR2_X1 U842 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n756) );
  NAND2_X1 U843 ( .A1(G105), .A2(n984), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n756), .B(n755), .ZN(n760) );
  NAND2_X1 U845 ( .A1(G129), .A2(n980), .ZN(n758) );
  NAND2_X1 U846 ( .A1(G141), .A2(n983), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n979), .A2(G117), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n999) );
  NAND2_X1 U851 ( .A1(G1996), .A2(n999), .ZN(n771) );
  NAND2_X1 U852 ( .A1(G119), .A2(n980), .ZN(n764) );
  NAND2_X1 U853 ( .A1(G95), .A2(n984), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n767) );
  NAND2_X1 U855 ( .A1(G131), .A2(n983), .ZN(n765) );
  XNOR2_X1 U856 ( .A(KEYINPUT91), .B(n765), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n979), .A2(G107), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n992) );
  NAND2_X1 U860 ( .A1(G1991), .A2(n992), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n907) );
  INV_X1 U862 ( .A(n907), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n880), .A2(n772), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G160), .A2(G40), .ZN(n773) );
  NOR2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n814) );
  NAND2_X1 U866 ( .A1(n775), .A2(n814), .ZN(n786) );
  NAND2_X1 U867 ( .A1(G140), .A2(n983), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G104), .A2(n984), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U870 ( .A(KEYINPUT34), .B(n778), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n979), .A2(G116), .ZN(n779) );
  XNOR2_X1 U872 ( .A(n779), .B(KEYINPUT90), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G128), .A2(n980), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U875 ( .A(KEYINPUT35), .B(n782), .Z(n783) );
  NOR2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U877 ( .A(KEYINPUT36), .B(n785), .ZN(n995) );
  XNOR2_X1 U878 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NOR2_X1 U879 ( .A1(n995), .A2(n811), .ZN(n908) );
  NAND2_X1 U880 ( .A1(n908), .A2(n814), .ZN(n809) );
  NAND2_X1 U881 ( .A1(n786), .A2(n809), .ZN(n803) );
  INV_X1 U882 ( .A(n803), .ZN(n787) );
  AND2_X1 U883 ( .A1(n889), .A2(n787), .ZN(n788) );
  AND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n819) );
  NAND2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n794) );
  NOR2_X1 U886 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  AND2_X1 U889 ( .A1(n798), .A2(n795), .ZN(n801) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U891 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  NOR2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT93), .B(n799), .Z(n800) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  OR2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n817) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n999), .ZN(n926) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n992), .ZN(n933) );
  NOR2_X1 U899 ( .A1(n804), .A2(n933), .ZN(n805) );
  XNOR2_X1 U900 ( .A(n805), .B(KEYINPUT102), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n907), .A2(n806), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n926), .A2(n807), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n995), .A2(n811), .ZN(n922) );
  NAND2_X1 U906 ( .A1(n812), .A2(n922), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U908 ( .A(n815), .B(KEYINPUT103), .Z(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U911 ( .A(KEYINPUT40), .B(n820), .Z(G329) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n1020), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U914 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(G188) );
  NAND2_X1 U918 ( .A1(n980), .A2(G124), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(KEYINPUT44), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G136), .A2(n983), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT109), .ZN(n829) );
  NAND2_X1 U923 ( .A1(G100), .A2(n984), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n979), .A2(G112), .ZN(n830) );
  XOR2_X1 U926 ( .A(KEYINPUT110), .B(n830), .Z(n831) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(G162) );
  INV_X1 U928 ( .A(KEYINPUT55), .ZN(n940) );
  XNOR2_X1 U929 ( .A(G2084), .B(G34), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n833), .B(KEYINPUT54), .ZN(n849) );
  XNOR2_X1 U931 ( .A(G2090), .B(G35), .ZN(n846) );
  XOR2_X1 U932 ( .A(G1991), .B(G25), .Z(n834) );
  NAND2_X1 U933 ( .A1(n834), .A2(G28), .ZN(n843) );
  XNOR2_X1 U934 ( .A(G2067), .B(G26), .ZN(n836) );
  XNOR2_X1 U935 ( .A(G33), .B(G2072), .ZN(n835) );
  NOR2_X1 U936 ( .A1(n836), .A2(n835), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n837), .B(G27), .ZN(n839) );
  XNOR2_X1 U938 ( .A(G1996), .B(G32), .ZN(n838) );
  NOR2_X1 U939 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U940 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U942 ( .A(KEYINPUT53), .B(n844), .ZN(n845) );
  NOR2_X1 U943 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT118), .B(n847), .Z(n848) );
  NOR2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n940), .B(n850), .ZN(n851) );
  NOR2_X1 U947 ( .A1(G29), .A2(n851), .ZN(n852) );
  XNOR2_X1 U948 ( .A(KEYINPUT119), .B(n852), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n853), .A2(G11), .ZN(n905) );
  XNOR2_X1 U950 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n854), .B(KEYINPUT123), .ZN(n877) );
  XNOR2_X1 U952 ( .A(G1348), .B(KEYINPUT59), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n855), .B(G4), .ZN(n859) );
  XNOR2_X1 U954 ( .A(G1981), .B(G6), .ZN(n857) );
  XNOR2_X1 U955 ( .A(G1956), .B(G20), .ZN(n856) );
  NOR2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n862) );
  XOR2_X1 U958 ( .A(KEYINPUT121), .B(G1341), .Z(n860) );
  XNOR2_X1 U959 ( .A(G19), .B(n860), .ZN(n861) );
  NOR2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U961 ( .A(KEYINPUT60), .B(n863), .ZN(n867) );
  XNOR2_X1 U962 ( .A(G1966), .B(G21), .ZN(n865) );
  XNOR2_X1 U963 ( .A(G5), .B(G1961), .ZN(n864) );
  NOR2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n866) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n875) );
  XNOR2_X1 U966 ( .A(G1976), .B(G23), .ZN(n869) );
  XNOR2_X1 U967 ( .A(G1971), .B(G22), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n872) );
  XOR2_X1 U969 ( .A(G1986), .B(KEYINPUT122), .Z(n870) );
  XNOR2_X1 U970 ( .A(G24), .B(n870), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(KEYINPUT58), .B(n873), .ZN(n874) );
  NOR2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U975 ( .A1(G16), .A2(n878), .ZN(n902) );
  XOR2_X1 U976 ( .A(G1341), .B(n1007), .Z(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n898) );
  XOR2_X1 U978 ( .A(G1956), .B(G299), .Z(n882) );
  NAND2_X1 U979 ( .A1(G1971), .A2(G303), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n886) );
  XNOR2_X1 U981 ( .A(G1348), .B(n1008), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U983 ( .A1(n886), .A2(n885), .ZN(n896) );
  XOR2_X1 U984 ( .A(G301), .B(G1961), .Z(n888) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n894) );
  XNOR2_X1 U986 ( .A(G1966), .B(G168), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n891), .B(KEYINPUT120), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT57), .B(n892), .Z(n893) );
  NOR2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n895) );
  NAND2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U992 ( .A1(n898), .A2(n897), .ZN(n900) );
  XOR2_X1 U993 ( .A(G16), .B(KEYINPUT56), .Z(n899) );
  NOR2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n901) );
  NOR2_X1 U995 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n903), .B(KEYINPUT125), .ZN(n904) );
  NOR2_X1 U997 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U998 ( .A(n906), .B(KEYINPUT126), .ZN(n944) );
  NOR2_X1 U999 ( .A1(n908), .A2(n907), .ZN(n931) );
  XNOR2_X1 U1000 ( .A(G164), .B(G2078), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n909), .B(KEYINPUT117), .ZN(n920) );
  XNOR2_X1 U1002 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n914) );
  NAND2_X1 U1003 ( .A1(G115), .A2(n979), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(G127), .A2(n980), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n912), .B(KEYINPUT47), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(n914), .B(n913), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n983), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(G103), .A2(n984), .ZN(n915) );
  NAND2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n990) );
  XOR2_X1 U1012 ( .A(G2072), .B(n990), .Z(n919) );
  NOR2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(n921), .B(KEYINPUT50), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n929) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n924) );
  XNOR2_X1 U1017 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NOR2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1019 ( .A(KEYINPUT51), .B(n927), .ZN(n928) );
  NOR2_X1 U1020 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1021 ( .A1(n931), .A2(n930), .ZN(n938) );
  XNOR2_X1 U1022 ( .A(G2084), .B(G160), .ZN(n932) );
  XNOR2_X1 U1023 ( .A(n932), .B(KEYINPUT114), .ZN(n935) );
  NOR2_X1 U1024 ( .A1(n933), .A2(n998), .ZN(n934) );
  NAND2_X1 U1025 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1026 ( .A(KEYINPUT115), .B(n936), .Z(n937) );
  NOR2_X1 U1027 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n939), .ZN(n941) );
  NAND2_X1 U1029 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1030 ( .A1(n942), .A2(G29), .ZN(n943) );
  NAND2_X1 U1031 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1032 ( .A(KEYINPUT62), .B(n945), .Z(G311) );
  XNOR2_X1 U1033 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1034 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1035 ( .A1(n947), .A2(n946), .ZN(G325) );
  INV_X1 U1036 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1037 ( .A(G2443), .B(G1341), .ZN(n956) );
  XNOR2_X1 U1038 ( .A(G2430), .B(G2446), .ZN(n954) );
  XOR2_X1 U1039 ( .A(G2454), .B(G2451), .Z(n949) );
  XNOR2_X1 U1040 ( .A(G2427), .B(G2435), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(n949), .B(n948), .ZN(n950) );
  XOR2_X1 U1042 ( .A(n950), .B(G2438), .Z(n952) );
  XNOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT104), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n952), .B(n951), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(n954), .B(n953), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(n956), .B(n955), .ZN(n957) );
  NAND2_X1 U1047 ( .A1(n957), .A2(G14), .ZN(n958) );
  XOR2_X1 U1048 ( .A(KEYINPUT105), .B(n958), .Z(n1013) );
  XOR2_X1 U1049 ( .A(KEYINPUT106), .B(n1013), .Z(G401) );
  XNOR2_X1 U1050 ( .A(n959), .B(G2096), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G2090), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n961), .B(n960), .ZN(n965) );
  XOR2_X1 U1053 ( .A(G2678), .B(KEYINPUT42), .Z(n963) );
  XNOR2_X1 U1054 ( .A(G2072), .B(KEYINPUT43), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n963), .B(n962), .ZN(n964) );
  XOR2_X1 U1056 ( .A(n965), .B(n964), .Z(n967) );
  XNOR2_X1 U1057 ( .A(G2084), .B(G2078), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n967), .B(n966), .ZN(G227) );
  XOR2_X1 U1059 ( .A(KEYINPUT41), .B(G1996), .Z(n969) );
  XNOR2_X1 U1060 ( .A(G1976), .B(G1961), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1062 ( .A(n970), .B(G2474), .Z(n972) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G1991), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n972), .B(n971), .ZN(n976) );
  XOR2_X1 U1065 ( .A(KEYINPUT108), .B(G1986), .Z(n974) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G1956), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1068 ( .A(n976), .B(n975), .Z(n978) );
  XNOR2_X1 U1069 ( .A(G1971), .B(KEYINPUT107), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n978), .B(n977), .ZN(G229) );
  NAND2_X1 U1071 ( .A1(G118), .A2(n979), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(G130), .A2(n980), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n989) );
  NAND2_X1 U1074 ( .A1(G142), .A2(n983), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(G106), .A2(n984), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1077 ( .A(KEYINPUT45), .B(n987), .Z(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n994) );
  XOR2_X1 U1079 ( .A(G162), .B(n990), .Z(n991) );
  XNOR2_X1 U1080 ( .A(n992), .B(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n994), .B(n993), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(n995), .B(G160), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(n997), .B(n996), .ZN(n1004) );
  XNOR2_X1 U1084 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(n999), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XOR2_X1 U1087 ( .A(G164), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1088 ( .A(n1004), .B(n1003), .ZN(n1005) );
  NOR2_X1 U1089 ( .A1(G37), .A2(n1005), .ZN(G395) );
  XNOR2_X1 U1090 ( .A(n1007), .B(n1006), .ZN(n1010) );
  XOR2_X1 U1091 ( .A(G301), .B(n1008), .Z(n1009) );
  XNOR2_X1 U1092 ( .A(n1010), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(G286), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1094 ( .A1(G37), .A2(n1012), .ZN(G397) );
  NAND2_X1 U1095 ( .A1(G319), .A2(n1013), .ZN(n1017) );
  NOR2_X1 U1096 ( .A1(G227), .A2(G229), .ZN(n1014) );
  XOR2_X1 U1097 ( .A(KEYINPUT113), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1098 ( .A(n1015), .B(KEYINPUT49), .ZN(n1016) );
  NOR2_X1 U1099 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NOR2_X1 U1100 ( .A1(G395), .A2(G397), .ZN(n1018) );
  NAND2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(G225) );
  INV_X1 U1102 ( .A(G225), .ZN(G308) );
  INV_X1 U1103 ( .A(G57), .ZN(G237) );
  INV_X1 U1104 ( .A(n1020), .ZN(G223) );
endmodule

